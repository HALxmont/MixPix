magic
tech sky130A
magscale 1 2
timestamp 1668464426
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 331214 702992 331220 703044
rect 331272 703032 331278 703044
rect 332502 703032 332508 703044
rect 331272 703004 332508 703032
rect 331272 702992 331278 703004
rect 332502 702992 332508 703004
rect 332560 702992 332566 703044
rect 410518 700408 410524 700460
rect 410576 700448 410582 700460
rect 429838 700448 429844 700460
rect 410576 700420 429844 700448
rect 410576 700408 410582 700420
rect 429838 700408 429844 700420
rect 429896 700408 429902 700460
rect 300118 700340 300124 700392
rect 300176 700380 300182 700392
rect 303246 700380 303252 700392
rect 300176 700352 303252 700380
rect 300176 700340 300182 700352
rect 303246 700340 303252 700352
rect 303304 700340 303310 700392
rect 409138 700340 409144 700392
rect 409196 700380 409202 700392
rect 494790 700380 494796 700392
rect 409196 700352 494796 700380
rect 409196 700340 409202 700352
rect 494790 700340 494796 700352
rect 494848 700340 494854 700392
rect 254578 700272 254584 700324
rect 254636 700312 254642 700324
rect 267642 700312 267648 700324
rect 254636 700284 267648 700312
rect 254636 700272 254642 700284
rect 267642 700272 267648 700284
rect 267700 700272 267706 700324
rect 407758 700272 407764 700324
rect 407816 700312 407822 700324
rect 559650 700312 559656 700324
rect 407816 700284 559656 700312
rect 407816 700272 407822 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 348786 699796 348792 699848
rect 348844 699836 348850 699848
rect 351178 699836 351184 699848
rect 348844 699808 351184 699836
rect 348844 699796 348850 699808
rect 351178 699796 351184 699808
rect 351236 699796 351242 699848
rect 152458 699660 152464 699712
rect 152516 699700 152522 699712
rect 154114 699700 154120 699712
rect 152516 699672 154120 699700
rect 152516 699660 152522 699672
rect 154114 699660 154120 699672
rect 154172 699660 154178 699712
rect 196618 699660 196624 699712
rect 196676 699700 196682 699712
rect 202782 699700 202788 699712
rect 196676 699672 202788 699700
rect 196676 699660 196682 699672
rect 202782 699660 202788 699672
rect 202840 699660 202846 699712
rect 217318 699660 217324 699712
rect 217376 699700 217382 699712
rect 218974 699700 218980 699712
rect 217376 699672 218980 699700
rect 217376 699660 217382 699672
rect 218974 699660 218980 699672
rect 219032 699660 219038 699712
rect 282178 697552 282184 697604
rect 282236 697592 282242 697604
rect 283834 697592 283840 697604
rect 282236 697564 283840 697592
rect 282236 697552 282242 697564
rect 283834 697552 283840 697564
rect 283892 697552 283898 697604
rect 303246 693404 303252 693456
rect 303304 693444 303310 693456
rect 316034 693444 316040 693456
rect 303304 693416 316040 693444
rect 303304 693404 303310 693416
rect 316034 693404 316040 693416
rect 316092 693404 316098 693456
rect 351178 692044 351184 692096
rect 351236 692084 351242 692096
rect 358078 692084 358084 692096
rect 351236 692056 358084 692084
rect 351236 692044 351242 692056
rect 358078 692044 358084 692056
rect 358136 692044 358142 692096
rect 364334 690412 364340 690464
rect 364392 690452 364398 690464
rect 369854 690452 369860 690464
rect 364392 690424 369860 690452
rect 364392 690412 364398 690424
rect 369854 690412 369860 690424
rect 369912 690412 369918 690464
rect 150434 689256 150440 689308
rect 150492 689296 150498 689308
rect 152458 689296 152464 689308
rect 150492 689268 152464 689296
rect 150492 689256 150498 689268
rect 152458 689256 152464 689268
rect 152516 689256 152522 689308
rect 239030 689256 239036 689308
rect 239088 689296 239094 689308
rect 254578 689296 254584 689308
rect 239088 689268 254584 689296
rect 239088 689256 239094 689268
rect 254578 689256 254584 689268
rect 254636 689256 254642 689308
rect 331214 688848 331220 688900
rect 331272 688888 331278 688900
rect 334618 688888 334624 688900
rect 331272 688860 334624 688888
rect 331272 688848 331278 688860
rect 334618 688848 334624 688860
rect 334676 688848 334682 688900
rect 217318 688684 217324 688696
rect 215312 688656 217324 688684
rect 213178 688576 213184 688628
rect 213236 688616 213242 688628
rect 215312 688616 215340 688656
rect 217318 688644 217324 688656
rect 217376 688644 217382 688696
rect 213236 688588 215340 688616
rect 213236 688576 213242 688588
rect 316034 688168 316040 688220
rect 316092 688208 316098 688220
rect 323578 688208 323584 688220
rect 316092 688180 323584 688208
rect 316092 688168 316098 688180
rect 323578 688168 323584 688180
rect 323636 688168 323642 688220
rect 369854 688168 369860 688220
rect 369912 688208 369918 688220
rect 372614 688208 372620 688220
rect 369912 688180 372620 688208
rect 369912 688168 369918 688180
rect 372614 688168 372620 688180
rect 372672 688168 372678 688220
rect 224218 685108 224224 685160
rect 224276 685148 224282 685160
rect 239030 685148 239036 685160
rect 224276 685120 239036 685148
rect 224276 685108 224282 685120
rect 239030 685108 239036 685120
rect 239088 685108 239094 685160
rect 2774 683680 2780 683732
rect 2832 683720 2838 683732
rect 4798 683720 4804 683732
rect 2832 683692 4804 683720
rect 2832 683680 2838 683692
rect 4798 683680 4804 683692
rect 4856 683680 4862 683732
rect 149054 683680 149060 683732
rect 149112 683720 149118 683732
rect 150434 683720 150440 683732
rect 149112 683692 150440 683720
rect 149112 683680 149118 683692
rect 150434 683680 150440 683692
rect 150492 683680 150498 683732
rect 372614 683612 372620 683664
rect 372672 683652 372678 683664
rect 375374 683652 375380 683664
rect 372672 683624 375380 683652
rect 372672 683612 372678 683624
rect 375374 683612 375380 683624
rect 375432 683612 375438 683664
rect 358078 681028 358084 681080
rect 358136 681068 358142 681080
rect 360470 681068 360476 681080
rect 358136 681040 360476 681068
rect 358136 681028 358142 681040
rect 360470 681028 360476 681040
rect 360528 681028 360534 681080
rect 261478 680960 261484 681012
rect 261536 681000 261542 681012
rect 282178 681000 282184 681012
rect 261536 680972 282184 681000
rect 261536 680960 261542 680972
rect 282178 680960 282184 680972
rect 282236 680960 282242 681012
rect 375374 680960 375380 681012
rect 375432 681000 375438 681012
rect 389174 681000 389180 681012
rect 375432 680972 389180 681000
rect 375432 680960 375438 680972
rect 389174 680960 389180 680972
rect 389232 680960 389238 681012
rect 360470 678240 360476 678292
rect 360528 678280 360534 678292
rect 369118 678280 369124 678292
rect 360528 678252 369124 678280
rect 360528 678240 360534 678252
rect 369118 678240 369124 678252
rect 369176 678240 369182 678292
rect 146202 676336 146208 676388
rect 146260 676376 146266 676388
rect 148962 676376 148968 676388
rect 146260 676348 148968 676376
rect 146260 676336 146266 676348
rect 148962 676336 148968 676348
rect 149020 676336 149026 676388
rect 369118 675452 369124 675504
rect 369176 675492 369182 675504
rect 378778 675492 378784 675504
rect 369176 675464 378784 675492
rect 369176 675452 369182 675464
rect 378778 675452 378784 675464
rect 378836 675452 378842 675504
rect 389174 675180 389180 675232
rect 389232 675220 389238 675232
rect 393314 675220 393320 675232
rect 389232 675192 393320 675220
rect 389232 675180 389238 675192
rect 393314 675180 393320 675192
rect 393372 675180 393378 675232
rect 143534 674432 143540 674484
rect 143592 674472 143598 674484
rect 146202 674472 146208 674484
rect 143592 674444 146208 674472
rect 143592 674432 143598 674444
rect 146202 674432 146208 674444
rect 146260 674432 146266 674484
rect 220814 673752 220820 673804
rect 220872 673792 220878 673804
rect 224218 673792 224224 673804
rect 220872 673764 224224 673792
rect 220872 673752 220878 673764
rect 224218 673752 224224 673764
rect 224276 673752 224282 673804
rect 393314 673208 393320 673260
rect 393372 673248 393378 673260
rect 396442 673248 396448 673260
rect 393372 673220 396448 673248
rect 393372 673208 393378 673220
rect 396442 673208 396448 673220
rect 396500 673208 396506 673260
rect 211522 672052 211528 672104
rect 211580 672092 211586 672104
rect 213178 672092 213184 672104
rect 211580 672064 213184 672092
rect 211580 672052 211586 672064
rect 213178 672052 213184 672064
rect 213236 672052 213242 672104
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 15838 670732 15844 670744
rect 3568 670704 15844 670732
rect 3568 670692 3574 670704
rect 15838 670692 15844 670704
rect 15896 670692 15902 670744
rect 208394 670692 208400 670744
rect 208452 670732 208458 670744
rect 211522 670732 211528 670744
rect 208452 670704 211528 670732
rect 208452 670692 208458 670704
rect 211522 670692 211528 670704
rect 211580 670692 211586 670744
rect 406378 670692 406384 670744
rect 406436 670732 406442 670744
rect 580166 670732 580172 670744
rect 406436 670704 580172 670732
rect 406436 670692 406442 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 143534 667944 143540 667956
rect 142126 667916 143540 667944
rect 140038 667836 140044 667888
rect 140096 667876 140102 667888
rect 142126 667876 142154 667916
rect 143534 667904 143540 667916
rect 143592 667904 143598 667956
rect 140096 667848 142154 667876
rect 140096 667836 140102 667848
rect 218698 667632 218704 667684
rect 218756 667672 218762 667684
rect 220814 667672 220820 667684
rect 218756 667644 220820 667672
rect 218756 667632 218762 667644
rect 220814 667632 220820 667644
rect 220872 667632 220878 667684
rect 261478 666584 261484 666596
rect 259472 666556 261484 666584
rect 258718 666476 258724 666528
rect 258776 666516 258782 666528
rect 259472 666516 259500 666556
rect 261478 666544 261484 666556
rect 261536 666544 261542 666596
rect 258776 666488 259500 666516
rect 258776 666476 258782 666488
rect 206278 665864 206284 665916
rect 206336 665904 206342 665916
rect 208302 665904 208308 665916
rect 206336 665876 208308 665904
rect 206336 665864 206342 665876
rect 208302 665864 208308 665876
rect 208360 665864 208366 665916
rect 378778 664436 378784 664488
rect 378836 664476 378842 664488
rect 387058 664476 387064 664488
rect 378836 664448 387064 664476
rect 378836 664436 378842 664448
rect 387058 664436 387064 664448
rect 387116 664436 387122 664488
rect 215294 662396 215300 662448
rect 215352 662436 215358 662448
rect 218698 662436 218704 662448
rect 215352 662408 218704 662436
rect 215352 662396 215358 662408
rect 218698 662396 218704 662408
rect 218756 662396 218762 662448
rect 323578 662328 323584 662380
rect 323636 662368 323642 662380
rect 326614 662368 326620 662380
rect 323636 662340 326620 662368
rect 323636 662328 323642 662340
rect 326614 662328 326620 662340
rect 326672 662328 326678 662380
rect 326614 659200 326620 659252
rect 326672 659240 326678 659252
rect 330018 659240 330024 659252
rect 326672 659212 330024 659240
rect 326672 659200 326678 659212
rect 330018 659200 330024 659212
rect 330076 659200 330082 659252
rect 211798 657568 211804 657620
rect 211856 657608 211862 657620
rect 215294 657608 215300 657620
rect 211856 657580 215300 657608
rect 211856 657568 211862 657580
rect 215294 657568 215300 657580
rect 215352 657568 215358 657620
rect 330018 656140 330024 656192
rect 330076 656180 330082 656192
rect 336734 656180 336740 656192
rect 330076 656152 336740 656180
rect 330076 656140 330082 656152
rect 336734 656140 336740 656152
rect 336792 656140 336798 656192
rect 257430 654100 257436 654152
rect 257488 654140 257494 654152
rect 258718 654140 258724 654152
rect 257488 654112 258724 654140
rect 257488 654100 257494 654112
rect 258718 654100 258724 654112
rect 258776 654100 258782 654152
rect 387058 652264 387064 652316
rect 387116 652304 387122 652316
rect 395338 652304 395344 652316
rect 387116 652276 395344 652304
rect 387116 652264 387122 652276
rect 395338 652264 395344 652276
rect 395396 652264 395402 652316
rect 138658 651380 138664 651432
rect 138716 651420 138722 651432
rect 140038 651420 140044 651432
rect 138716 651392 140044 651420
rect 138716 651380 138722 651392
rect 140038 651380 140044 651392
rect 140096 651380 140102 651432
rect 255314 651380 255320 651432
rect 255372 651420 255378 651432
rect 257430 651420 257436 651432
rect 255372 651392 257436 651420
rect 255372 651380 255378 651392
rect 257430 651380 257436 651392
rect 257488 651380 257494 651432
rect 336734 649272 336740 649324
rect 336792 649312 336798 649324
rect 345658 649312 345664 649324
rect 336792 649284 345664 649312
rect 336792 649272 336798 649284
rect 345658 649272 345664 649284
rect 345716 649272 345722 649324
rect 201402 647844 201408 647896
rect 201460 647884 201466 647896
rect 211798 647884 211804 647896
rect 201460 647856 211804 647884
rect 201460 647844 201466 647856
rect 211798 647844 211804 647856
rect 211856 647844 211862 647896
rect 204898 647164 204904 647216
rect 204956 647204 204962 647216
rect 206278 647204 206284 647216
rect 204956 647176 206284 647204
rect 204956 647164 204962 647176
rect 206278 647164 206284 647176
rect 206336 647164 206342 647216
rect 334618 646484 334624 646536
rect 334676 646524 334682 646536
rect 342898 646524 342904 646536
rect 334676 646496 342904 646524
rect 334676 646484 334682 646496
rect 342898 646484 342904 646496
rect 342956 646484 342962 646536
rect 189718 645124 189724 645176
rect 189776 645164 189782 645176
rect 201402 645164 201408 645176
rect 189776 645136 201408 645164
rect 189776 645124 189782 645136
rect 201402 645124 201408 645136
rect 201460 645124 201466 645176
rect 245562 645124 245568 645176
rect 245620 645164 245626 645176
rect 255314 645164 255320 645176
rect 245620 645136 255320 645164
rect 245620 645124 245626 645136
rect 255314 645124 255320 645136
rect 255372 645124 255378 645176
rect 345658 644308 345664 644360
rect 345716 644348 345722 644360
rect 353938 644348 353944 644360
rect 345716 644320 353944 644348
rect 345716 644308 345722 644320
rect 353938 644308 353944 644320
rect 353996 644308 354002 644360
rect 135898 641724 135904 641776
rect 135956 641764 135962 641776
rect 138658 641764 138664 641776
rect 135956 641736 138664 641764
rect 135956 641724 135962 641736
rect 138658 641724 138664 641736
rect 138716 641724 138722 641776
rect 243538 640296 243544 640348
rect 243596 640336 243602 640348
rect 245562 640336 245568 640348
rect 243596 640308 245568 640336
rect 243596 640296 243602 640308
rect 245562 640296 245568 640308
rect 245620 640296 245626 640348
rect 179414 636828 179420 636880
rect 179472 636868 179478 636880
rect 189718 636868 189724 636880
rect 179472 636840 189724 636868
rect 179472 636828 179478 636840
rect 189718 636828 189724 636840
rect 189776 636828 189782 636880
rect 2774 632068 2780 632120
rect 2832 632108 2838 632120
rect 4890 632108 4896 632120
rect 2832 632080 4896 632108
rect 2832 632068 2838 632080
rect 4890 632068 4896 632080
rect 4948 632068 4954 632120
rect 174446 630640 174452 630692
rect 174504 630680 174510 630692
rect 179414 630680 179420 630692
rect 174504 630652 179420 630680
rect 174504 630640 174510 630652
rect 179414 630640 179420 630652
rect 179472 630640 179478 630692
rect 171778 629008 171784 629060
rect 171836 629048 171842 629060
rect 174446 629048 174452 629060
rect 171836 629020 174452 629048
rect 171836 629008 171842 629020
rect 174446 629008 174452 629020
rect 174504 629008 174510 629060
rect 193858 623772 193864 623824
rect 193916 623812 193922 623824
rect 196618 623812 196624 623824
rect 193916 623784 196624 623812
rect 193916 623772 193922 623784
rect 196618 623772 196624 623784
rect 196676 623772 196682 623824
rect 243538 623812 243544 623824
rect 241532 623784 243544 623812
rect 239950 623704 239956 623756
rect 240008 623744 240014 623756
rect 241532 623744 241560 623784
rect 243538 623772 243544 623784
rect 243596 623772 243602 623824
rect 240008 623716 241560 623744
rect 240008 623704 240014 623716
rect 353938 622344 353944 622396
rect 353996 622384 354002 622396
rect 356698 622384 356704 622396
rect 353996 622356 356704 622384
rect 353996 622344 354002 622356
rect 356698 622344 356704 622356
rect 356756 622344 356762 622396
rect 237374 620984 237380 621036
rect 237432 621024 237438 621036
rect 239950 621024 239956 621036
rect 237432 620996 239956 621024
rect 237432 620984 237438 620996
rect 239950 620984 239956 620996
rect 240008 620984 240014 621036
rect 3510 618264 3516 618316
rect 3568 618304 3574 618316
rect 19978 618304 19984 618316
rect 3568 618276 19984 618304
rect 3568 618264 3574 618276
rect 19978 618264 19984 618276
rect 20036 618264 20042 618316
rect 237374 616876 237380 616888
rect 236012 616848 237380 616876
rect 233878 616768 233884 616820
rect 233936 616808 233942 616820
rect 236012 616808 236040 616848
rect 237374 616836 237380 616848
rect 237432 616836 237438 616888
rect 404998 616836 405004 616888
rect 405056 616876 405062 616888
rect 579706 616876 579712 616888
rect 405056 616848 579712 616876
rect 405056 616836 405062 616848
rect 579706 616836 579712 616848
rect 579764 616836 579770 616888
rect 233936 616780 236040 616808
rect 233936 616768 233942 616780
rect 342898 616088 342904 616140
rect 342956 616128 342962 616140
rect 360838 616128 360844 616140
rect 342956 616100 360844 616128
rect 342956 616088 342962 616100
rect 360838 616088 360844 616100
rect 360896 616088 360902 616140
rect 191098 610648 191104 610700
rect 191156 610688 191162 610700
rect 193858 610688 193864 610700
rect 191156 610660 193864 610688
rect 191156 610648 191162 610660
rect 193858 610648 193864 610660
rect 193916 610648 193922 610700
rect 232590 610240 232596 610292
rect 232648 610280 232654 610292
rect 234614 610280 234620 610292
rect 232648 610252 234620 610280
rect 232648 610240 232654 610252
rect 234614 610240 234620 610252
rect 234672 610240 234678 610292
rect 356698 607860 356704 607912
rect 356756 607900 356762 607912
rect 369118 607900 369124 607912
rect 356756 607872 369124 607900
rect 356756 607860 356762 607872
rect 369118 607860 369124 607872
rect 369176 607860 369182 607912
rect 153838 605072 153844 605124
rect 153896 605112 153902 605124
rect 171778 605112 171784 605124
rect 153896 605084 171784 605112
rect 153896 605072 153902 605084
rect 171778 605072 171784 605084
rect 171836 605072 171842 605124
rect 134518 603100 134524 603152
rect 134576 603140 134582 603152
rect 135898 603140 135904 603152
rect 134576 603112 135904 603140
rect 134576 603100 134582 603112
rect 135898 603100 135904 603112
rect 135956 603100 135962 603152
rect 232498 603100 232504 603152
rect 232556 603140 232562 603152
rect 233878 603140 233884 603152
rect 232556 603112 233884 603140
rect 232556 603100 232562 603112
rect 233878 603100 233884 603112
rect 233936 603100 233942 603152
rect 203610 601672 203616 601724
rect 203668 601712 203674 601724
rect 204898 601712 204904 601724
rect 203668 601684 204904 601712
rect 203668 601672 203674 601684
rect 204898 601672 204904 601684
rect 204956 601672 204962 601724
rect 224402 600924 224408 600976
rect 224460 600964 224466 600976
rect 232590 600964 232596 600976
rect 224460 600936 232596 600964
rect 224460 600924 224466 600936
rect 232590 600924 232596 600936
rect 232648 600924 232654 600976
rect 184198 599836 184204 599888
rect 184256 599876 184262 599888
rect 191098 599876 191104 599888
rect 184256 599848 191104 599876
rect 184256 599836 184262 599848
rect 191098 599836 191104 599848
rect 191156 599836 191162 599888
rect 202138 599632 202144 599684
rect 202196 599672 202202 599684
rect 203610 599672 203616 599684
rect 202196 599644 203616 599672
rect 202196 599632 202202 599644
rect 203610 599632 203616 599644
rect 203668 599632 203674 599684
rect 220814 598136 220820 598188
rect 220872 598176 220878 598188
rect 224402 598176 224408 598188
rect 220872 598148 224408 598176
rect 220872 598136 220878 598148
rect 224402 598136 224408 598148
rect 224460 598136 224466 598188
rect 214558 594804 214564 594856
rect 214616 594844 214622 594856
rect 220814 594844 220820 594856
rect 214616 594816 220820 594844
rect 214616 594804 214622 594816
rect 220814 594804 220820 594816
rect 220872 594804 220878 594856
rect 360838 594396 360844 594448
rect 360896 594436 360902 594448
rect 366358 594436 366364 594448
rect 360896 594408 366364 594436
rect 360896 594396 360902 594408
rect 366358 594396 366364 594408
rect 366416 594396 366422 594448
rect 181438 592016 181444 592068
rect 181496 592056 181502 592068
rect 184198 592056 184204 592068
rect 181496 592028 184204 592056
rect 181496 592016 181502 592028
rect 184198 592016 184204 592028
rect 184256 592016 184262 592068
rect 369118 590588 369124 590640
rect 369176 590628 369182 590640
rect 371878 590628 371884 590640
rect 369176 590600 371884 590628
rect 369176 590588 369182 590600
rect 371878 590588 371884 590600
rect 371936 590588 371942 590640
rect 371878 585760 371884 585812
rect 371936 585800 371942 585812
rect 380158 585800 380164 585812
rect 371936 585772 380164 585800
rect 371936 585760 371942 585772
rect 380158 585760 380164 585772
rect 380216 585760 380222 585812
rect 134518 583760 134524 583772
rect 132466 583732 134524 583760
rect 130378 583652 130384 583704
rect 130436 583692 130442 583704
rect 132466 583692 132494 583732
rect 134518 583720 134524 583732
rect 134576 583720 134582 583772
rect 130436 583664 132494 583692
rect 130436 583652 130442 583664
rect 3510 579640 3516 579692
rect 3568 579680 3574 579692
rect 10318 579680 10324 579692
rect 3568 579652 10324 579680
rect 3568 579640 3574 579652
rect 10318 579640 10324 579652
rect 10376 579640 10382 579692
rect 211798 578144 211804 578196
rect 211856 578184 211862 578196
rect 214558 578184 214564 578196
rect 211856 578156 214564 578184
rect 211856 578144 211862 578156
rect 214558 578144 214564 578156
rect 214616 578144 214622 578196
rect 149054 575220 149060 575272
rect 149112 575260 149118 575272
rect 153838 575260 153844 575272
rect 149112 575232 153844 575260
rect 149112 575220 149118 575232
rect 153838 575220 153844 575232
rect 153896 575220 153902 575272
rect 366358 574064 366364 574116
rect 366416 574104 366422 574116
rect 369118 574104 369124 574116
rect 366416 574076 369124 574104
rect 366416 574064 366422 574076
rect 369118 574064 369124 574076
rect 369176 574064 369182 574116
rect 231118 572704 231124 572756
rect 231176 572744 231182 572756
rect 232498 572744 232504 572756
rect 231176 572716 232504 572744
rect 231176 572704 231182 572716
rect 232498 572704 232504 572716
rect 232556 572704 232562 572756
rect 137278 571956 137284 572008
rect 137336 571996 137342 572008
rect 149054 571996 149060 572008
rect 137336 571968 149060 571996
rect 137336 571956 137342 571968
rect 149054 571956 149060 571968
rect 149112 571956 149118 572008
rect 380158 570596 380164 570648
rect 380216 570636 380222 570648
rect 392578 570636 392584 570648
rect 380216 570608 392584 570636
rect 380216 570596 380222 570608
rect 392578 570596 392584 570608
rect 392636 570596 392642 570648
rect 127618 567808 127624 567860
rect 127676 567848 127682 567860
rect 137278 567848 137284 567860
rect 127676 567820 137284 567848
rect 127676 567808 127682 567820
rect 137278 567808 137284 567820
rect 137336 567808 137342 567860
rect 3050 565836 3056 565888
rect 3108 565876 3114 565888
rect 37918 565876 37924 565888
rect 3108 565848 37924 565876
rect 3108 565836 3114 565848
rect 37918 565836 37924 565848
rect 37976 565836 37982 565888
rect 209038 564952 209044 565004
rect 209096 564992 209102 565004
rect 211798 564992 211804 565004
rect 209096 564964 211804 564992
rect 209096 564952 209102 564964
rect 211798 564952 211804 564964
rect 211856 564952 211862 565004
rect 229922 564680 229928 564732
rect 229980 564720 229986 564732
rect 231118 564720 231124 564732
rect 229980 564692 231124 564720
rect 229980 564680 229986 564692
rect 231118 564680 231124 564692
rect 231176 564680 231182 564732
rect 392578 564340 392584 564392
rect 392636 564380 392642 564392
rect 395430 564380 395436 564392
rect 392636 564352 395436 564380
rect 392636 564340 392642 564352
rect 395430 564340 395436 564352
rect 395488 564340 395494 564392
rect 403618 563048 403624 563100
rect 403676 563088 403682 563100
rect 580166 563088 580172 563100
rect 403676 563060 580172 563088
rect 403676 563048 403682 563060
rect 580166 563048 580172 563060
rect 580224 563048 580230 563100
rect 228358 562640 228364 562692
rect 228416 562680 228422 562692
rect 229922 562680 229928 562692
rect 228416 562652 229928 562680
rect 228416 562640 228422 562652
rect 229922 562640 229928 562652
rect 229980 562640 229986 562692
rect 189074 560940 189080 560992
rect 189132 560980 189138 560992
rect 202138 560980 202144 560992
rect 189132 560952 202144 560980
rect 189132 560940 189138 560952
rect 202138 560940 202144 560952
rect 202196 560940 202202 560992
rect 184934 558968 184940 559020
rect 184992 559008 184998 559020
rect 189074 559008 189080 559020
rect 184992 558980 189080 559008
rect 184992 558968 184998 558980
rect 189074 558968 189080 558980
rect 189132 558968 189138 559020
rect 124858 558832 124864 558884
rect 124916 558872 124922 558884
rect 127618 558872 127624 558884
rect 124916 558844 127624 558872
rect 124916 558832 124922 558844
rect 127618 558832 127624 558844
rect 127676 558832 127682 558884
rect 201218 556180 201224 556232
rect 201276 556220 201282 556232
rect 209038 556220 209044 556232
rect 201276 556192 209044 556220
rect 201276 556180 201282 556192
rect 209038 556180 209044 556192
rect 209096 556180 209102 556232
rect 163498 554004 163504 554056
rect 163556 554044 163562 554056
rect 181438 554044 181444 554056
rect 163556 554016 181444 554044
rect 163556 554004 163562 554016
rect 181438 554004 181444 554016
rect 181496 554004 181502 554056
rect 193858 552848 193864 552900
rect 193916 552888 193922 552900
rect 201218 552888 201224 552900
rect 193916 552860 201224 552888
rect 193916 552848 193922 552860
rect 201218 552848 201224 552860
rect 201276 552848 201282 552900
rect 183186 552644 183192 552696
rect 183244 552684 183250 552696
rect 184842 552684 184848 552696
rect 183244 552656 184848 552684
rect 183244 552644 183250 552656
rect 184842 552644 184848 552656
rect 184900 552644 184906 552696
rect 226978 552644 226984 552696
rect 227036 552684 227042 552696
rect 228358 552684 228364 552696
rect 227036 552656 228364 552684
rect 227036 552644 227042 552656
rect 228358 552644 228364 552656
rect 228416 552644 228422 552696
rect 181438 550400 181444 550452
rect 181496 550440 181502 550452
rect 183186 550440 183192 550452
rect 181496 550412 183192 550440
rect 181496 550400 181502 550412
rect 183186 550400 183192 550412
rect 183244 550400 183250 550452
rect 128998 550196 129004 550248
rect 129056 550236 129062 550248
rect 130378 550236 130384 550248
rect 129056 550208 130384 550236
rect 129056 550196 129062 550208
rect 130378 550196 130384 550208
rect 130436 550196 130442 550248
rect 146110 547136 146116 547188
rect 146168 547176 146174 547188
rect 163498 547176 163504 547188
rect 146168 547148 163504 547176
rect 146168 547136 146174 547148
rect 163498 547136 163504 547148
rect 163556 547136 163562 547188
rect 224954 546456 224960 546508
rect 225012 546496 225018 546508
rect 226978 546496 226984 546508
rect 225012 546468 226984 546496
rect 225012 546456 225018 546468
rect 226978 546456 226984 546468
rect 227036 546456 227042 546508
rect 170398 545708 170404 545760
rect 170456 545748 170462 545760
rect 193858 545748 193864 545760
rect 170456 545720 193864 545748
rect 170456 545708 170462 545720
rect 193858 545708 193864 545720
rect 193916 545708 193922 545760
rect 122098 545572 122104 545624
rect 122156 545612 122162 545624
rect 124858 545612 124864 545624
rect 122156 545584 124864 545612
rect 122156 545572 122162 545584
rect 124858 545572 124864 545584
rect 124916 545572 124922 545624
rect 133138 544348 133144 544400
rect 133196 544388 133202 544400
rect 146110 544388 146116 544400
rect 133196 544360 146116 544388
rect 133196 544348 133202 544360
rect 146110 544348 146116 544360
rect 146168 544348 146174 544400
rect 223022 540064 223028 540116
rect 223080 540104 223086 540116
rect 224862 540104 224868 540116
rect 223080 540076 224868 540104
rect 223080 540064 223086 540076
rect 224862 540064 224868 540076
rect 224920 540064 224926 540116
rect 156598 537480 156604 537532
rect 156656 537520 156662 537532
rect 170398 537520 170404 537532
rect 156656 537492 170404 537520
rect 156656 537480 156662 537492
rect 170398 537480 170404 537492
rect 170456 537480 170462 537532
rect 123478 536052 123484 536104
rect 123536 536092 123542 536104
rect 133138 536092 133144 536104
rect 123536 536064 133144 536092
rect 123536 536052 123542 536064
rect 133138 536052 133144 536064
rect 133196 536052 133202 536104
rect 220354 535440 220360 535492
rect 220412 535480 220418 535492
rect 223022 535480 223028 535492
rect 220412 535452 223028 535480
rect 220412 535440 220418 535452
rect 223022 535440 223028 535452
rect 223080 535440 223086 535492
rect 180058 534012 180064 534064
rect 180116 534052 180122 534064
rect 181438 534052 181444 534064
rect 180116 534024 181444 534052
rect 180116 534012 180122 534024
rect 181438 534012 181444 534024
rect 181496 534012 181502 534064
rect 218698 532312 218704 532364
rect 218756 532352 218762 532364
rect 220354 532352 220360 532364
rect 218756 532324 220360 532352
rect 218756 532312 218762 532324
rect 220354 532312 220360 532324
rect 220412 532312 220418 532364
rect 117130 527144 117136 527196
rect 117188 527184 117194 527196
rect 122098 527184 122104 527196
rect 117188 527156 122104 527184
rect 117188 527144 117194 527156
rect 122098 527144 122104 527156
rect 122156 527144 122162 527196
rect 106918 525036 106924 525088
rect 106976 525076 106982 525088
rect 128998 525076 129004 525088
rect 106976 525048 129004 525076
rect 106976 525036 106982 525048
rect 128998 525036 129004 525048
rect 129056 525036 129062 525088
rect 101398 519528 101404 519580
rect 101456 519568 101462 519580
rect 117130 519568 117136 519580
rect 101456 519540 117136 519568
rect 101456 519528 101462 519540
rect 117130 519528 117136 519540
rect 117188 519528 117194 519580
rect 127618 516740 127624 516792
rect 127676 516780 127682 516792
rect 156598 516780 156604 516792
rect 127676 516752 156604 516780
rect 127676 516740 127682 516752
rect 156598 516740 156604 516752
rect 156656 516740 156662 516792
rect 3326 514768 3332 514820
rect 3384 514808 3390 514820
rect 43438 514808 43444 514820
rect 3384 514780 43444 514808
rect 3384 514768 3390 514780
rect 43438 514768 43444 514780
rect 43496 514768 43502 514820
rect 105538 514020 105544 514072
rect 105596 514060 105602 514072
rect 106918 514060 106924 514072
rect 105596 514032 106924 514060
rect 105596 514020 105602 514032
rect 106918 514020 106924 514032
rect 106976 514020 106982 514072
rect 98638 511912 98644 511964
rect 98696 511952 98702 511964
rect 101398 511952 101404 511964
rect 98696 511924 101404 511952
rect 98696 511912 98702 511924
rect 101398 511912 101404 511924
rect 101456 511912 101462 511964
rect 400858 510620 400864 510672
rect 400916 510660 400922 510672
rect 580166 510660 580172 510672
rect 400916 510632 580172 510660
rect 400916 510620 400922 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 113818 508512 113824 508564
rect 113876 508552 113882 508564
rect 123478 508552 123484 508564
rect 113876 508524 123484 508552
rect 113876 508512 113882 508524
rect 123478 508512 123484 508524
rect 123536 508512 123542 508564
rect 178678 505112 178684 505164
rect 178736 505152 178742 505164
rect 180058 505152 180064 505164
rect 178736 505124 180064 505152
rect 178736 505112 178742 505124
rect 180058 505112 180064 505124
rect 180116 505112 180122 505164
rect 102778 499536 102784 499588
rect 102836 499576 102842 499588
rect 105538 499576 105544 499588
rect 102836 499548 105544 499576
rect 102836 499536 102842 499548
rect 105538 499536 105544 499548
rect 105596 499536 105602 499588
rect 175274 498176 175280 498228
rect 175332 498216 175338 498228
rect 178678 498216 178684 498228
rect 175332 498188 178684 498216
rect 175332 498176 175338 498188
rect 178678 498176 178684 498188
rect 178736 498176 178742 498228
rect 173158 493280 173164 493332
rect 173216 493320 173222 493332
rect 175182 493320 175188 493332
rect 173216 493292 175188 493320
rect 173216 493280 173222 493292
rect 175182 493280 175188 493292
rect 175240 493280 175246 493332
rect 217318 493280 217324 493332
rect 217376 493320 217382 493332
rect 218698 493320 218704 493332
rect 217376 493292 218704 493320
rect 217376 493280 217382 493292
rect 218698 493280 218704 493292
rect 218756 493280 218762 493332
rect 369118 490356 369124 490408
rect 369176 490396 369182 490408
rect 376018 490396 376024 490408
rect 369176 490368 376024 490396
rect 369176 490356 369182 490368
rect 376018 490356 376024 490368
rect 376076 490356 376082 490408
rect 171134 482808 171140 482860
rect 171192 482848 171198 482860
rect 173158 482848 173164 482860
rect 171192 482820 173164 482848
rect 171192 482808 171198 482820
rect 173158 482808 173164 482820
rect 173216 482808 173222 482860
rect 215938 482672 215944 482724
rect 215996 482712 216002 482724
rect 217318 482712 217324 482724
rect 215996 482684 217324 482712
rect 215996 482672 216002 482684
rect 217318 482672 217324 482684
rect 217376 482672 217382 482724
rect 119338 482264 119344 482316
rect 119396 482304 119402 482316
rect 127618 482304 127624 482316
rect 119396 482276 127624 482304
rect 119396 482264 119402 482276
rect 127618 482264 127624 482276
rect 127676 482264 127682 482316
rect 171134 478904 171140 478916
rect 171106 478864 171140 478904
rect 171192 478864 171198 478916
rect 167638 478796 167644 478848
rect 167696 478836 167702 478848
rect 171106 478836 171134 478864
rect 167696 478808 171134 478836
rect 167696 478796 167702 478808
rect 101398 477504 101404 477556
rect 101456 477544 101462 477556
rect 102778 477544 102784 477556
rect 101456 477516 102784 477544
rect 101456 477504 101462 477516
rect 102778 477504 102784 477516
rect 102836 477504 102842 477556
rect 116578 469208 116584 469260
rect 116636 469248 116642 469260
rect 119338 469248 119344 469260
rect 116636 469220 119344 469248
rect 116636 469208 116642 469220
rect 119338 469208 119344 469220
rect 119396 469208 119402 469260
rect 213178 469208 213184 469260
rect 213236 469248 213242 469260
rect 215938 469248 215944 469260
rect 213236 469220 215944 469248
rect 213236 469208 213242 469220
rect 215938 469208 215944 469220
rect 215996 469208 216002 469260
rect 95878 466420 95884 466472
rect 95936 466460 95942 466472
rect 98638 466460 98644 466472
rect 95936 466432 98644 466460
rect 95936 466420 95942 466432
rect 98638 466420 98644 466432
rect 98696 466420 98702 466472
rect 2774 462544 2780 462596
rect 2832 462584 2838 462596
rect 4982 462584 4988 462596
rect 2832 462556 4988 462584
rect 2832 462544 2838 462556
rect 4982 462544 4988 462556
rect 5040 462544 5046 462596
rect 399478 456764 399484 456816
rect 399536 456804 399542 456816
rect 580166 456804 580172 456816
rect 399536 456776 580172 456804
rect 399536 456764 399542 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 376018 456016 376024 456068
rect 376076 456056 376082 456068
rect 385678 456056 385684 456068
rect 376076 456028 385684 456056
rect 376076 456016 376082 456028
rect 385678 456016 385684 456028
rect 385736 456016 385742 456068
rect 213178 454084 213184 454096
rect 211172 454056 213184 454084
rect 210510 453976 210516 454028
rect 210568 454016 210574 454028
rect 211172 454016 211200 454056
rect 213178 454044 213184 454056
rect 213236 454044 213242 454096
rect 210568 453988 211200 454016
rect 210568 453976 210574 453988
rect 101398 452656 101404 452668
rect 99392 452628 101404 452656
rect 97258 452548 97264 452600
rect 97316 452588 97322 452600
rect 99392 452588 99420 452628
rect 101398 452616 101404 452628
rect 101456 452616 101462 452668
rect 97316 452560 99420 452588
rect 97316 452548 97322 452560
rect 108298 447720 108304 447772
rect 108356 447760 108362 447772
rect 113818 447760 113824 447772
rect 108356 447732 113824 447760
rect 108356 447720 108362 447732
rect 113818 447720 113824 447732
rect 113876 447720 113882 447772
rect 209038 446360 209044 446412
rect 209096 446400 209102 446412
rect 210510 446400 210516 446412
rect 209096 446372 210516 446400
rect 209096 446360 209102 446372
rect 210510 446360 210516 446372
rect 210568 446360 210574 446412
rect 207658 438880 207664 438932
rect 207716 438920 207722 438932
rect 209038 438920 209044 438932
rect 207716 438892 209044 438920
rect 207716 438880 207722 438892
rect 209038 438880 209044 438892
rect 209096 438880 209102 438932
rect 204898 430584 204904 430636
rect 204956 430624 204962 430636
rect 207658 430624 207664 430636
rect 204956 430596 207664 430624
rect 204956 430584 204962 430596
rect 207658 430584 207664 430596
rect 207716 430584 207722 430636
rect 396718 430584 396724 430636
rect 396776 430624 396782 430636
rect 579982 430624 579988 430636
rect 396776 430596 579988 430624
rect 396776 430584 396782 430596
rect 579982 430584 579988 430596
rect 580040 430584 580046 430636
rect 93118 429700 93124 429752
rect 93176 429740 93182 429752
rect 95878 429740 95884 429752
rect 93176 429712 95884 429740
rect 93176 429700 93182 429712
rect 95878 429700 95884 429712
rect 95936 429700 95942 429752
rect 100018 424328 100024 424380
rect 100076 424368 100082 424380
rect 108298 424368 108304 424380
rect 100076 424340 108304 424368
rect 100076 424328 100082 424340
rect 108298 424328 108304 424340
rect 108356 424328 108362 424380
rect 166258 423580 166264 423632
rect 166316 423620 166322 423632
rect 167638 423620 167644 423632
rect 166316 423592 167644 423620
rect 166316 423580 166322 423592
rect 167638 423580 167644 423592
rect 167696 423580 167702 423632
rect 3142 422900 3148 422952
rect 3200 422940 3206 422952
rect 6178 422940 6184 422952
rect 3200 422912 6184 422940
rect 3200 422900 3206 422912
rect 6178 422900 6184 422912
rect 6236 422900 6242 422952
rect 398098 418140 398104 418192
rect 398156 418180 398162 418192
rect 580166 418180 580172 418192
rect 398156 418152 580172 418180
rect 398156 418140 398162 418152
rect 580166 418140 580172 418152
rect 580224 418140 580230 418192
rect 164786 415080 164792 415132
rect 164844 415120 164850 415132
rect 166258 415120 166264 415132
rect 164844 415092 166264 415120
rect 164844 415080 164850 415092
rect 166258 415080 166264 415092
rect 166316 415080 166322 415132
rect 95878 415012 95884 415064
rect 95936 415052 95942 415064
rect 97258 415052 97264 415064
rect 95936 415024 97264 415052
rect 95936 415012 95942 415024
rect 97258 415012 97264 415024
rect 97316 415012 97322 415064
rect 108298 411884 108304 411936
rect 108356 411924 108362 411936
rect 116578 411924 116584 411936
rect 108356 411896 116584 411924
rect 108356 411884 108362 411896
rect 116578 411884 116584 411896
rect 116636 411884 116642 411936
rect 3326 409912 3332 409964
rect 3384 409952 3390 409964
rect 8938 409952 8944 409964
rect 3384 409924 8944 409952
rect 3384 409912 3390 409924
rect 8938 409912 8944 409924
rect 8996 409912 9002 409964
rect 161842 407124 161848 407176
rect 161900 407164 161906 407176
rect 164786 407164 164792 407176
rect 161900 407136 164792 407164
rect 161900 407124 161906 407136
rect 164786 407124 164792 407136
rect 164844 407124 164850 407176
rect 93210 406376 93216 406428
rect 93268 406416 93274 406428
rect 100018 406416 100024 406428
rect 93268 406388 100024 406416
rect 93268 406376 93274 406388
rect 100018 406376 100024 406388
rect 100076 406376 100082 406428
rect 160094 406376 160100 406428
rect 160152 406416 160158 406428
rect 161842 406416 161848 406428
rect 160152 406388 161848 406416
rect 160152 406376 160158 406388
rect 161842 406376 161848 406388
rect 161900 406376 161906 406428
rect 160094 404376 160100 404388
rect 158732 404348 160100 404376
rect 157334 404268 157340 404320
rect 157392 404308 157398 404320
rect 158732 404308 158760 404348
rect 160094 404336 160100 404348
rect 160152 404336 160158 404388
rect 421558 404336 421564 404388
rect 421616 404376 421622 404388
rect 580166 404376 580172 404388
rect 421616 404348 580172 404376
rect 421616 404336 421622 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 157392 404280 158760 404308
rect 157392 404268 157398 404280
rect 157334 400228 157340 400240
rect 155972 400200 157340 400228
rect 153838 400120 153844 400172
rect 153896 400160 153902 400172
rect 155972 400160 156000 400200
rect 157334 400188 157340 400200
rect 157392 400188 157398 400240
rect 153896 400132 156000 400160
rect 153896 400120 153902 400132
rect 69658 396720 69664 396772
rect 69716 396760 69722 396772
rect 136634 396760 136640 396772
rect 69716 396732 136640 396760
rect 69716 396720 69722 396732
rect 136634 396720 136640 396732
rect 136692 396720 136698 396772
rect 105538 394612 105544 394664
rect 105596 394652 105602 394664
rect 108298 394652 108304 394664
rect 105596 394624 108304 394652
rect 105596 394612 105602 394624
rect 108298 394612 108304 394624
rect 108356 394612 108362 394664
rect 93302 393320 93308 393372
rect 93360 393360 93366 393372
rect 95878 393360 95884 393372
rect 93360 393332 95884 393360
rect 93360 393320 93366 393332
rect 95878 393320 95884 393332
rect 95936 393320 95942 393372
rect 153838 392000 153844 392012
rect 151786 391972 153844 392000
rect 146938 391892 146944 391944
rect 146996 391932 147002 391944
rect 151786 391932 151814 391972
rect 153838 391960 153844 391972
rect 153896 391960 153902 392012
rect 146996 391904 151814 391932
rect 146996 391892 147002 391904
rect 385678 388492 385684 388544
rect 385736 388532 385742 388544
rect 389266 388532 389272 388544
rect 385736 388504 389272 388532
rect 385736 388492 385742 388504
rect 389266 388492 389272 388504
rect 389324 388492 389330 388544
rect 199378 388424 199384 388476
rect 199436 388464 199442 388476
rect 204898 388464 204904 388476
rect 199436 388436 204904 388464
rect 199436 388424 199442 388436
rect 204898 388424 204904 388436
rect 204956 388424 204962 388476
rect 97534 385024 97540 385076
rect 97592 385064 97598 385076
rect 105538 385064 105544 385076
rect 97592 385036 105544 385064
rect 97592 385024 97598 385036
rect 105538 385024 105544 385036
rect 105596 385024 105602 385076
rect 68278 384956 68284 385008
rect 68336 384996 68342 385008
rect 69658 384996 69664 385008
rect 68336 384968 69664 384996
rect 68336 384956 68342 384968
rect 69658 384956 69664 384968
rect 69716 384956 69722 385008
rect 389266 384956 389272 385008
rect 389324 384996 389330 385008
rect 392762 384996 392768 385008
rect 389324 384968 392768 384996
rect 389324 384956 389330 384968
rect 392762 384956 392768 384968
rect 392820 384956 392826 385008
rect 88978 384412 88984 384464
rect 89036 384452 89042 384464
rect 93210 384452 93216 384464
rect 89036 384424 93216 384452
rect 89036 384412 89042 384424
rect 93210 384412 93216 384424
rect 93268 384412 93274 384464
rect 86862 382916 86868 382968
rect 86920 382956 86926 382968
rect 97534 382956 97540 382968
rect 86920 382928 97540 382956
rect 86920 382916 86926 382928
rect 97534 382916 97540 382928
rect 97592 382916 97598 382968
rect 392762 382168 392768 382220
rect 392820 382208 392826 382220
rect 395522 382208 395528 382220
rect 392820 382180 395528 382208
rect 392820 382168 392826 382180
rect 395522 382168 395528 382180
rect 395580 382168 395586 382220
rect 91922 379516 91928 379568
rect 91980 379556 91986 379568
rect 93302 379556 93308 379568
rect 91980 379528 93308 379556
rect 91980 379516 91986 379528
rect 93302 379516 93308 379528
rect 93360 379516 93366 379568
rect 79318 379040 79324 379092
rect 79376 379080 79382 379092
rect 86862 379080 86868 379092
rect 79376 379052 86868 379080
rect 79376 379040 79382 379052
rect 86862 379040 86868 379052
rect 86920 379040 86926 379092
rect 396902 378156 396908 378208
rect 396960 378196 396966 378208
rect 579798 378196 579804 378208
rect 396960 378168 579804 378196
rect 396960 378156 396966 378168
rect 579798 378156 579804 378168
rect 579856 378156 579862 378208
rect 90358 377816 90364 377868
rect 90416 377856 90422 377868
rect 91922 377856 91928 377868
rect 90416 377828 91928 377856
rect 90416 377816 90422 377828
rect 91922 377816 91928 377828
rect 91980 377816 91986 377868
rect 197354 372580 197360 372632
rect 197412 372620 197418 372632
rect 199378 372620 199384 372632
rect 197412 372592 199384 372620
rect 197412 372580 197418 372592
rect 199378 372580 199384 372592
rect 199436 372580 199442 372632
rect 3326 371220 3332 371272
rect 3384 371260 3390 371272
rect 10410 371260 10416 371272
rect 3384 371232 10416 371260
rect 3384 371220 3390 371232
rect 10410 371220 10416 371232
rect 10468 371220 10474 371272
rect 197354 369900 197360 369912
rect 193232 369872 197360 369900
rect 192478 369792 192484 369844
rect 192536 369832 192542 369844
rect 193232 369832 193260 369872
rect 197354 369860 197360 369872
rect 197412 369860 197418 369912
rect 192536 369804 193260 369832
rect 192536 369792 192542 369804
rect 87506 364488 87512 364540
rect 87564 364528 87570 364540
rect 90358 364528 90364 364540
rect 87564 364500 90364 364528
rect 87564 364488 87570 364500
rect 90358 364488 90364 364500
rect 90416 364488 90422 364540
rect 73798 359456 73804 359508
rect 73856 359496 73862 359508
rect 88978 359496 88984 359508
rect 73856 359468 88984 359496
rect 73856 359456 73862 359468
rect 88978 359456 88984 359468
rect 89036 359456 89042 359508
rect 65702 359048 65708 359100
rect 65760 359088 65766 359100
rect 68278 359088 68284 359100
rect 65760 359060 68284 359088
rect 65760 359048 65766 359060
rect 68278 359048 68284 359060
rect 68336 359048 68342 359100
rect 86218 358912 86224 358964
rect 86276 358952 86282 358964
rect 87506 358952 87512 358964
rect 86276 358924 87512 358952
rect 86276 358912 86282 358924
rect 87506 358912 87512 358924
rect 87564 358912 87570 358964
rect 146938 358816 146944 358828
rect 144932 358788 146944 358816
rect 142798 358708 142804 358760
rect 142856 358748 142862 358760
rect 144932 358748 144960 358788
rect 146938 358776 146944 358788
rect 146996 358776 147002 358828
rect 142856 358720 144960 358748
rect 142856 358708 142862 358720
rect 64138 358164 64144 358216
rect 64196 358204 64202 358216
rect 65702 358204 65708 358216
rect 64196 358176 65708 358204
rect 64196 358164 64202 358176
rect 65702 358164 65708 358176
rect 65760 358164 65766 358216
rect 54478 358028 54484 358080
rect 54536 358068 54542 358080
rect 79318 358068 79324 358080
rect 54536 358040 79324 358068
rect 54536 358028 54542 358040
rect 79318 358028 79324 358040
rect 79376 358028 79382 358080
rect 3326 357416 3332 357468
rect 3384 357456 3390 357468
rect 24118 357456 24124 357468
rect 3384 357428 24124 357456
rect 3384 357416 3390 357428
rect 24118 357416 24124 357428
rect 24176 357416 24182 357468
rect 85022 353268 85028 353320
rect 85080 353308 85086 353320
rect 86218 353308 86224 353320
rect 85080 353280 86224 353308
rect 85080 353268 85086 353280
rect 86218 353268 86224 353280
rect 86276 353268 86282 353320
rect 140774 353268 140780 353320
rect 140832 353308 140838 353320
rect 142798 353308 142804 353320
rect 140832 353280 142804 353308
rect 140832 353268 140838 353280
rect 142798 353268 142804 353280
rect 142856 353268 142862 353320
rect 418798 351908 418804 351960
rect 418856 351948 418862 351960
rect 580074 351948 580080 351960
rect 418856 351920 580080 351948
rect 418856 351908 418862 351920
rect 580074 351908 580080 351920
rect 580132 351908 580138 351960
rect 82814 351296 82820 351348
rect 82872 351336 82878 351348
rect 85022 351336 85028 351348
rect 82872 351308 85028 351336
rect 82872 351296 82878 351308
rect 85022 351296 85028 351308
rect 85080 351296 85086 351348
rect 137278 350548 137284 350600
rect 137336 350588 137342 350600
rect 140774 350588 140780 350600
rect 137336 350560 140780 350588
rect 137336 350548 137342 350560
rect 140774 350548 140780 350560
rect 140832 350548 140838 350600
rect 51718 349460 51724 349512
rect 51776 349500 51782 349512
rect 54478 349500 54484 349512
rect 51776 349472 54484 349500
rect 51776 349460 51782 349472
rect 54478 349460 54484 349472
rect 54536 349460 54542 349512
rect 82814 346440 82820 346452
rect 80072 346412 82820 346440
rect 78674 346332 78680 346384
rect 78732 346372 78738 346384
rect 80072 346372 80100 346412
rect 82814 346400 82820 346412
rect 82872 346400 82878 346452
rect 78732 346344 80100 346372
rect 78732 346332 78738 346344
rect 2774 345176 2780 345228
rect 2832 345216 2838 345228
rect 5074 345216 5080 345228
rect 2832 345188 5080 345216
rect 2832 345176 2838 345188
rect 5074 345176 5080 345188
rect 5132 345176 5138 345228
rect 189718 345040 189724 345092
rect 189776 345080 189782 345092
rect 192478 345080 192484 345092
rect 189776 345052 192484 345080
rect 189776 345040 189782 345052
rect 192478 345040 192484 345052
rect 192536 345040 192542 345092
rect 395522 343612 395528 343664
rect 395580 343652 395586 343664
rect 397546 343652 397552 343664
rect 395580 343624 397552 343652
rect 395580 343612 395586 343624
rect 397546 343612 397552 343624
rect 397604 343612 397610 343664
rect 75914 340892 75920 340944
rect 75972 340932 75978 340944
rect 78582 340932 78588 340944
rect 75972 340904 78588 340932
rect 75972 340892 75978 340904
rect 78582 340892 78588 340904
rect 78640 340892 78646 340944
rect 62114 340144 62120 340196
rect 62172 340184 62178 340196
rect 73798 340184 73804 340196
rect 62172 340156 73804 340184
rect 62172 340144 62178 340156
rect 73798 340144 73804 340156
rect 73856 340144 73862 340196
rect 53834 337356 53840 337408
rect 53892 337396 53898 337408
rect 62114 337396 62120 337408
rect 53892 337368 62120 337396
rect 53892 337356 53898 337368
rect 62114 337356 62120 337368
rect 62172 337356 62178 337408
rect 73154 336744 73160 336796
rect 73212 336784 73218 336796
rect 75822 336784 75828 336796
rect 73212 336756 75828 336784
rect 73212 336744 73218 336756
rect 75822 336744 75828 336756
rect 75880 336744 75886 336796
rect 189718 336784 189724 336796
rect 186332 336756 189724 336784
rect 186222 336676 186228 336728
rect 186280 336716 186286 336728
rect 186332 336716 186360 336756
rect 189718 336744 189724 336756
rect 189776 336744 189782 336796
rect 186280 336688 186360 336716
rect 186280 336676 186286 336688
rect 46382 333956 46388 334008
rect 46440 333996 46446 334008
rect 53834 333996 53840 334008
rect 46440 333968 53840 333996
rect 46440 333956 46446 333968
rect 53834 333956 53840 333968
rect 53892 333956 53898 334008
rect 73062 332636 73068 332648
rect 70412 332608 73068 332636
rect 70302 332528 70308 332580
rect 70360 332568 70366 332580
rect 70412 332568 70440 332608
rect 73062 332596 73068 332608
rect 73120 332596 73126 332648
rect 70360 332540 70440 332568
rect 70360 332528 70366 332540
rect 62850 331848 62856 331900
rect 62908 331888 62914 331900
rect 88334 331888 88340 331900
rect 62908 331860 88340 331888
rect 62908 331848 62914 331860
rect 88334 331848 88340 331860
rect 88392 331848 88398 331900
rect 44910 331508 44916 331560
rect 44968 331548 44974 331560
rect 46382 331548 46388 331560
rect 44968 331520 46388 331548
rect 44968 331508 44974 331520
rect 46382 331508 46388 331520
rect 46440 331508 46446 331560
rect 45002 330488 45008 330540
rect 45060 330528 45066 330540
rect 51718 330528 51724 330540
rect 45060 330500 51724 330528
rect 45060 330488 45066 330500
rect 51718 330488 51724 330500
rect 51776 330488 51782 330540
rect 183554 330012 183560 330064
rect 183612 330052 183618 330064
rect 186222 330052 186228 330064
rect 183612 330024 186228 330052
rect 183612 330012 183618 330024
rect 186222 330012 186228 330024
rect 186280 330012 186286 330064
rect 134518 329536 134524 329588
rect 134576 329576 134582 329588
rect 137278 329576 137284 329588
rect 134576 329548 137284 329576
rect 134576 329536 134582 329548
rect 137278 329536 137284 329548
rect 137336 329536 137342 329588
rect 68186 328040 68192 328092
rect 68244 328080 68250 328092
rect 70302 328080 70308 328092
rect 68244 328052 70308 328080
rect 68244 328040 68250 328052
rect 70302 328040 70308 328052
rect 70360 328040 70366 328092
rect 182818 326408 182824 326460
rect 182876 326448 182882 326460
rect 183554 326448 183560 326460
rect 182876 326420 183560 326448
rect 182876 326408 182882 326420
rect 183554 326408 183560 326420
rect 183612 326408 183618 326460
rect 397086 324300 397092 324352
rect 397144 324340 397150 324352
rect 580074 324340 580080 324352
rect 397144 324312 580080 324340
rect 397144 324300 397150 324312
rect 580074 324300 580080 324312
rect 580132 324300 580138 324352
rect 134518 320192 134524 320204
rect 132466 320164 134524 320192
rect 66898 320084 66904 320136
rect 66956 320124 66962 320136
rect 68186 320124 68192 320136
rect 66956 320096 68192 320124
rect 66956 320084 66962 320096
rect 68186 320084 68192 320096
rect 68244 320084 68250 320136
rect 126238 320084 126244 320136
rect 126296 320124 126302 320136
rect 132466 320124 132494 320164
rect 134518 320152 134524 320164
rect 134576 320152 134582 320204
rect 126296 320096 132494 320124
rect 126296 320084 126302 320096
rect 62758 319404 62764 319456
rect 62816 319444 62822 319456
rect 64138 319444 64144 319456
rect 62816 319416 64144 319444
rect 62816 319404 62822 319416
rect 64138 319404 64144 319416
rect 64196 319404 64202 319456
rect 3142 318792 3148 318844
rect 3200 318832 3206 318844
rect 33778 318832 33784 318844
rect 3200 318804 33784 318832
rect 3200 318792 3206 318804
rect 33778 318792 33784 318804
rect 33836 318792 33842 318844
rect 61470 318384 61476 318436
rect 61528 318424 61534 318436
rect 62850 318424 62856 318436
rect 61528 318396 62856 318424
rect 61528 318384 61534 318396
rect 62850 318384 62856 318396
rect 62908 318384 62914 318436
rect 84838 315256 84844 315308
rect 84896 315296 84902 315308
rect 104894 315296 104900 315308
rect 84896 315268 104900 315296
rect 84896 315256 84902 315268
rect 104894 315256 104900 315268
rect 104952 315256 104958 315308
rect 62114 312128 62120 312180
rect 62172 312168 62178 312180
rect 66898 312168 66904 312180
rect 62172 312140 66904 312168
rect 62172 312128 62178 312140
rect 66898 312128 66904 312140
rect 66956 312128 66962 312180
rect 90358 311856 90364 311908
rect 90416 311896 90422 311908
rect 93118 311896 93124 311908
rect 90416 311868 93124 311896
rect 90416 311856 90422 311868
rect 93118 311856 93124 311868
rect 93176 311856 93182 311908
rect 398190 311856 398196 311908
rect 398248 311896 398254 311908
rect 580074 311896 580080 311908
rect 398248 311868 580080 311896
rect 398248 311856 398254 311868
rect 580074 311856 580080 311868
rect 580132 311856 580138 311908
rect 59998 311176 60004 311228
rect 60056 311216 60062 311228
rect 61470 311216 61476 311228
rect 60056 311188 61476 311216
rect 60056 311176 60062 311188
rect 61470 311176 61476 311188
rect 61528 311176 61534 311228
rect 60090 307232 60096 307284
rect 60148 307272 60154 307284
rect 62114 307272 62120 307284
rect 60148 307244 62120 307272
rect 60148 307232 60154 307244
rect 62114 307232 62120 307244
rect 62172 307232 62178 307284
rect 179598 306348 179604 306400
rect 179656 306388 179662 306400
rect 182818 306388 182824 306400
rect 179656 306360 182824 306388
rect 179656 306348 179662 306360
rect 182818 306348 182824 306360
rect 182876 306348 182882 306400
rect 178678 301384 178684 301436
rect 178736 301424 178742 301436
rect 179598 301424 179604 301436
rect 178736 301396 179604 301424
rect 178736 301384 178742 301396
rect 179598 301384 179604 301396
rect 179656 301384 179662 301436
rect 61562 299072 61568 299124
rect 61620 299112 61626 299124
rect 62758 299112 62764 299124
rect 61620 299084 62764 299112
rect 61620 299072 61626 299084
rect 62758 299072 62764 299084
rect 62816 299072 62822 299124
rect 417418 298120 417424 298172
rect 417476 298160 417482 298172
rect 580074 298160 580080 298172
rect 417476 298132 580080 298160
rect 417476 298120 417482 298132
rect 580074 298120 580080 298132
rect 580132 298120 580138 298172
rect 73154 294584 73160 294636
rect 73212 294624 73218 294636
rect 90358 294624 90364 294636
rect 73212 294596 90364 294624
rect 73212 294584 73218 294596
rect 90358 294584 90364 294596
rect 90416 294584 90422 294636
rect 60182 293972 60188 294024
rect 60240 294012 60246 294024
rect 61562 294012 61568 294024
rect 60240 293984 61568 294012
rect 60240 293972 60246 293984
rect 61562 293972 61568 293984
rect 61620 293972 61626 294024
rect 175274 293972 175280 294024
rect 175332 294012 175338 294024
rect 178678 294012 178684 294024
rect 175332 293984 178684 294012
rect 175332 293972 175338 293984
rect 178678 293972 178684 293984
rect 178736 293972 178742 294024
rect 124858 292544 124864 292596
rect 124916 292584 124922 292596
rect 126238 292584 126244 292596
rect 124916 292556 126244 292584
rect 124916 292544 124922 292556
rect 126238 292544 126244 292556
rect 126296 292544 126302 292596
rect 66990 291184 66996 291236
rect 67048 291224 67054 291236
rect 73154 291224 73160 291236
rect 67048 291196 73160 291224
rect 67048 291184 67054 291196
rect 73154 291184 73160 291196
rect 73212 291184 73218 291236
rect 58618 291116 58624 291168
rect 58676 291156 58682 291168
rect 59998 291156 60004 291168
rect 58676 291128 60004 291156
rect 58676 291116 58682 291128
rect 59998 291116 60004 291128
rect 60056 291116 60062 291168
rect 60090 289864 60096 289876
rect 57992 289836 60096 289864
rect 55214 289756 55220 289808
rect 55272 289796 55278 289808
rect 57992 289796 58020 289836
rect 60090 289824 60096 289836
rect 60148 289824 60154 289876
rect 55272 289768 58020 289796
rect 55272 289756 55278 289768
rect 55858 289076 55864 289128
rect 55916 289116 55922 289128
rect 66990 289116 66996 289128
rect 55916 289088 66996 289116
rect 55916 289076 55922 289088
rect 66990 289076 66996 289088
rect 67048 289076 67054 289128
rect 57238 287648 57244 287700
rect 57296 287688 57302 287700
rect 71774 287688 71780 287700
rect 57296 287660 71780 287688
rect 57296 287648 57302 287660
rect 71774 287648 71780 287660
rect 71832 287648 71838 287700
rect 58618 284356 58624 284368
rect 56612 284328 58624 284356
rect 56502 284248 56508 284300
rect 56560 284288 56566 284300
rect 56612 284288 56640 284328
rect 58618 284316 58624 284328
rect 58676 284316 58682 284368
rect 84838 284356 84844 284368
rect 84166 284328 84844 284356
rect 56560 284260 56640 284288
rect 56560 284248 56566 284260
rect 82078 284248 82084 284300
rect 82136 284288 82142 284300
rect 84166 284288 84194 284328
rect 84838 284316 84844 284328
rect 84896 284316 84902 284368
rect 82136 284260 84194 284288
rect 82136 284248 82142 284260
rect 57974 282888 57980 282940
rect 58032 282928 58038 282940
rect 60182 282928 60188 282940
rect 58032 282900 60188 282928
rect 58032 282888 58038 282900
rect 60182 282888 60188 282900
rect 60240 282888 60246 282940
rect 173158 281800 173164 281852
rect 173216 281840 173222 281852
rect 174906 281840 174912 281852
rect 173216 281812 174912 281840
rect 173216 281800 173222 281812
rect 174906 281800 174912 281812
rect 174964 281800 174970 281852
rect 54202 281392 54208 281444
rect 54260 281432 54266 281444
rect 56502 281432 56508 281444
rect 54260 281404 56508 281432
rect 54260 281392 54266 281404
rect 56502 281392 56508 281404
rect 56560 281392 56566 281444
rect 53282 280780 53288 280832
rect 53340 280820 53346 280832
rect 169754 280820 169760 280832
rect 53340 280792 169760 280820
rect 53340 280780 53346 280792
rect 169754 280780 169760 280792
rect 169812 280780 169818 280832
rect 53374 280168 53380 280220
rect 53432 280208 53438 280220
rect 55122 280208 55128 280220
rect 53432 280180 55128 280208
rect 53432 280168 53438 280180
rect 55122 280168 55128 280180
rect 55180 280168 55186 280220
rect 53098 279420 53104 279472
rect 53156 279460 53162 279472
rect 54202 279460 54208 279472
rect 53156 279432 54208 279460
rect 53156 279420 53162 279432
rect 54202 279420 54208 279432
rect 54260 279420 54266 279472
rect 54478 278740 54484 278792
rect 54536 278780 54542 278792
rect 57882 278780 57888 278792
rect 54536 278752 57888 278780
rect 54536 278740 54542 278752
rect 57882 278740 57888 278752
rect 57940 278740 57946 278792
rect 57238 277420 57244 277432
rect 55232 277392 57244 277420
rect 53834 277312 53840 277364
rect 53892 277352 53898 277364
rect 55232 277352 55260 277392
rect 57238 277380 57244 277392
rect 57296 277380 57302 277432
rect 53892 277324 55260 277352
rect 53892 277312 53898 277324
rect 55950 276632 55956 276684
rect 56008 276672 56014 276684
rect 82078 276672 82084 276684
rect 56008 276644 82084 276672
rect 56008 276632 56014 276644
rect 82078 276632 82084 276644
rect 82136 276632 82142 276684
rect 50338 274864 50344 274916
rect 50396 274904 50402 274916
rect 55858 274904 55864 274916
rect 50396 274876 55864 274904
rect 50396 274864 50402 274876
rect 55858 274864 55864 274876
rect 55916 274864 55922 274916
rect 50430 274728 50436 274780
rect 50488 274768 50494 274780
rect 53374 274768 53380 274780
rect 50488 274740 53380 274768
rect 50488 274728 50494 274740
rect 53374 274728 53380 274740
rect 53432 274728 53438 274780
rect 53190 274660 53196 274712
rect 53248 274700 53254 274712
rect 53834 274700 53840 274712
rect 53248 274672 53840 274700
rect 53248 274660 53254 274672
rect 53834 274660 53840 274672
rect 53892 274660 53898 274712
rect 124858 273272 124864 273284
rect 122806 273244 124864 273272
rect 118694 273164 118700 273216
rect 118752 273204 118758 273216
rect 122806 273204 122834 273244
rect 124858 273232 124864 273244
rect 124916 273232 124922 273284
rect 118752 273176 122834 273204
rect 118752 273164 118758 273176
rect 51718 272008 51724 272060
rect 51776 272048 51782 272060
rect 53098 272048 53104 272060
rect 51776 272020 53104 272048
rect 51776 272008 51782 272020
rect 53098 272008 53104 272020
rect 53156 272008 53162 272060
rect 396810 271872 396816 271924
rect 396868 271912 396874 271924
rect 579798 271912 579804 271924
rect 396868 271884 579804 271912
rect 396868 271872 396874 271884
rect 579798 271872 579804 271884
rect 579856 271872 579862 271924
rect 167638 271804 167644 271856
rect 167696 271844 167702 271856
rect 173158 271844 173164 271856
rect 167696 271816 173164 271844
rect 167696 271804 167702 271816
rect 173158 271804 173164 271816
rect 173216 271804 173222 271856
rect 116762 270512 116768 270564
rect 116820 270552 116826 270564
rect 118694 270552 118700 270564
rect 116820 270524 118700 270552
rect 116820 270512 116826 270524
rect 118694 270512 118700 270524
rect 118752 270512 118758 270564
rect 51074 270444 51080 270496
rect 51132 270484 51138 270496
rect 53282 270484 53288 270496
rect 51132 270456 53288 270484
rect 51132 270444 51138 270456
rect 53282 270444 53288 270456
rect 53340 270444 53346 270496
rect 45278 268336 45284 268388
rect 45336 268376 45342 268388
rect 50338 268376 50344 268388
rect 45336 268348 50344 268376
rect 45336 268336 45342 268348
rect 50338 268336 50344 268348
rect 50396 268336 50402 268388
rect 112162 268336 112168 268388
rect 112220 268376 112226 268388
rect 116762 268376 116768 268388
rect 112220 268348 116768 268376
rect 112220 268336 112226 268348
rect 116762 268336 116768 268348
rect 116820 268336 116826 268388
rect 3142 266704 3148 266756
rect 3200 266744 3206 266756
rect 9030 266744 9036 266756
rect 3200 266716 9036 266744
rect 3200 266704 3206 266716
rect 9030 266704 9036 266716
rect 9088 266704 9094 266756
rect 165614 266568 165620 266620
rect 165672 266608 165678 266620
rect 167638 266608 167644 266620
rect 165672 266580 167644 266608
rect 165672 266568 165678 266580
rect 167638 266568 167644 266580
rect 167696 266568 167702 266620
rect 53190 266432 53196 266484
rect 53248 266472 53254 266484
rect 54478 266472 54484 266484
rect 53248 266444 54484 266472
rect 53248 266432 53254 266444
rect 54478 266432 54484 266444
rect 54536 266432 54542 266484
rect 50430 266404 50436 266416
rect 46952 266376 50436 266404
rect 46198 266296 46204 266348
rect 46256 266336 46262 266348
rect 46952 266336 46980 266376
rect 50430 266364 50436 266376
rect 50488 266364 50494 266416
rect 51074 266404 51080 266416
rect 50540 266376 51080 266404
rect 46256 266308 46980 266336
rect 46256 266296 46262 266308
rect 48314 266296 48320 266348
rect 48372 266336 48378 266348
rect 50540 266336 50568 266376
rect 51074 266364 51080 266376
rect 51132 266364 51138 266416
rect 54202 266364 54208 266416
rect 54260 266404 54266 266416
rect 55950 266404 55956 266416
rect 54260 266376 55956 266404
rect 54260 266364 54266 266376
rect 55950 266364 55956 266376
rect 56008 266364 56014 266416
rect 109034 266364 109040 266416
rect 109092 266404 109098 266416
rect 112162 266404 112168 266416
rect 109092 266376 112168 266404
rect 109092 266364 109098 266376
rect 112162 266364 112168 266376
rect 112220 266364 112226 266416
rect 48372 266308 50568 266336
rect 48372 266296 48378 266308
rect 158714 265616 158720 265668
rect 158772 265656 158778 265668
rect 165614 265656 165620 265668
rect 158772 265628 165620 265656
rect 158772 265616 158778 265628
rect 165614 265616 165620 265628
rect 165672 265616 165678 265668
rect 49694 263576 49700 263628
rect 49752 263616 49758 263628
rect 51718 263616 51724 263628
rect 49752 263588 51724 263616
rect 49752 263576 49758 263588
rect 51718 263576 51724 263588
rect 51776 263576 51782 263628
rect 53282 263576 53288 263628
rect 53340 263616 53346 263628
rect 54202 263616 54208 263628
rect 53340 263588 54208 263616
rect 53340 263576 53346 263588
rect 54202 263576 54208 263588
rect 54260 263576 54266 263628
rect 107010 260448 107016 260500
rect 107068 260488 107074 260500
rect 108942 260488 108948 260500
rect 107068 260460 108948 260488
rect 107068 260448 107074 260460
rect 108942 260448 108948 260460
rect 109000 260448 109006 260500
rect 151814 259224 151820 259276
rect 151872 259264 151878 259276
rect 158714 259264 158720 259276
rect 151872 259236 158720 259264
rect 151872 259224 151878 259236
rect 158714 259224 158720 259236
rect 158772 259224 158778 259276
rect 45738 259088 45744 259140
rect 45796 259128 45802 259140
rect 48222 259128 48228 259140
rect 45796 259100 48228 259128
rect 45796 259088 45802 259100
rect 48222 259088 48228 259100
rect 48280 259088 48286 259140
rect 46934 258544 46940 258596
rect 46992 258584 46998 258596
rect 49694 258584 49700 258596
rect 46992 258556 49700 258584
rect 46992 258544 46998 258556
rect 49694 258544 49700 258556
rect 49752 258544 49758 258596
rect 418890 258068 418896 258120
rect 418948 258108 418954 258120
rect 579982 258108 579988 258120
rect 418948 258080 579988 258108
rect 418948 258068 418954 258080
rect 579982 258068 579988 258080
rect 580040 258068 580046 258120
rect 45186 256708 45192 256760
rect 45244 256748 45250 256760
rect 46198 256748 46204 256760
rect 45244 256720 46204 256748
rect 45244 256708 45250 256720
rect 46198 256708 46204 256720
rect 46256 256708 46262 256760
rect 53282 256748 53288 256760
rect 51092 256720 53288 256748
rect 50430 256640 50436 256692
rect 50488 256680 50494 256692
rect 51092 256680 51120 256720
rect 53282 256708 53288 256720
rect 53340 256708 53346 256760
rect 104894 256708 104900 256760
rect 104952 256748 104958 256760
rect 107010 256748 107016 256760
rect 104952 256720 107016 256748
rect 104952 256708 104958 256720
rect 107010 256708 107016 256720
rect 107068 256708 107074 256760
rect 50488 256652 51120 256680
rect 50488 256640 50494 256652
rect 45646 255280 45652 255332
rect 45704 255320 45710 255332
rect 46934 255320 46940 255332
rect 45704 255292 46940 255320
rect 45704 255280 45710 255292
rect 46934 255280 46940 255292
rect 46992 255280 46998 255332
rect 104894 255320 104900 255332
rect 103486 255292 104900 255320
rect 101398 255212 101404 255264
rect 101456 255252 101462 255264
rect 103486 255252 103514 255292
rect 104894 255280 104900 255292
rect 104952 255280 104958 255332
rect 101456 255224 103514 255252
rect 101456 255212 101462 255224
rect 53190 254028 53196 254040
rect 46952 254000 53196 254028
rect 3142 253920 3148 253972
rect 3200 253960 3206 253972
rect 22738 253960 22744 253972
rect 3200 253932 22744 253960
rect 3200 253920 3206 253932
rect 22738 253920 22744 253932
rect 22796 253920 22802 253972
rect 46198 253852 46204 253904
rect 46256 253892 46262 253904
rect 46952 253892 46980 254000
rect 53190 253988 53196 254000
rect 53248 253988 53254 254040
rect 47578 253920 47584 253972
rect 47636 253960 47642 253972
rect 50430 253960 50436 253972
rect 47636 253932 50436 253960
rect 47636 253920 47642 253932
rect 50430 253920 50436 253932
rect 50488 253920 50494 253972
rect 151722 253960 151728 253972
rect 147692 253932 151728 253960
rect 46256 253864 46980 253892
rect 46256 253852 46262 253864
rect 146938 253852 146944 253904
rect 146996 253892 147002 253904
rect 147692 253892 147720 253932
rect 151722 253920 151728 253932
rect 151780 253920 151786 253972
rect 146996 253864 147720 253892
rect 146996 253852 147002 253864
rect 51074 252832 51080 252884
rect 51132 252872 51138 252884
rect 53098 252872 53104 252884
rect 51132 252844 53104 252872
rect 51132 252832 51138 252844
rect 53098 252832 53104 252844
rect 53156 252832 53162 252884
rect 50338 250384 50344 250436
rect 50396 250424 50402 250436
rect 51074 250424 51080 250436
rect 50396 250396 51080 250424
rect 50396 250384 50402 250396
rect 51074 250384 51080 250396
rect 51132 250384 51138 250436
rect 143258 247052 143264 247104
rect 143316 247092 143322 247104
rect 146938 247092 146944 247104
rect 143316 247064 146944 247092
rect 143316 247052 143322 247064
rect 146938 247052 146944 247064
rect 146996 247052 147002 247104
rect 45830 245624 45836 245676
rect 45888 245664 45894 245676
rect 47578 245664 47584 245676
rect 45888 245636 47584 245664
rect 45888 245624 45894 245636
rect 47578 245624 47584 245636
rect 47636 245624 47642 245676
rect 44818 244944 44824 244996
rect 44876 244984 44882 244996
rect 46198 244984 46204 244996
rect 44876 244956 46204 244984
rect 44876 244944 44882 244956
rect 46198 244944 46204 244956
rect 46256 244944 46262 244996
rect 414658 244264 414664 244316
rect 414716 244304 414722 244316
rect 579982 244304 579988 244316
rect 414716 244276 579988 244304
rect 414716 244264 414722 244276
rect 579982 244264 579988 244276
rect 580040 244264 580046 244316
rect 45094 240796 45100 240848
rect 45152 240836 45158 240848
rect 101398 240836 101404 240848
rect 45152 240808 101404 240836
rect 45152 240796 45158 240808
rect 101398 240796 101404 240808
rect 101456 240796 101462 240848
rect 45462 240728 45468 240780
rect 45520 240768 45526 240780
rect 143258 240768 143264 240780
rect 45520 240740 143264 240768
rect 45520 240728 45526 240740
rect 143258 240728 143264 240740
rect 143316 240728 143322 240780
rect 45646 240524 45652 240576
rect 45704 240564 45710 240576
rect 50338 240564 50344 240576
rect 45704 240536 50344 240564
rect 45704 240524 45710 240536
rect 50338 240524 50344 240536
rect 50396 240524 50402 240576
rect 2774 240184 2780 240236
rect 2832 240224 2838 240236
rect 5166 240224 5172 240236
rect 2832 240196 5172 240224
rect 2832 240184 2838 240196
rect 5166 240184 5172 240196
rect 5224 240184 5230 240236
rect 395430 240048 395436 240100
rect 395488 240088 395494 240100
rect 396534 240088 396540 240100
rect 395488 240060 396540 240088
rect 395488 240048 395494 240060
rect 396534 240048 396540 240060
rect 396592 240048 396598 240100
rect 395338 239776 395344 239828
rect 395396 239816 395402 239828
rect 395396 239788 395936 239816
rect 395396 239776 395402 239788
rect 45370 238756 45376 238808
rect 45428 238796 45434 238808
rect 45830 238796 45836 238808
rect 45428 238768 45836 238796
rect 45428 238756 45434 238768
rect 45830 238756 45836 238768
rect 45888 238756 45894 238808
rect 395908 238660 395936 239788
rect 396534 238796 396540 238808
rect 396046 238768 396540 238796
rect 396046 238728 396074 238768
rect 396534 238756 396540 238768
rect 396592 238756 396598 238808
rect 396626 238728 396632 238740
rect 396046 238700 396632 238728
rect 396626 238688 396632 238700
rect 396684 238688 396690 238740
rect 396534 238660 396540 238672
rect 395908 238632 396540 238660
rect 396534 238620 396540 238632
rect 396592 238620 396598 238672
rect 45738 233316 45744 233368
rect 45796 233356 45802 233368
rect 45796 233328 46060 233356
rect 45796 233316 45802 233328
rect 45554 233248 45560 233300
rect 45612 233288 45618 233300
rect 45612 233260 45968 233288
rect 45612 233248 45618 233260
rect 45370 233180 45376 233232
rect 45428 233220 45434 233232
rect 45428 233192 45692 233220
rect 45428 233180 45434 233192
rect 45094 233112 45100 233164
rect 45152 233152 45158 233164
rect 45664 233152 45692 233192
rect 45830 233152 45836 233164
rect 45152 233124 45554 233152
rect 45664 233124 45836 233152
rect 45152 233112 45158 233124
rect 45526 232892 45554 233124
rect 45830 233112 45836 233124
rect 45888 233112 45894 233164
rect 45940 233016 45968 233260
rect 46032 233084 46060 233328
rect 46032 233056 64874 233084
rect 45940 232988 58940 233016
rect 45526 232852 45560 232892
rect 45554 232840 45560 232852
rect 45612 232840 45618 232892
rect 45462 232772 45468 232824
rect 45520 232812 45526 232824
rect 45738 232812 45744 232824
rect 45520 232784 45744 232812
rect 45520 232772 45526 232784
rect 45738 232772 45744 232784
rect 45796 232772 45802 232824
rect 58912 232812 58940 232988
rect 58912 232784 62804 232812
rect 62776 232416 62804 232784
rect 62758 232364 62764 232416
rect 62816 232364 62822 232416
rect 64846 232404 64874 233056
rect 82078 232404 82084 232416
rect 64846 232376 82084 232404
rect 82078 232364 82084 232376
rect 82136 232364 82142 232416
rect 395430 232364 395436 232416
rect 395488 232404 395494 232416
rect 396626 232404 396632 232416
rect 395488 232376 396632 232404
rect 395488 232364 395494 232376
rect 396626 232364 396632 232376
rect 396684 232364 396690 232416
rect 395338 232296 395344 232348
rect 395396 232336 395402 232348
rect 396442 232336 396448 232348
rect 395396 232308 396448 232336
rect 395396 232296 395402 232308
rect 396442 232296 396448 232308
rect 396500 232296 396506 232348
rect 391198 232228 391204 232280
rect 391256 232268 391262 232280
rect 396534 232268 396540 232280
rect 391256 232240 396540 232268
rect 391256 232228 391262 232240
rect 396534 232228 396540 232240
rect 396592 232228 396598 232280
rect 393958 231820 393964 231872
rect 394016 231860 394022 231872
rect 580074 231860 580080 231872
rect 394016 231832 580080 231860
rect 394016 231820 394022 231832
rect 580074 231820 580080 231832
rect 580132 231820 580138 231872
rect 45830 231140 45836 231192
rect 45888 231180 45894 231192
rect 134150 231180 134156 231192
rect 45888 231152 134156 231180
rect 45888 231140 45894 231152
rect 134150 231140 134156 231152
rect 134208 231140 134214 231192
rect 4062 231072 4068 231124
rect 4120 231112 4126 231124
rect 180794 231112 180800 231124
rect 4120 231084 180800 231112
rect 4120 231072 4126 231084
rect 180794 231072 180800 231084
rect 180852 231072 180858 231124
rect 44818 231004 44824 231056
rect 44876 231044 44882 231056
rect 84838 231044 84844 231056
rect 44876 231016 84844 231044
rect 44876 231004 44882 231016
rect 84838 231004 84844 231016
rect 84896 231004 84902 231056
rect 44910 230528 44916 230580
rect 44968 230568 44974 230580
rect 47670 230568 47676 230580
rect 44968 230540 47676 230568
rect 44968 230528 44974 230540
rect 47670 230528 47676 230540
rect 47728 230528 47734 230580
rect 45738 230392 45744 230444
rect 45796 230432 45802 230444
rect 47578 230432 47584 230444
rect 45796 230404 47584 230432
rect 45796 230392 45802 230404
rect 47578 230392 47584 230404
rect 47636 230392 47642 230444
rect 45554 230324 45560 230376
rect 45612 230364 45618 230376
rect 55122 230364 55128 230376
rect 45612 230336 55128 230364
rect 45612 230324 45618 230336
rect 55122 230324 55128 230336
rect 55180 230324 55186 230376
rect 134150 230052 134156 230104
rect 134208 230092 134214 230104
rect 136358 230092 136364 230104
rect 134208 230064 136364 230092
rect 134208 230052 134214 230064
rect 136358 230052 136364 230064
rect 136416 230052 136422 230104
rect 3878 229712 3884 229764
rect 3936 229752 3942 229764
rect 179414 229752 179420 229764
rect 3936 229724 179420 229752
rect 3936 229712 3942 229724
rect 179414 229712 179420 229724
rect 179472 229712 179478 229764
rect 45002 228352 45008 228404
rect 45060 228392 45066 228404
rect 49970 228392 49976 228404
rect 45060 228364 49976 228392
rect 45060 228352 45066 228364
rect 49970 228352 49976 228364
rect 50028 228352 50034 228404
rect 157978 228352 157984 228404
rect 158036 228392 158042 228404
rect 266538 228392 266544 228404
rect 158036 228364 266544 228392
rect 158036 228352 158042 228364
rect 266538 228352 266544 228364
rect 266596 228352 266602 228404
rect 266998 228352 267004 228404
rect 267056 228392 267062 228404
rect 356514 228392 356520 228404
rect 267056 228364 356520 228392
rect 267056 228352 267062 228364
rect 356514 228352 356520 228364
rect 356572 228352 356578 228404
rect 3142 227740 3148 227792
rect 3200 227780 3206 227792
rect 138658 227780 138664 227792
rect 3200 227752 138664 227780
rect 3200 227740 3206 227752
rect 138658 227740 138664 227752
rect 138716 227740 138722 227792
rect 388438 227740 388444 227792
rect 388496 227780 388502 227792
rect 391198 227780 391204 227792
rect 388496 227752 391204 227780
rect 388496 227740 388502 227752
rect 391198 227740 391204 227752
rect 391256 227740 391262 227792
rect 391290 227740 391296 227792
rect 391348 227780 391354 227792
rect 395430 227780 395436 227792
rect 391348 227752 395436 227780
rect 391348 227740 391354 227752
rect 395430 227740 395436 227752
rect 395488 227740 395494 227792
rect 82078 227672 82084 227724
rect 82136 227712 82142 227724
rect 85482 227712 85488 227724
rect 82136 227684 85488 227712
rect 82136 227672 82142 227684
rect 85482 227672 85488 227684
rect 85540 227672 85546 227724
rect 62758 227128 62764 227180
rect 62816 227168 62822 227180
rect 65794 227168 65800 227180
rect 62816 227140 65800 227168
rect 62816 227128 62822 227140
rect 65794 227128 65800 227140
rect 65852 227128 65858 227180
rect 45186 226244 45192 226296
rect 45244 226284 45250 226296
rect 48222 226284 48228 226296
rect 45244 226256 48228 226284
rect 45244 226244 45250 226256
rect 48222 226244 48228 226256
rect 48280 226244 48286 226296
rect 136358 225156 136364 225208
rect 136416 225196 136422 225208
rect 138750 225196 138756 225208
rect 136416 225168 138756 225196
rect 136416 225156 136422 225168
rect 138750 225156 138756 225168
rect 138808 225156 138814 225208
rect 49970 224952 49976 225004
rect 50028 224992 50034 225004
rect 53834 224992 53840 225004
rect 50028 224964 53840 224992
rect 50028 224952 50034 224964
rect 53834 224952 53840 224964
rect 53892 224952 53898 225004
rect 389082 224952 389088 225004
rect 389140 224992 389146 225004
rect 391290 224992 391296 225004
rect 389140 224964 391296 224992
rect 389140 224952 389146 224964
rect 391290 224952 391296 224964
rect 391348 224952 391354 225004
rect 85482 224204 85488 224256
rect 85540 224244 85546 224256
rect 100018 224244 100024 224256
rect 85540 224216 100024 224244
rect 85540 224204 85546 224216
rect 100018 224204 100024 224216
rect 100076 224204 100082 224256
rect 55214 224136 55220 224188
rect 55272 224176 55278 224188
rect 59354 224176 59360 224188
rect 55272 224148 59360 224176
rect 55272 224136 55278 224148
rect 59354 224136 59360 224148
rect 59412 224136 59418 224188
rect 394050 223524 394056 223576
rect 394108 223564 394114 223576
rect 395338 223564 395344 223576
rect 394108 223536 395344 223564
rect 394108 223524 394114 223536
rect 395338 223524 395344 223536
rect 395396 223524 395402 223576
rect 118694 222844 118700 222896
rect 118752 222884 118758 222896
rect 580166 222884 580172 222896
rect 118752 222856 580172 222884
rect 118752 222844 118758 222856
rect 580166 222844 580172 222856
rect 580224 222844 580230 222896
rect 48222 222164 48228 222216
rect 48280 222204 48286 222216
rect 48280 222176 51120 222204
rect 48280 222164 48286 222176
rect 47578 222096 47584 222148
rect 47636 222136 47642 222148
rect 48314 222136 48320 222148
rect 47636 222108 48320 222136
rect 47636 222096 47642 222108
rect 48314 222096 48320 222108
rect 48372 222096 48378 222148
rect 51092 222136 51120 222176
rect 53190 222136 53196 222148
rect 51092 222108 53196 222136
rect 53190 222096 53196 222108
rect 53248 222096 53254 222148
rect 65794 222096 65800 222148
rect 65852 222136 65858 222148
rect 69658 222136 69664 222148
rect 65852 222108 69664 222136
rect 65852 222096 65858 222108
rect 69658 222096 69664 222108
rect 69716 222096 69722 222148
rect 53834 221416 53840 221468
rect 53892 221456 53898 221468
rect 59262 221456 59268 221468
rect 53892 221428 59268 221456
rect 53892 221416 53898 221428
rect 59262 221416 59268 221428
rect 59320 221416 59326 221468
rect 59354 220736 59360 220788
rect 59412 220776 59418 220788
rect 62758 220776 62764 220788
rect 59412 220748 62764 220776
rect 59412 220736 59418 220748
rect 62758 220736 62764 220748
rect 62816 220736 62822 220788
rect 84838 220736 84844 220788
rect 84896 220776 84902 220788
rect 85758 220776 85764 220788
rect 84896 220748 85764 220776
rect 84896 220736 84902 220748
rect 85758 220736 85764 220748
rect 85816 220736 85822 220788
rect 385034 220736 385040 220788
rect 385092 220776 385098 220788
rect 389082 220776 389088 220788
rect 385092 220748 389088 220776
rect 385092 220736 385098 220748
rect 389082 220736 389088 220748
rect 389140 220736 389146 220788
rect 48314 219444 48320 219496
rect 48372 219484 48378 219496
rect 48372 219456 52500 219484
rect 48372 219444 48378 219456
rect 52472 219416 52500 219456
rect 55122 219416 55128 219428
rect 52472 219388 55128 219416
rect 55122 219376 55128 219388
rect 55180 219376 55186 219428
rect 138750 218696 138756 218748
rect 138808 218736 138814 218748
rect 158714 218736 158720 218748
rect 138808 218708 158720 218736
rect 138808 218696 138814 218708
rect 158714 218696 158720 218708
rect 158772 218696 158778 218748
rect 394418 218084 394424 218136
rect 394476 218124 394482 218136
rect 397546 218124 397552 218136
rect 394476 218096 397552 218124
rect 394476 218084 394482 218096
rect 397546 218084 397552 218096
rect 397604 218084 397610 218136
rect 85758 218016 85764 218068
rect 85816 218056 85822 218068
rect 87598 218056 87604 218068
rect 85816 218028 87604 218056
rect 85816 218016 85822 218028
rect 87598 218016 87604 218028
rect 87656 218016 87662 218068
rect 118602 218016 118608 218068
rect 118660 218056 118666 218068
rect 579982 218056 579988 218068
rect 118660 218028 579988 218056
rect 118660 218016 118666 218028
rect 579982 218016 579988 218028
rect 580040 218016 580046 218068
rect 380894 217880 380900 217932
rect 380952 217920 380958 217932
rect 385034 217920 385040 217932
rect 380952 217892 385040 217920
rect 380952 217880 380958 217892
rect 385034 217880 385040 217892
rect 385092 217880 385098 217932
rect 45278 217608 45284 217660
rect 45336 217648 45342 217660
rect 47578 217648 47584 217660
rect 45336 217620 47584 217648
rect 45336 217608 45342 217620
rect 47578 217608 47584 217620
rect 47636 217608 47642 217660
rect 47670 216724 47676 216776
rect 47728 216764 47734 216776
rect 50338 216764 50344 216776
rect 47728 216736 50344 216764
rect 47728 216724 47734 216736
rect 50338 216724 50344 216736
rect 50396 216724 50402 216776
rect 158714 215976 158720 216028
rect 158772 216016 158778 216028
rect 162762 216016 162768 216028
rect 158772 215988 162768 216016
rect 158772 215976 158778 215988
rect 162762 215976 162768 215988
rect 162820 215976 162826 216028
rect 100018 215908 100024 215960
rect 100076 215948 100082 215960
rect 111058 215948 111064 215960
rect 100076 215920 111064 215948
rect 100076 215908 100082 215920
rect 111058 215908 111064 215920
rect 111116 215908 111122 215960
rect 59262 215704 59268 215756
rect 59320 215744 59326 215756
rect 61378 215744 61384 215756
rect 59320 215716 61384 215744
rect 59320 215704 59326 215716
rect 61378 215704 61384 215716
rect 61436 215704 61442 215756
rect 375466 215432 375472 215484
rect 375524 215472 375530 215484
rect 380894 215472 380900 215484
rect 375524 215444 380900 215472
rect 375524 215432 375530 215444
rect 380894 215432 380900 215444
rect 380952 215432 380958 215484
rect 53190 215228 53196 215280
rect 53248 215268 53254 215280
rect 53834 215268 53840 215280
rect 53248 215240 53840 215268
rect 53248 215228 53254 215240
rect 53834 215228 53840 215240
rect 53892 215228 53898 215280
rect 3142 213936 3148 213988
rect 3200 213976 3206 213988
rect 179506 213976 179512 213988
rect 3200 213948 179512 213976
rect 3200 213936 3206 213948
rect 179506 213936 179512 213948
rect 179564 213936 179570 213988
rect 375466 213976 375472 213988
rect 373966 213948 375472 213976
rect 371878 213868 371884 213920
rect 371936 213908 371942 213920
rect 373966 213908 373994 213948
rect 375466 213936 375472 213948
rect 375524 213936 375530 213988
rect 371936 213880 373994 213908
rect 371936 213868 371942 213880
rect 55214 213188 55220 213240
rect 55272 213228 55278 213240
rect 68278 213228 68284 213240
rect 55272 213200 68284 213228
rect 55272 213188 55278 213200
rect 68278 213188 68284 213200
rect 68336 213188 68342 213240
rect 391198 213120 391204 213172
rect 391256 213160 391262 213172
rect 394418 213160 394424 213172
rect 391256 213132 394424 213160
rect 391256 213120 391262 213132
rect 394418 213120 394424 213132
rect 394476 213120 394482 213172
rect 162762 212848 162768 212900
rect 162820 212888 162826 212900
rect 164878 212888 164884 212900
rect 162820 212860 164884 212888
rect 162820 212848 162826 212860
rect 164878 212848 164884 212860
rect 164936 212848 164942 212900
rect 53834 211692 53840 211744
rect 53892 211732 53898 211744
rect 55214 211732 55220 211744
rect 53892 211704 55220 211732
rect 53892 211692 53898 211704
rect 55214 211692 55220 211704
rect 55272 211692 55278 211744
rect 69658 209516 69664 209568
rect 69716 209556 69722 209568
rect 77018 209556 77024 209568
rect 69716 209528 77024 209556
rect 69716 209516 69722 209528
rect 77018 209516 77024 209528
rect 77076 209516 77082 209568
rect 55214 208836 55220 208888
rect 55272 208876 55278 208888
rect 56870 208876 56876 208888
rect 55272 208848 56876 208876
rect 55272 208836 55278 208848
rect 56870 208836 56876 208848
rect 56928 208836 56934 208888
rect 164878 208360 164884 208412
rect 164936 208400 164942 208412
rect 166258 208400 166264 208412
rect 164936 208372 166264 208400
rect 164936 208360 164942 208372
rect 166258 208360 166264 208372
rect 166316 208360 166322 208412
rect 45554 207612 45560 207664
rect 45612 207652 45618 207664
rect 50430 207652 50436 207664
rect 45612 207624 50436 207652
rect 45612 207612 45618 207624
rect 50430 207612 50436 207624
rect 50488 207612 50494 207664
rect 77018 205776 77024 205828
rect 77076 205816 77082 205828
rect 78674 205816 78680 205828
rect 77076 205788 78680 205816
rect 77076 205776 77082 205788
rect 78674 205776 78680 205788
rect 78732 205776 78738 205828
rect 50338 205708 50344 205760
rect 50396 205748 50402 205760
rect 54478 205748 54484 205760
rect 50396 205720 54484 205748
rect 50396 205708 50402 205720
rect 54478 205708 54484 205720
rect 54536 205708 54542 205760
rect 370498 205708 370504 205760
rect 370556 205748 370562 205760
rect 371878 205748 371884 205760
rect 370556 205720 371884 205748
rect 370556 205708 370562 205720
rect 371878 205708 371884 205720
rect 371936 205708 371942 205760
rect 56870 205640 56876 205692
rect 56928 205680 56934 205692
rect 56928 205652 58020 205680
rect 56928 205640 56934 205652
rect 57992 205612 58020 205652
rect 188338 205640 188344 205692
rect 188396 205680 188402 205692
rect 580166 205680 580172 205692
rect 188396 205652 580172 205680
rect 188396 205640 188402 205652
rect 580166 205640 580172 205652
rect 580224 205640 580230 205692
rect 59998 205612 60004 205624
rect 57992 205584 60004 205612
rect 59998 205572 60004 205584
rect 60056 205572 60062 205624
rect 384390 205436 384396 205488
rect 384448 205476 384454 205488
rect 388438 205476 388444 205488
rect 384448 205448 388444 205476
rect 384448 205436 384454 205448
rect 388438 205436 388444 205448
rect 388496 205436 388502 205488
rect 61378 204892 61384 204944
rect 61436 204932 61442 204944
rect 75178 204932 75184 204944
rect 61436 204904 75184 204932
rect 61436 204892 61442 204904
rect 75178 204892 75184 204904
rect 75236 204892 75242 204944
rect 68278 204212 68284 204264
rect 68336 204252 68342 204264
rect 69658 204252 69664 204264
rect 68336 204224 69664 204252
rect 68336 204212 68342 204224
rect 69658 204212 69664 204224
rect 69716 204212 69722 204264
rect 385678 204212 385684 204264
rect 385736 204252 385742 204264
rect 391198 204252 391204 204264
rect 385736 204224 391204 204252
rect 385736 204212 385742 204224
rect 391198 204212 391204 204224
rect 391256 204212 391262 204264
rect 382918 203328 382924 203380
rect 382976 203368 382982 203380
rect 384390 203368 384396 203380
rect 382976 203340 384396 203368
rect 382976 203328 382982 203340
rect 384390 203328 384396 203340
rect 384448 203328 384454 203380
rect 87598 202784 87604 202836
rect 87656 202824 87662 202836
rect 93118 202824 93124 202836
rect 87656 202796 93124 202824
rect 87656 202784 87662 202796
rect 93118 202784 93124 202796
rect 93176 202784 93182 202836
rect 78674 202104 78680 202156
rect 78732 202144 78738 202156
rect 88058 202144 88064 202156
rect 78732 202116 88064 202144
rect 78732 202104 78738 202116
rect 88058 202104 88064 202116
rect 88116 202104 88122 202156
rect 111058 202104 111064 202156
rect 111116 202144 111122 202156
rect 126882 202144 126888 202156
rect 111116 202116 126888 202144
rect 111116 202104 111122 202116
rect 126882 202104 126888 202116
rect 126940 202104 126946 202156
rect 147766 202104 147772 202156
rect 147824 202144 147830 202156
rect 176654 202144 176660 202156
rect 147824 202116 176660 202144
rect 147824 202104 147830 202116
rect 176654 202104 176660 202116
rect 176712 202104 176718 202156
rect 50430 201900 50436 201952
rect 50488 201940 50494 201952
rect 57238 201940 57244 201952
rect 50488 201912 57244 201940
rect 50488 201900 50494 201912
rect 57238 201900 57244 201912
rect 57296 201900 57302 201952
rect 3142 201832 3148 201884
rect 3200 201872 3206 201884
rect 7558 201872 7564 201884
rect 3200 201844 7564 201872
rect 3200 201832 3206 201844
rect 7558 201832 7564 201844
rect 7616 201832 7622 201884
rect 155954 199384 155960 199436
rect 156012 199424 156018 199436
rect 296714 199424 296720 199436
rect 156012 199396 296720 199424
rect 156012 199384 156018 199396
rect 296714 199384 296720 199396
rect 296772 199384 296778 199436
rect 88058 198704 88064 198756
rect 88116 198744 88122 198756
rect 90358 198744 90364 198756
rect 88116 198716 90364 198744
rect 88116 198704 88122 198716
rect 90358 198704 90364 198716
rect 90416 198704 90422 198756
rect 148962 197956 148968 198008
rect 149020 197996 149026 198008
rect 207014 197996 207020 198008
rect 149020 197968 207020 197996
rect 149020 197956 149026 197968
rect 207014 197956 207020 197968
rect 207072 197956 207078 198008
rect 154482 197412 154488 197464
rect 154540 197452 154546 197464
rect 155954 197452 155960 197464
rect 154540 197424 155960 197452
rect 154540 197412 154546 197424
rect 155954 197412 155960 197424
rect 156012 197412 156018 197464
rect 166258 197344 166264 197396
rect 166316 197384 166322 197396
rect 167638 197384 167644 197396
rect 166316 197356 167644 197384
rect 166316 197344 166322 197356
rect 167638 197344 167644 197356
rect 167696 197344 167702 197396
rect 59998 197276 60004 197328
rect 60056 197316 60062 197328
rect 65518 197316 65524 197328
rect 60056 197288 65524 197316
rect 60056 197276 60062 197288
rect 65518 197276 65524 197288
rect 65576 197276 65582 197328
rect 152734 197276 152740 197328
rect 152792 197316 152798 197328
rect 157978 197316 157984 197328
rect 152792 197288 157984 197316
rect 152792 197276 152798 197288
rect 157978 197276 157984 197288
rect 158036 197276 158042 197328
rect 380894 196868 380900 196920
rect 380952 196908 380958 196920
rect 382918 196908 382924 196920
rect 380952 196880 382924 196908
rect 380952 196868 380958 196880
rect 382918 196868 382924 196880
rect 382976 196868 382982 196920
rect 138658 196732 138664 196784
rect 138716 196772 138722 196784
rect 164234 196772 164240 196784
rect 138716 196744 164240 196772
rect 138716 196732 138722 196744
rect 164234 196732 164240 196744
rect 164292 196732 164298 196784
rect 151170 196664 151176 196716
rect 151228 196704 151234 196716
rect 235994 196704 236000 196716
rect 151228 196676 236000 196704
rect 151228 196664 151234 196676
rect 235994 196664 236000 196676
rect 236052 196664 236058 196716
rect 155954 196596 155960 196648
rect 156012 196636 156018 196648
rect 327074 196636 327080 196648
rect 156012 196608 327080 196636
rect 156012 196596 156018 196608
rect 327074 196596 327080 196608
rect 327132 196596 327138 196648
rect 126882 196324 126888 196376
rect 126940 196364 126946 196376
rect 128998 196364 129004 196376
rect 126940 196336 129004 196364
rect 126940 196324 126946 196336
rect 128998 196324 129004 196336
rect 129056 196324 129062 196376
rect 56594 195916 56600 195968
rect 56652 195956 56658 195968
rect 138106 195956 138112 195968
rect 56652 195928 138112 195956
rect 56652 195916 56658 195928
rect 138106 195916 138112 195928
rect 138164 195916 138170 195968
rect 160094 195916 160100 195968
rect 160152 195956 160158 195968
rect 386414 195956 386420 195968
rect 160152 195928 386420 195956
rect 160152 195916 160158 195928
rect 386414 195916 386420 195928
rect 386472 195916 386478 195968
rect 86954 195848 86960 195900
rect 87012 195888 87018 195900
rect 139394 195888 139400 195900
rect 87012 195860 139400 195888
rect 87012 195848 87018 195860
rect 139394 195848 139400 195860
rect 139452 195848 139458 195900
rect 157610 195848 157616 195900
rect 157668 195888 157674 195900
rect 266998 195888 267004 195900
rect 157668 195860 267004 195888
rect 157668 195848 157674 195860
rect 266998 195848 267004 195860
rect 267056 195848 267062 195900
rect 115934 194556 115940 194608
rect 115992 194596 115998 194608
rect 140774 194596 140780 194608
rect 115992 194568 140780 194596
rect 115992 194556 115998 194568
rect 140774 194556 140780 194568
rect 140832 194556 140838 194608
rect 47578 194488 47584 194540
rect 47636 194528 47642 194540
rect 54570 194528 54576 194540
rect 47636 194500 54576 194528
rect 47636 194488 47642 194500
rect 54570 194488 54576 194500
rect 54628 194488 54634 194540
rect 380158 193944 380164 193996
rect 380216 193984 380222 193996
rect 385678 193984 385684 193996
rect 380216 193956 385684 193984
rect 380216 193944 380222 193956
rect 385678 193944 385684 193956
rect 385736 193944 385742 193996
rect 166166 193808 166172 193860
rect 166224 193848 166230 193860
rect 380894 193848 380900 193860
rect 166224 193820 380900 193848
rect 166224 193808 166230 193820
rect 380894 193808 380900 193820
rect 380952 193808 380958 193860
rect 54478 192448 54484 192500
rect 54536 192488 54542 192500
rect 58618 192488 58624 192500
rect 54536 192460 58624 192488
rect 54536 192448 54542 192460
rect 58618 192448 58624 192460
rect 58676 192448 58682 192500
rect 180058 191836 180064 191888
rect 180116 191876 180122 191888
rect 580166 191876 580172 191888
rect 180116 191848 580172 191876
rect 180116 191836 180122 191848
rect 580166 191836 580172 191848
rect 580224 191836 580230 191888
rect 144730 190476 144736 190528
rect 144788 190516 144794 190528
rect 144788 190488 144960 190516
rect 144788 190476 144794 190488
rect 144932 190312 144960 190488
rect 145006 190312 145012 190324
rect 144932 190284 145012 190312
rect 145006 190272 145012 190284
rect 145064 190272 145070 190324
rect 54570 189728 54576 189780
rect 54628 189768 54634 189780
rect 60734 189768 60740 189780
rect 54628 189740 60740 189768
rect 54628 189728 54634 189740
rect 60734 189728 60740 189740
rect 60792 189728 60798 189780
rect 93118 189252 93124 189304
rect 93176 189292 93182 189304
rect 94498 189292 94504 189304
rect 93176 189264 94504 189292
rect 93176 189252 93182 189264
rect 94498 189252 94504 189264
rect 94556 189252 94562 189304
rect 387058 189048 387064 189100
rect 387116 189088 387122 189100
rect 394050 189088 394056 189100
rect 387116 189060 394056 189088
rect 387116 189048 387122 189060
rect 394050 189048 394056 189060
rect 394108 189048 394114 189100
rect 144730 188912 144736 188964
rect 144788 188952 144794 188964
rect 145006 188952 145012 188964
rect 144788 188924 145012 188952
rect 144788 188912 144794 188924
rect 145006 188912 145012 188924
rect 145064 188912 145070 188964
rect 75178 187756 75184 187808
rect 75236 187796 75242 187808
rect 80054 187796 80060 187808
rect 75236 187768 80060 187796
rect 75236 187756 75242 187768
rect 80054 187756 80060 187768
rect 80112 187756 80118 187808
rect 2774 187688 2780 187740
rect 2832 187728 2838 187740
rect 5258 187728 5264 187740
rect 2832 187700 5264 187728
rect 2832 187688 2838 187700
rect 5258 187688 5264 187700
rect 5316 187688 5322 187740
rect 69658 186328 69664 186380
rect 69716 186368 69722 186380
rect 71130 186368 71136 186380
rect 69716 186340 71136 186368
rect 69716 186328 69722 186340
rect 71130 186328 71136 186340
rect 71188 186328 71194 186380
rect 62758 186056 62764 186108
rect 62816 186096 62822 186108
rect 64138 186096 64144 186108
rect 62816 186068 64144 186096
rect 62816 186056 62822 186068
rect 64138 186056 64144 186068
rect 64196 186056 64202 186108
rect 128998 185580 129004 185632
rect 129056 185620 129062 185632
rect 132402 185620 132408 185632
rect 129056 185592 132408 185620
rect 129056 185580 129062 185592
rect 132402 185580 132408 185592
rect 132460 185580 132466 185632
rect 60734 184832 60740 184884
rect 60792 184872 60798 184884
rect 65610 184872 65616 184884
rect 60792 184844 65616 184872
rect 60792 184832 60798 184844
rect 65610 184832 65616 184844
rect 65668 184832 65674 184884
rect 94498 184832 94504 184884
rect 94556 184872 94562 184884
rect 97258 184872 97264 184884
rect 94556 184844 97264 184872
rect 94556 184832 94562 184844
rect 97258 184832 97264 184844
rect 97316 184832 97322 184884
rect 57238 184152 57244 184204
rect 57296 184192 57302 184204
rect 65794 184192 65800 184204
rect 57296 184164 65800 184192
rect 57296 184152 57302 184164
rect 65794 184152 65800 184164
rect 65852 184152 65858 184204
rect 71130 183472 71136 183524
rect 71188 183512 71194 183524
rect 72510 183512 72516 183524
rect 71188 183484 72516 183512
rect 71188 183472 71194 183484
rect 72510 183472 72516 183484
rect 72568 183472 72574 183524
rect 167638 183472 167644 183524
rect 167696 183512 167702 183524
rect 169110 183512 169116 183524
rect 167696 183484 169116 183512
rect 167696 183472 167702 183484
rect 169110 183472 169116 183484
rect 169168 183472 169174 183524
rect 132402 183268 132408 183320
rect 132460 183308 132466 183320
rect 135898 183308 135904 183320
rect 132460 183280 135904 183308
rect 132460 183268 132466 183280
rect 135898 183268 135904 183280
rect 135956 183268 135962 183320
rect 80054 182792 80060 182844
rect 80112 182832 80118 182844
rect 88978 182832 88984 182844
rect 80112 182804 88984 182832
rect 80112 182792 80118 182804
rect 88978 182792 88984 182804
rect 89036 182792 89042 182844
rect 58618 182452 58624 182504
rect 58676 182492 58682 182504
rect 64874 182492 64880 182504
rect 58676 182464 64880 182492
rect 58676 182452 58682 182464
rect 64874 182452 64880 182464
rect 64932 182452 64938 182504
rect 90358 181432 90364 181484
rect 90416 181472 90422 181484
rect 100018 181472 100024 181484
rect 90416 181444 100024 181472
rect 90416 181432 90422 181444
rect 100018 181432 100024 181444
rect 100076 181432 100082 181484
rect 144914 180956 144920 181008
rect 144972 180996 144978 181008
rect 144972 180968 153194 180996
rect 144972 180956 144978 180968
rect 153166 180792 153194 180968
rect 153930 180792 153936 180804
rect 153166 180764 153936 180792
rect 153930 180752 153936 180764
rect 153988 180752 153994 180804
rect 154390 180616 154396 180668
rect 154448 180616 154454 180668
rect 65794 180548 65800 180600
rect 65852 180588 65858 180600
rect 68370 180588 68376 180600
rect 65852 180560 68376 180588
rect 65852 180548 65858 180560
rect 68370 180548 68376 180560
rect 68428 180548 68434 180600
rect 154408 180180 154436 180616
rect 154408 180152 154574 180180
rect 121454 180072 121460 180124
rect 121512 180112 121518 180124
rect 136358 180112 136364 180124
rect 121512 180084 136364 180112
rect 121512 180072 121518 180084
rect 136358 180072 136364 180084
rect 136416 180072 136422 180124
rect 154546 180112 154574 180152
rect 157794 180112 157800 180124
rect 154546 180084 157800 180112
rect 157794 180072 157800 180084
rect 157852 180072 157858 180124
rect 158622 180072 158628 180124
rect 158680 180112 158686 180124
rect 165614 180112 165620 180124
rect 158680 180084 165620 180112
rect 158680 180072 158686 180084
rect 165614 180072 165620 180084
rect 165672 180072 165678 180124
rect 65518 179868 65524 179920
rect 65576 179908 65582 179920
rect 66990 179908 66996 179920
rect 65576 179880 66996 179908
rect 65576 179868 65582 179880
rect 66990 179868 66996 179880
rect 67048 179868 67054 179920
rect 135990 178848 135996 178900
rect 136048 178888 136054 178900
rect 136542 178888 136548 178900
rect 136048 178860 136548 178888
rect 136048 178848 136054 178860
rect 136542 178848 136548 178860
rect 136600 178848 136606 178900
rect 122834 178644 122840 178696
rect 122892 178684 122898 178696
rect 136450 178684 136456 178696
rect 122892 178656 136456 178684
rect 122892 178644 122898 178656
rect 136450 178644 136456 178656
rect 136508 178644 136514 178696
rect 72510 178032 72516 178084
rect 72568 178072 72574 178084
rect 73798 178072 73804 178084
rect 72568 178044 73804 178072
rect 72568 178032 72574 178044
rect 73798 178032 73804 178044
rect 73856 178032 73862 178084
rect 166534 178032 166540 178084
rect 166592 178072 166598 178084
rect 580166 178072 580172 178084
rect 166592 178044 580172 178072
rect 166592 178032 166598 178044
rect 580166 178032 580172 178044
rect 580224 178032 580230 178084
rect 159450 177828 159456 177880
rect 159508 177868 159514 177880
rect 167638 177868 167644 177880
rect 159508 177840 167644 177868
rect 159508 177828 159514 177840
rect 167638 177828 167644 177840
rect 167696 177828 167702 177880
rect 124214 177284 124220 177336
rect 124272 177324 124278 177336
rect 135990 177324 135996 177336
rect 124272 177296 135996 177324
rect 124272 177284 124278 177296
rect 135990 177284 135996 177296
rect 136048 177284 136054 177336
rect 64874 177148 64880 177200
rect 64932 177188 64938 177200
rect 68462 177188 68468 177200
rect 64932 177160 68468 177188
rect 64932 177148 64938 177160
rect 68462 177148 68468 177160
rect 68520 177148 68526 177200
rect 149330 176468 149336 176520
rect 149388 176508 149394 176520
rect 149388 176480 153976 176508
rect 149388 176468 149394 176480
rect 153948 176452 153976 176480
rect 153930 176400 153936 176452
rect 153988 176400 153994 176452
rect 154390 176400 154396 176452
rect 154448 176400 154454 176452
rect 126974 176060 126980 176112
rect 127032 176100 127038 176112
rect 136266 176100 136272 176112
rect 127032 176072 136272 176100
rect 127032 176060 127038 176072
rect 136266 176060 136272 176072
rect 136324 176060 136330 176112
rect 125594 175924 125600 175976
rect 125652 175964 125658 175976
rect 136174 175964 136180 175976
rect 125652 175936 136180 175964
rect 125652 175924 125658 175936
rect 136174 175924 136180 175936
rect 136232 175924 136238 175976
rect 144086 175924 144092 175976
rect 144144 175964 144150 175976
rect 149330 175964 149336 175976
rect 144144 175936 149336 175964
rect 144144 175924 144150 175936
rect 149330 175924 149336 175936
rect 149388 175924 149394 175976
rect 154408 175964 154436 176400
rect 169110 176332 169116 176384
rect 169168 176372 169174 176384
rect 169754 176372 169760 176384
rect 169168 176344 169760 176372
rect 169168 176332 169174 176344
rect 169754 176332 169760 176344
rect 169812 176332 169818 176384
rect 162486 175964 162492 175976
rect 154408 175936 162492 175964
rect 162486 175924 162492 175936
rect 162544 175924 162550 175976
rect 144454 175516 144460 175568
rect 144512 175556 144518 175568
rect 149974 175556 149980 175568
rect 144512 175528 149980 175556
rect 144512 175516 144518 175528
rect 149974 175516 149980 175528
rect 150032 175516 150038 175568
rect 128354 175176 128360 175228
rect 128412 175216 128418 175228
rect 136358 175216 136364 175228
rect 128412 175188 136364 175216
rect 128412 175176 128418 175188
rect 136358 175176 136364 175188
rect 136416 175176 136422 175228
rect 141602 174700 141608 174752
rect 141660 174700 141666 174752
rect 143074 174700 143080 174752
rect 143132 174740 143138 174752
rect 143132 174712 143534 174740
rect 143132 174700 143138 174712
rect 141620 174468 141648 174700
rect 143506 174536 143534 174712
rect 152458 174632 152464 174684
rect 152516 174672 152522 174684
rect 156506 174672 156512 174684
rect 152516 174644 156512 174672
rect 152516 174632 152522 174644
rect 156506 174632 156512 174644
rect 156564 174632 156570 174684
rect 161474 174536 161480 174548
rect 143506 174508 161480 174536
rect 161474 174496 161480 174508
rect 161532 174496 161538 174548
rect 366358 174496 366364 174548
rect 366416 174536 366422 174548
rect 380158 174536 380164 174548
rect 366416 174508 380164 174536
rect 366416 174496 366422 174508
rect 380158 174496 380164 174508
rect 380216 174496 380222 174548
rect 385678 174496 385684 174548
rect 385736 174536 385742 174548
rect 387058 174536 387064 174548
rect 385736 174508 387064 174536
rect 385736 174496 385742 174508
rect 387058 174496 387064 174508
rect 387116 174496 387122 174548
rect 141620 174440 142154 174468
rect 142126 174332 142154 174440
rect 166994 174332 167000 174344
rect 142126 174304 167000 174332
rect 166994 174292 167000 174304
rect 167052 174292 167058 174344
rect 133874 173884 133880 173936
rect 133932 173924 133938 173936
rect 137370 173924 137376 173936
rect 133932 173896 137376 173924
rect 133932 173884 133938 173896
rect 137370 173884 137376 173896
rect 137428 173884 137434 173936
rect 135898 173136 135904 173188
rect 135956 173176 135962 173188
rect 135956 173148 142154 173176
rect 135956 173136 135962 173148
rect 142126 172904 142154 173148
rect 148318 172932 148324 172984
rect 148376 172972 148382 172984
rect 149054 172972 149060 172984
rect 148376 172944 149060 172972
rect 148376 172932 148382 172944
rect 149054 172932 149060 172944
rect 149112 172932 149118 172984
rect 149330 172932 149336 172984
rect 149388 172972 149394 172984
rect 151446 172972 151452 172984
rect 149388 172944 151452 172972
rect 149388 172932 149394 172944
rect 151446 172932 151452 172944
rect 151504 172932 151510 172984
rect 162486 172932 162492 172984
rect 162544 172972 162550 172984
rect 165430 172972 165436 172984
rect 162544 172944 165436 172972
rect 162544 172932 162550 172944
rect 165430 172932 165436 172944
rect 165488 172932 165494 172984
rect 148962 172904 148968 172916
rect 142126 172876 148968 172904
rect 148962 172864 148968 172876
rect 149020 172864 149026 172916
rect 131114 172524 131120 172576
rect 131172 172564 131178 172576
rect 136542 172564 136548 172576
rect 131172 172536 136548 172564
rect 131172 172524 131178 172536
rect 136542 172524 136548 172536
rect 136600 172524 136606 172576
rect 66990 172456 66996 172508
rect 67048 172496 67054 172508
rect 68278 172496 68284 172508
rect 67048 172468 68284 172496
rect 67048 172456 67054 172468
rect 68278 172456 68284 172468
rect 68336 172456 68342 172508
rect 65610 172388 65616 172440
rect 65668 172428 65674 172440
rect 71038 172428 71044 172440
rect 65668 172400 71044 172428
rect 65668 172388 65674 172400
rect 71038 172388 71044 172400
rect 71096 172388 71102 172440
rect 138014 172116 138020 172168
rect 138072 172156 138078 172168
rect 140774 172156 140780 172168
rect 138072 172128 140780 172156
rect 138072 172116 138078 172128
rect 140774 172116 140780 172128
rect 140832 172116 140838 172168
rect 135254 171640 135260 171692
rect 135312 171680 135318 171692
rect 138658 171680 138664 171692
rect 135312 171652 138664 171680
rect 135312 171640 135318 171652
rect 138658 171640 138664 171652
rect 138716 171640 138722 171692
rect 169754 171368 169760 171420
rect 169812 171408 169818 171420
rect 171778 171408 171784 171420
rect 169812 171380 171784 171408
rect 169812 171368 169818 171380
rect 171778 171368 171784 171380
rect 171836 171368 171842 171420
rect 132494 171096 132500 171148
rect 132552 171136 132558 171148
rect 136726 171136 136732 171148
rect 132552 171108 136732 171136
rect 132552 171096 132558 171108
rect 136726 171096 136732 171108
rect 136784 171096 136790 171148
rect 148962 170348 148968 170400
rect 149020 170388 149026 170400
rect 162670 170388 162676 170400
rect 149020 170360 162676 170388
rect 149020 170348 149026 170360
rect 162670 170348 162676 170360
rect 162728 170348 162734 170400
rect 118418 168988 118424 169040
rect 118476 169028 118482 169040
rect 158438 169028 158444 169040
rect 118476 169000 158444 169028
rect 118476 168988 118482 169000
rect 158438 168988 158444 169000
rect 158496 168988 158502 169040
rect 68462 168036 68468 168088
rect 68520 168076 68526 168088
rect 71498 168076 71504 168088
rect 68520 168048 71504 168076
rect 68520 168036 68526 168048
rect 71498 168036 71504 168048
rect 71556 168036 71562 168088
rect 162670 167696 162676 167748
rect 162728 167736 162734 167748
rect 172238 167736 172244 167748
rect 162728 167708 172244 167736
rect 162728 167696 162734 167708
rect 172238 167696 172244 167708
rect 172296 167696 172302 167748
rect 118786 167628 118792 167680
rect 118844 167668 118850 167680
rect 580258 167668 580264 167680
rect 118844 167640 580264 167668
rect 118844 167628 118850 167640
rect 580258 167628 580264 167640
rect 580316 167628 580322 167680
rect 384298 167084 384304 167136
rect 384356 167124 384362 167136
rect 385678 167124 385684 167136
rect 384356 167096 385684 167124
rect 384356 167084 384362 167096
rect 385678 167084 385684 167096
rect 385736 167084 385742 167136
rect 68370 166948 68376 167000
rect 68428 166988 68434 167000
rect 71774 166988 71780 167000
rect 68428 166960 71780 166988
rect 68428 166948 68434 166960
rect 71774 166948 71780 166960
rect 71832 166948 71838 167000
rect 142430 166268 142436 166320
rect 142488 166308 142494 166320
rect 142614 166308 142620 166320
rect 142488 166280 142620 166308
rect 142488 166268 142494 166280
rect 142614 166268 142620 166280
rect 142672 166268 142678 166320
rect 226978 165588 226984 165640
rect 227036 165628 227042 165640
rect 580166 165628 580172 165640
rect 227036 165600 580172 165628
rect 227036 165588 227042 165600
rect 580166 165588 580172 165600
rect 580224 165588 580230 165640
rect 97258 165520 97264 165572
rect 97316 165560 97322 165572
rect 98638 165560 98644 165572
rect 97316 165532 98644 165560
rect 97316 165520 97322 165532
rect 98638 165520 98644 165532
rect 98696 165520 98702 165572
rect 380894 165248 380900 165300
rect 380952 165288 380958 165300
rect 384298 165288 384304 165300
rect 380952 165260 384304 165288
rect 380952 165248 380958 165260
rect 384298 165248 384304 165260
rect 384356 165248 384362 165300
rect 172238 164160 172244 164212
rect 172296 164200 172302 164212
rect 175182 164200 175188 164212
rect 172296 164172 175188 164200
rect 172296 164160 172302 164172
rect 175182 164160 175188 164172
rect 175240 164160 175246 164212
rect 71498 163548 71504 163600
rect 71556 163588 71562 163600
rect 82814 163588 82820 163600
rect 71556 163560 82820 163588
rect 71556 163548 71562 163560
rect 82814 163548 82820 163560
rect 82872 163548 82878 163600
rect 71774 163480 71780 163532
rect 71832 163520 71838 163532
rect 86218 163520 86224 163532
rect 71832 163492 86224 163520
rect 71832 163480 71838 163492
rect 86218 163480 86224 163492
rect 86276 163480 86282 163532
rect 380250 163072 380256 163124
rect 380308 163112 380314 163124
rect 380894 163112 380900 163124
rect 380308 163084 380900 163112
rect 380308 163072 380314 163084
rect 380894 163072 380900 163084
rect 380952 163072 380958 163124
rect 3142 162868 3148 162920
rect 3200 162908 3206 162920
rect 180886 162908 180892 162920
rect 3200 162880 180892 162908
rect 3200 162868 3206 162880
rect 180886 162868 180892 162880
rect 180944 162868 180950 162920
rect 9030 162120 9036 162172
rect 9088 162160 9094 162172
rect 182174 162160 182180 162172
rect 9088 162132 182180 162160
rect 9088 162120 9094 162132
rect 182174 162120 182180 162132
rect 182232 162120 182238 162172
rect 118878 160692 118884 160744
rect 118936 160732 118942 160744
rect 580442 160732 580448 160744
rect 118936 160704 580448 160732
rect 118936 160692 118942 160704
rect 580442 160692 580448 160704
rect 580500 160692 580506 160744
rect 73798 160080 73804 160132
rect 73856 160120 73862 160132
rect 73856 160092 74534 160120
rect 73856 160080 73862 160092
rect 74506 160052 74534 160092
rect 76558 160052 76564 160064
rect 74506 160024 76564 160052
rect 76558 160012 76564 160024
rect 76616 160012 76622 160064
rect 64138 159332 64144 159384
rect 64196 159372 64202 159384
rect 66162 159372 66168 159384
rect 64196 159344 66168 159372
rect 64196 159332 64202 159344
rect 66162 159332 66168 159344
rect 66220 159332 66226 159384
rect 82814 159060 82820 159112
rect 82872 159100 82878 159112
rect 86586 159100 86592 159112
rect 82872 159072 86592 159100
rect 82872 159060 82878 159072
rect 86586 159060 86592 159072
rect 86644 159060 86650 159112
rect 175182 158856 175188 158908
rect 175240 158896 175246 158908
rect 177298 158896 177304 158908
rect 175240 158868 177304 158896
rect 175240 158856 175246 158868
rect 177298 158856 177304 158868
rect 177356 158856 177362 158908
rect 88978 158652 88984 158704
rect 89036 158692 89042 158704
rect 96522 158692 96528 158704
rect 89036 158664 96528 158692
rect 89036 158652 89042 158664
rect 96522 158652 96528 158664
rect 96580 158652 96586 158704
rect 154482 157972 154488 158024
rect 154540 158012 154546 158024
rect 165614 158012 165620 158024
rect 154540 157984 165620 158012
rect 154540 157972 154546 157984
rect 165614 157972 165620 157984
rect 165672 157972 165678 158024
rect 378870 157360 378876 157412
rect 378928 157400 378934 157412
rect 380250 157400 380256 157412
rect 378928 157372 380256 157400
rect 378928 157360 378934 157372
rect 380250 157360 380256 157372
rect 380308 157360 380314 157412
rect 71038 154504 71044 154556
rect 71096 154544 71102 154556
rect 74166 154544 74172 154556
rect 71096 154516 74172 154544
rect 71096 154504 71102 154516
rect 74166 154504 74172 154516
rect 74224 154504 74230 154556
rect 165614 154504 165620 154556
rect 165672 154544 165678 154556
rect 168374 154544 168380 154556
rect 165672 154516 168380 154544
rect 165672 154504 165678 154516
rect 168374 154504 168380 154516
rect 168432 154504 168438 154556
rect 377398 154096 377404 154148
rect 377456 154136 377462 154148
rect 378870 154136 378876 154148
rect 377456 154108 378876 154136
rect 377456 154096 377462 154108
rect 378870 154096 378876 154108
rect 378928 154096 378934 154148
rect 96522 153824 96528 153876
rect 96580 153864 96586 153876
rect 109678 153864 109684 153876
rect 96580 153836 109684 153864
rect 96580 153824 96586 153836
rect 109678 153824 109684 153836
rect 109736 153824 109742 153876
rect 118970 153824 118976 153876
rect 119028 153864 119034 153876
rect 580626 153864 580632 153876
rect 119028 153836 580632 153864
rect 119028 153824 119034 153836
rect 580626 153824 580632 153836
rect 580684 153824 580690 153876
rect 86586 153144 86592 153196
rect 86644 153184 86650 153196
rect 89622 153184 89628 153196
rect 86644 153156 89628 153184
rect 86644 153144 86650 153156
rect 89622 153144 89628 153156
rect 89680 153144 89686 153196
rect 180150 151784 180156 151836
rect 180208 151824 180214 151836
rect 580166 151824 580172 151836
rect 180208 151796 580172 151824
rect 180208 151784 180214 151796
rect 580166 151784 580172 151796
rect 580224 151784 580230 151836
rect 66254 151444 66260 151496
rect 66312 151484 66318 151496
rect 68370 151484 68376 151496
rect 66312 151456 68376 151484
rect 66312 151444 66318 151456
rect 68370 151444 68376 151456
rect 68428 151444 68434 151496
rect 3234 149676 3240 149728
rect 3292 149716 3298 149728
rect 22830 149716 22836 149728
rect 3292 149688 22836 149716
rect 3292 149676 3298 149688
rect 22830 149676 22836 149688
rect 22888 149676 22894 149728
rect 118510 148316 118516 148368
rect 118568 148356 118574 148368
rect 166442 148356 166448 148368
rect 118568 148328 166448 148356
rect 118568 148316 118574 148328
rect 166442 148316 166448 148328
rect 166500 148316 166506 148368
rect 86218 147908 86224 147960
rect 86276 147948 86282 147960
rect 88978 147948 88984 147960
rect 86276 147920 88984 147948
rect 86276 147908 86282 147920
rect 88978 147908 88984 147920
rect 89036 147908 89042 147960
rect 76558 147568 76564 147620
rect 76616 147608 76622 147620
rect 79962 147608 79968 147620
rect 76616 147580 79968 147608
rect 76616 147568 76622 147580
rect 79962 147568 79968 147580
rect 80020 147568 80026 147620
rect 171778 146956 171784 147008
rect 171836 146996 171842 147008
rect 172514 146996 172520 147008
rect 171836 146968 172520 146996
rect 171836 146956 171842 146968
rect 172514 146956 172520 146968
rect 172572 146956 172578 147008
rect 89622 146888 89628 146940
rect 89680 146928 89686 146940
rect 105998 146928 106004 146940
rect 89680 146900 106004 146928
rect 89680 146888 89686 146900
rect 105998 146888 106004 146900
rect 106056 146888 106062 146940
rect 141694 146208 141700 146260
rect 141752 146248 141758 146260
rect 142430 146248 142436 146260
rect 141752 146220 142436 146248
rect 141752 146208 141758 146220
rect 142430 146208 142436 146220
rect 142488 146208 142494 146260
rect 139486 146072 139492 146124
rect 139544 146112 139550 146124
rect 142246 146112 142252 146124
rect 139544 146084 142252 146112
rect 139544 146072 139550 146084
rect 142246 146072 142252 146084
rect 142304 146072 142310 146124
rect 74166 145528 74172 145580
rect 74224 145568 74230 145580
rect 78674 145568 78680 145580
rect 74224 145540 78680 145568
rect 74224 145528 74230 145540
rect 78674 145528 78680 145540
rect 78732 145528 78738 145580
rect 177298 144848 177304 144900
rect 177356 144888 177362 144900
rect 180242 144888 180248 144900
rect 177356 144860 180248 144888
rect 177356 144848 177362 144860
rect 180242 144848 180248 144860
rect 180300 144848 180306 144900
rect 105998 144576 106004 144628
rect 106056 144616 106062 144628
rect 109770 144616 109776 144628
rect 106056 144588 109776 144616
rect 106056 144576 106062 144588
rect 109770 144576 109776 144588
rect 109828 144576 109834 144628
rect 33778 144440 33784 144492
rect 33836 144480 33842 144492
rect 182266 144480 182272 144492
rect 33836 144452 182272 144480
rect 33836 144440 33842 144452
rect 182266 144440 182272 144452
rect 182324 144440 182330 144492
rect 10410 144372 10416 144424
rect 10468 144412 10474 144424
rect 182542 144412 182548 144424
rect 10468 144384 182548 144412
rect 10468 144372 10474 144384
rect 182542 144372 182548 144384
rect 182600 144372 182606 144424
rect 6178 144304 6184 144356
rect 6236 144344 6242 144356
rect 182450 144344 182456 144356
rect 6236 144316 182456 144344
rect 6236 144304 6242 144316
rect 182450 144304 182456 144316
rect 182508 144304 182514 144356
rect 118050 144236 118056 144288
rect 118108 144276 118114 144288
rect 398098 144276 398104 144288
rect 118108 144248 398104 144276
rect 118108 144236 118114 144248
rect 398098 144236 398104 144248
rect 398156 144236 398162 144288
rect 119246 144168 119252 144220
rect 119304 144208 119310 144220
rect 477494 144208 477500 144220
rect 119304 144180 477500 144208
rect 119304 144168 119310 144180
rect 477494 144168 477500 144180
rect 477552 144168 477558 144220
rect 79962 143556 79968 143608
rect 80020 143596 80026 143608
rect 80020 143568 82216 143596
rect 80020 143556 80026 143568
rect 78674 143488 78680 143540
rect 78732 143528 78738 143540
rect 82078 143528 82084 143540
rect 78732 143500 82084 143528
rect 78732 143488 78738 143500
rect 82078 143488 82084 143500
rect 82136 143488 82142 143540
rect 82188 143528 82216 143568
rect 84194 143528 84200 143540
rect 82188 143500 84200 143528
rect 84194 143488 84200 143500
rect 84252 143488 84258 143540
rect 146478 143488 146484 143540
rect 146536 143528 146542 143540
rect 148042 143528 148048 143540
rect 146536 143500 148048 143528
rect 146536 143488 146542 143500
rect 148042 143488 148048 143500
rect 148100 143488 148106 143540
rect 153470 143488 153476 143540
rect 153528 143528 153534 143540
rect 158990 143528 158996 143540
rect 153528 143500 158996 143528
rect 153528 143488 153534 143500
rect 158990 143488 158996 143500
rect 159048 143488 159054 143540
rect 167638 143488 167644 143540
rect 167696 143528 167702 143540
rect 169938 143528 169944 143540
rect 167696 143500 169944 143528
rect 167696 143488 167702 143500
rect 169938 143488 169944 143500
rect 169996 143488 170002 143540
rect 172514 143488 172520 143540
rect 172572 143528 172578 143540
rect 176470 143528 176476 143540
rect 172572 143500 176476 143528
rect 172572 143488 172578 143500
rect 176470 143488 176476 143500
rect 176528 143488 176534 143540
rect 137738 143420 137744 143472
rect 137796 143460 137802 143472
rect 139578 143460 139584 143472
rect 137796 143432 139584 143460
rect 137796 143420 137802 143432
rect 139578 143420 139584 143432
rect 139636 143420 139642 143472
rect 152458 143420 152464 143472
rect 152516 143460 152522 143472
rect 157426 143460 157432 143472
rect 152516 143432 157432 143460
rect 152516 143420 152522 143432
rect 157426 143420 157432 143432
rect 157484 143420 157490 143472
rect 163590 143148 163596 143200
rect 163648 143188 163654 143200
rect 174630 143188 174636 143200
rect 163648 143160 174636 143188
rect 163648 143148 163654 143160
rect 174630 143148 174636 143160
rect 174688 143148 174694 143200
rect 150526 143080 150532 143132
rect 150584 143120 150590 143132
rect 154574 143120 154580 143132
rect 150584 143092 154580 143120
rect 150584 143080 150590 143092
rect 154574 143080 154580 143092
rect 154632 143080 154638 143132
rect 164510 143080 164516 143132
rect 164568 143120 164574 143132
rect 176194 143120 176200 143132
rect 164568 143092 176200 143120
rect 164568 143080 164574 143092
rect 176194 143080 176200 143092
rect 176252 143080 176258 143132
rect 144454 143012 144460 143064
rect 144512 143052 144518 143064
rect 160554 143052 160560 143064
rect 144512 143024 160560 143052
rect 144512 143012 144518 143024
rect 160554 143012 160560 143024
rect 160612 143012 160618 143064
rect 163498 143012 163504 143064
rect 163556 143052 163562 143064
rect 178034 143052 178040 143064
rect 163556 143024 178040 143052
rect 163556 143012 163562 143024
rect 178034 143012 178040 143024
rect 178092 143012 178098 143064
rect 142522 142944 142528 142996
rect 142580 142984 142586 142996
rect 173066 142984 173072 142996
rect 142580 142956 173072 142984
rect 142580 142944 142586 142956
rect 173066 142944 173072 142956
rect 173124 142944 173130 142996
rect 118142 142876 118148 142928
rect 118200 142916 118206 142928
rect 398190 142916 398196 142928
rect 118200 142888 398196 142916
rect 118200 142876 118206 142888
rect 398190 142876 398196 142888
rect 398248 142876 398254 142928
rect 118234 142808 118240 142860
rect 118292 142848 118298 142860
rect 418890 142848 418896 142860
rect 118292 142820 418896 142848
rect 118292 142808 118298 142820
rect 418890 142808 418896 142820
rect 418948 142808 418954 142860
rect 149514 142196 149520 142248
rect 149572 142196 149578 142248
rect 149532 142168 149560 142196
rect 152734 142168 152740 142180
rect 149532 142140 152740 142168
rect 152734 142128 152740 142140
rect 152792 142128 152798 142180
rect 157334 142128 157340 142180
rect 157392 142168 157398 142180
rect 163682 142168 163688 142180
rect 157392 142140 163688 142168
rect 157392 142128 157398 142140
rect 163682 142128 163688 142140
rect 163740 142128 163746 142180
rect 40034 141720 40040 141772
rect 40092 141760 40098 141772
rect 181162 141760 181168 141772
rect 40092 141732 181168 141760
rect 40092 141720 40098 141732
rect 181162 141720 181168 141732
rect 181220 141720 181226 141772
rect 4890 141652 4896 141704
rect 4948 141692 4954 141704
rect 182818 141692 182824 141704
rect 4948 141664 182824 141692
rect 4948 141652 4954 141664
rect 182818 141652 182824 141664
rect 182876 141652 182882 141704
rect 119338 141584 119344 141636
rect 119396 141624 119402 141636
rect 412634 141624 412640 141636
rect 119396 141596 412640 141624
rect 119396 141584 119402 141596
rect 412634 141584 412640 141596
rect 412692 141584 412698 141636
rect 120718 141516 120724 141568
rect 120776 141556 120782 141568
rect 542354 141556 542360 141568
rect 120776 141528 542360 141556
rect 120776 141516 120782 141528
rect 542354 141516 542360 141528
rect 542412 141516 542418 141568
rect 119154 141448 119160 141500
rect 119212 141488 119218 141500
rect 580810 141488 580816 141500
rect 119212 141460 580816 141488
rect 119212 141448 119218 141460
rect 580810 141448 580816 141460
rect 580868 141448 580874 141500
rect 119062 141380 119068 141432
rect 119120 141420 119126 141432
rect 580902 141420 580908 141432
rect 119120 141392 580908 141420
rect 119120 141380 119126 141392
rect 580902 141380 580908 141392
rect 580960 141380 580966 141432
rect 176470 141312 176476 141364
rect 176528 141352 176534 141364
rect 181070 141352 181076 141364
rect 176528 141324 181076 141352
rect 176528 141312 176534 141324
rect 181070 141312 181076 141324
rect 181128 141312 181134 141364
rect 367370 140768 367376 140820
rect 367428 140808 367434 140820
rect 370498 140808 370504 140820
rect 367428 140780 370504 140808
rect 367428 140768 367434 140780
rect 370498 140768 370504 140780
rect 370556 140768 370562 140820
rect 109678 140156 109684 140208
rect 109736 140196 109742 140208
rect 180334 140196 180340 140208
rect 109736 140168 180340 140196
rect 109736 140156 109742 140168
rect 180334 140156 180340 140168
rect 180392 140156 180398 140208
rect 10318 140088 10324 140140
rect 10376 140128 10382 140140
rect 182726 140128 182732 140140
rect 10376 140100 182732 140128
rect 10376 140088 10382 140100
rect 182726 140088 182732 140100
rect 182784 140088 182790 140140
rect 4798 140020 4804 140072
rect 4856 140060 4862 140072
rect 182634 140060 182640 140072
rect 4856 140032 182640 140060
rect 4856 140020 4862 140032
rect 182634 140020 182640 140032
rect 182692 140020 182698 140072
rect 375006 139816 375012 139868
rect 375064 139856 375070 139868
rect 377398 139856 377404 139868
rect 375064 139828 377404 139856
rect 375064 139816 375070 139828
rect 377398 139816 377404 139828
rect 377456 139816 377462 139868
rect 98638 139612 98644 139664
rect 98696 139652 98702 139664
rect 100846 139652 100852 139664
rect 98696 139624 100852 139652
rect 98696 139612 98702 139624
rect 100846 139612 100852 139624
rect 100904 139612 100910 139664
rect 62758 139476 62764 139528
rect 62816 139516 62822 139528
rect 182358 139516 182364 139528
rect 62816 139488 182364 139516
rect 62816 139476 62822 139488
rect 182358 139476 182364 139488
rect 182416 139476 182422 139528
rect 118326 139408 118332 139460
rect 118384 139448 118390 139460
rect 580166 139448 580172 139460
rect 118384 139420 580172 139448
rect 118384 139408 118390 139420
rect 580166 139408 580172 139420
rect 580224 139408 580230 139460
rect 3878 138660 3884 138712
rect 3936 138700 3942 138712
rect 25498 138700 25504 138712
rect 3936 138672 25504 138700
rect 3936 138660 3942 138672
rect 25498 138660 25504 138672
rect 25556 138660 25562 138712
rect 88978 138660 88984 138712
rect 89036 138700 89042 138712
rect 97258 138700 97264 138712
rect 89036 138672 97264 138700
rect 89036 138660 89042 138672
rect 97258 138660 97264 138672
rect 97316 138660 97322 138712
rect 373258 137368 373264 137420
rect 373316 137408 373322 137420
rect 375006 137408 375012 137420
rect 373316 137380 375012 137408
rect 373316 137368 373322 137380
rect 375006 137368 375012 137380
rect 375064 137368 375070 137420
rect 84194 137300 84200 137352
rect 84252 137340 84258 137352
rect 87598 137340 87604 137352
rect 84252 137312 87604 137340
rect 84252 137300 84258 137312
rect 87598 137300 87604 137312
rect 87656 137300 87662 137352
rect 3234 136688 3240 136740
rect 3292 136728 3298 136740
rect 116578 136728 116584 136740
rect 3292 136700 116584 136728
rect 3292 136688 3298 136700
rect 116578 136688 116584 136700
rect 116636 136688 116642 136740
rect 3878 136620 3884 136672
rect 3936 136660 3942 136672
rect 117314 136660 117320 136672
rect 3936 136632 117320 136660
rect 3936 136620 3942 136632
rect 117314 136620 117320 136632
rect 117372 136620 117378 136672
rect 365530 136212 365536 136264
rect 365588 136252 365594 136264
rect 367370 136252 367376 136264
rect 365588 136224 367376 136252
rect 365588 136212 365594 136224
rect 367370 136212 367376 136224
rect 367428 136212 367434 136264
rect 4062 135260 4068 135312
rect 4120 135300 4126 135312
rect 117314 135300 117320 135312
rect 4120 135272 117320 135300
rect 4120 135260 4126 135272
rect 117314 135260 117320 135272
rect 117372 135260 117378 135312
rect 100846 135192 100852 135244
rect 100904 135232 100910 135244
rect 102870 135232 102876 135244
rect 100904 135204 102876 135232
rect 100904 135192 100910 135204
rect 102870 135192 102876 135204
rect 102928 135192 102934 135244
rect 182358 134444 182364 134496
rect 182416 134484 182422 134496
rect 182634 134484 182640 134496
rect 182416 134456 182640 134484
rect 182416 134444 182422 134456
rect 182634 134444 182640 134456
rect 182692 134444 182698 134496
rect 3234 133900 3240 133952
rect 3292 133940 3298 133952
rect 117314 133940 117320 133952
rect 3292 133912 117320 133940
rect 3292 133900 3298 133912
rect 117314 133900 117320 133912
rect 117372 133900 117378 133952
rect 362218 133900 362224 133952
rect 362276 133940 362282 133952
rect 365530 133940 365536 133952
rect 362276 133912 365536 133940
rect 362276 133900 362282 133912
rect 365530 133900 365536 133912
rect 365588 133900 365594 133952
rect 25498 132404 25504 132456
rect 25556 132444 25562 132456
rect 117314 132444 117320 132456
rect 25556 132416 117320 132444
rect 25556 132404 25562 132416
rect 117314 132404 117320 132416
rect 117372 132404 117378 132456
rect 68278 132132 68284 132184
rect 68336 132172 68342 132184
rect 69014 132172 69020 132184
rect 68336 132144 69020 132172
rect 68336 132132 68342 132144
rect 69014 132132 69020 132144
rect 69072 132132 69078 132184
rect 109770 131724 109776 131776
rect 109828 131764 109834 131776
rect 117958 131764 117964 131776
rect 109828 131736 117964 131764
rect 109828 131724 109834 131736
rect 117958 131724 117964 131736
rect 118016 131724 118022 131776
rect 7558 131044 7564 131096
rect 7616 131084 7622 131096
rect 117314 131084 117320 131096
rect 7616 131056 117320 131084
rect 7616 131044 7622 131056
rect 117314 131044 117320 131056
rect 117372 131044 117378 131096
rect 69014 130976 69020 131028
rect 69072 131016 69078 131028
rect 74902 131016 74908 131028
rect 69072 130988 74908 131016
rect 69072 130976 69078 130988
rect 74902 130976 74908 130988
rect 74960 130976 74966 131028
rect 87598 129752 87604 129804
rect 87656 129792 87662 129804
rect 90358 129792 90364 129804
rect 87656 129764 90364 129792
rect 87656 129752 87662 129764
rect 90358 129752 90364 129764
rect 90416 129752 90422 129804
rect 373258 129792 373264 129804
rect 371252 129764 373264 129792
rect 22738 129684 22744 129736
rect 22796 129724 22802 129736
rect 117314 129724 117320 129736
rect 22796 129696 117320 129724
rect 22796 129684 22802 129696
rect 117314 129684 117320 129696
rect 117372 129684 117378 129736
rect 369854 129684 369860 129736
rect 369912 129724 369918 129736
rect 371252 129724 371280 129764
rect 373258 129752 373264 129764
rect 373316 129752 373322 129804
rect 369912 129696 371280 129724
rect 369912 129684 369918 129696
rect 102870 129616 102876 129668
rect 102928 129656 102934 129668
rect 104158 129656 104164 129668
rect 102928 129628 104164 129656
rect 102928 129616 102934 129628
rect 104158 129616 104164 129628
rect 104216 129616 104222 129668
rect 68370 129004 68376 129056
rect 68428 129044 68434 129056
rect 69658 129044 69664 129056
rect 68428 129016 69664 129044
rect 68428 129004 68434 129016
rect 69658 129004 69664 129016
rect 69716 129004 69722 129056
rect 74902 129004 74908 129056
rect 74960 129044 74966 129056
rect 84838 129044 84844 129056
rect 74960 129016 84844 129044
rect 74960 129004 74966 129016
rect 84838 129004 84844 129016
rect 84896 129004 84902 129056
rect 22830 128256 22836 128308
rect 22888 128296 22894 128308
rect 117314 128296 117320 128308
rect 22888 128268 117320 128296
rect 22888 128256 22894 128268
rect 117314 128256 117320 128268
rect 117372 128256 117378 128308
rect 180334 128256 180340 128308
rect 180392 128296 180398 128308
rect 182174 128296 182180 128308
rect 180392 128268 182180 128296
rect 180392 128256 180398 128268
rect 182174 128256 182180 128268
rect 182232 128256 182238 128308
rect 24118 126896 24124 126948
rect 24176 126936 24182 126948
rect 117314 126936 117320 126948
rect 24176 126908 117320 126936
rect 24176 126896 24182 126908
rect 117314 126896 117320 126908
rect 117372 126896 117378 126948
rect 184198 125604 184204 125656
rect 184256 125644 184262 125656
rect 580074 125644 580080 125656
rect 184256 125616 580080 125644
rect 184256 125604 184262 125616
rect 580074 125604 580080 125616
rect 580132 125604 580138 125656
rect 8938 125536 8944 125588
rect 8996 125576 9002 125588
rect 117314 125576 117320 125588
rect 8996 125548 117320 125576
rect 8996 125536 9002 125548
rect 117314 125536 117320 125548
rect 117372 125536 117378 125588
rect 367738 125128 367744 125180
rect 367796 125168 367802 125180
rect 369762 125168 369768 125180
rect 367796 125140 369768 125168
rect 367796 125128 367802 125140
rect 369762 125128 369768 125140
rect 369820 125128 369826 125180
rect 4982 124108 4988 124160
rect 5040 124148 5046 124160
rect 117314 124148 117320 124160
rect 5040 124120 117320 124148
rect 5040 124108 5046 124120
rect 117314 124108 117320 124120
rect 117372 124108 117378 124160
rect 97258 124040 97264 124092
rect 97316 124080 97322 124092
rect 100110 124080 100116 124092
rect 97316 124052 100116 124080
rect 97316 124040 97322 124052
rect 100110 124040 100116 124052
rect 100168 124040 100174 124092
rect 82078 123428 82084 123480
rect 82136 123468 82142 123480
rect 90450 123468 90456 123480
rect 82136 123440 90456 123468
rect 82136 123428 82142 123440
rect 90450 123428 90456 123440
rect 90508 123428 90514 123480
rect 43438 122748 43444 122800
rect 43496 122788 43502 122800
rect 117314 122788 117320 122800
rect 43496 122760 117320 122788
rect 43496 122748 43502 122760
rect 117314 122748 117320 122760
rect 117372 122748 117378 122800
rect 100018 122068 100024 122120
rect 100076 122108 100082 122120
rect 110414 122108 110420 122120
rect 100076 122080 110420 122108
rect 100076 122068 100082 122080
rect 110414 122068 110420 122080
rect 110472 122068 110478 122120
rect 37918 121388 37924 121440
rect 37976 121428 37982 121440
rect 117314 121428 117320 121440
rect 37976 121400 117320 121428
rect 37976 121388 37982 121400
rect 117314 121388 117320 121400
rect 117372 121388 117378 121440
rect 69658 120844 69664 120896
rect 69716 120884 69722 120896
rect 71682 120884 71688 120896
rect 69716 120856 71688 120884
rect 69716 120844 69722 120856
rect 71682 120844 71688 120856
rect 71740 120844 71746 120896
rect 19978 120028 19984 120080
rect 20036 120068 20042 120080
rect 117314 120068 117320 120080
rect 20036 120040 117320 120068
rect 20036 120028 20042 120040
rect 117314 120028 117320 120040
rect 117372 120028 117378 120080
rect 180242 120028 180248 120080
rect 180300 120068 180306 120080
rect 182266 120068 182272 120080
rect 180300 120040 182272 120068
rect 180300 120028 180306 120040
rect 182266 120028 182272 120040
rect 182324 120028 182330 120080
rect 110414 119960 110420 120012
rect 110472 120000 110478 120012
rect 114462 120000 114468 120012
rect 110472 119972 114468 120000
rect 110472 119960 110478 119972
rect 114462 119960 114468 119972
rect 114520 119960 114526 120012
rect 71682 119892 71688 119944
rect 71740 119932 71746 119944
rect 73154 119932 73160 119944
rect 71740 119904 73160 119932
rect 71740 119892 71746 119904
rect 73154 119892 73160 119904
rect 73212 119892 73218 119944
rect 355962 119348 355968 119400
rect 356020 119388 356026 119400
rect 366358 119388 366364 119400
rect 356020 119360 366364 119388
rect 356020 119348 356026 119360
rect 366358 119348 366364 119360
rect 366416 119348 366422 119400
rect 15838 118600 15844 118652
rect 15896 118640 15902 118652
rect 117314 118640 117320 118652
rect 15896 118612 117320 118640
rect 15896 118600 15902 118612
rect 117314 118600 117320 118612
rect 117372 118600 117378 118652
rect 104158 118532 104164 118584
rect 104216 118572 104222 118584
rect 108298 118572 108304 118584
rect 104216 118544 108304 118572
rect 104216 118532 104222 118544
rect 108298 118532 108304 118544
rect 108356 118532 108362 118584
rect 23474 117240 23480 117292
rect 23532 117280 23538 117292
rect 117314 117280 117320 117292
rect 23532 117252 117320 117280
rect 23532 117240 23538 117252
rect 117314 117240 117320 117252
rect 117372 117240 117378 117292
rect 352558 116832 352564 116884
rect 352616 116872 352622 116884
rect 355962 116872 355968 116884
rect 352616 116844 355968 116872
rect 352616 116832 352622 116844
rect 355962 116832 355968 116844
rect 356020 116832 356026 116884
rect 73154 114860 73160 114912
rect 73212 114900 73218 114912
rect 74902 114900 74908 114912
rect 73212 114872 74908 114900
rect 73212 114860 73218 114872
rect 74902 114860 74908 114872
rect 74960 114860 74966 114912
rect 114462 114452 114468 114504
rect 114520 114492 114526 114504
rect 117314 114492 117320 114504
rect 114520 114464 117320 114492
rect 114520 114452 114526 114464
rect 117314 114452 117320 114464
rect 117372 114452 117378 114504
rect 100110 113772 100116 113824
rect 100168 113812 100174 113824
rect 111794 113812 111800 113824
rect 100168 113784 111800 113812
rect 100168 113772 100174 113784
rect 111794 113772 111800 113784
rect 111852 113772 111858 113824
rect 84838 113092 84844 113144
rect 84896 113132 84902 113144
rect 117314 113132 117320 113144
rect 84896 113104 117320 113132
rect 84896 113092 84902 113104
rect 117314 113092 117320 113104
rect 117372 113092 117378 113144
rect 90358 112140 90364 112192
rect 90416 112180 90422 112192
rect 91830 112180 91836 112192
rect 90416 112152 91836 112180
rect 90416 112140 90422 112152
rect 91830 112140 91836 112152
rect 91888 112140 91894 112192
rect 74902 111800 74908 111852
rect 74960 111840 74966 111852
rect 74960 111812 75960 111840
rect 74960 111800 74966 111812
rect 3142 111732 3148 111784
rect 3200 111772 3206 111784
rect 62758 111772 62764 111784
rect 3200 111744 62764 111772
rect 3200 111732 3206 111744
rect 62758 111732 62764 111744
rect 62816 111732 62822 111784
rect 75932 111772 75960 111812
rect 180242 111800 180248 111852
rect 180300 111840 180306 111852
rect 580166 111840 580172 111852
rect 180300 111812 580172 111840
rect 180300 111800 180306 111812
rect 580166 111800 580172 111812
rect 580224 111800 580230 111852
rect 117314 111772 117320 111784
rect 75932 111744 117320 111772
rect 117314 111732 117320 111744
rect 117372 111732 117378 111784
rect 183278 111732 183284 111784
rect 183336 111772 183342 111784
rect 362218 111772 362224 111784
rect 183336 111744 362224 111772
rect 183336 111732 183342 111744
rect 362218 111732 362224 111744
rect 362276 111732 362282 111784
rect 91830 111052 91836 111104
rect 91888 111092 91894 111104
rect 97902 111092 97908 111104
rect 91888 111064 97908 111092
rect 91888 111052 91894 111064
rect 97902 111052 97908 111064
rect 97960 111052 97966 111104
rect 90450 110508 90456 110560
rect 90508 110548 90514 110560
rect 93118 110548 93124 110560
rect 90508 110520 93124 110548
rect 90508 110508 90514 110520
rect 93118 110508 93124 110520
rect 93176 110508 93182 110560
rect 349522 110440 349528 110492
rect 349580 110480 349586 110492
rect 352558 110480 352564 110492
rect 349580 110452 352564 110480
rect 349580 110440 349586 110452
rect 352558 110440 352564 110452
rect 352616 110440 352622 110492
rect 97902 110372 97908 110424
rect 97960 110412 97966 110424
rect 117314 110412 117320 110424
rect 97960 110384 117320 110412
rect 97960 110372 97966 110384
rect 117314 110372 117320 110384
rect 117372 110372 117378 110424
rect 183462 110372 183468 110424
rect 183520 110412 183526 110424
rect 367738 110412 367744 110424
rect 183520 110384 367744 110412
rect 183520 110372 183526 110384
rect 367738 110372 367744 110384
rect 367796 110372 367802 110424
rect 182266 108944 182272 108996
rect 182324 108984 182330 108996
rect 410518 108984 410524 108996
rect 182324 108956 410524 108984
rect 182324 108944 182330 108956
rect 410518 108944 410524 108956
rect 410576 108944 410582 108996
rect 108298 108264 108304 108316
rect 108356 108304 108362 108316
rect 109770 108304 109776 108316
rect 108356 108276 109776 108304
rect 108356 108264 108362 108276
rect 109770 108264 109776 108276
rect 109828 108264 109834 108316
rect 111794 106904 111800 106956
rect 111852 106944 111858 106956
rect 119430 106944 119436 106956
rect 111852 106916 119436 106944
rect 111852 106904 111858 106916
rect 119430 106904 119436 106916
rect 119488 106904 119494 106956
rect 183462 106224 183468 106276
rect 183520 106264 183526 106276
rect 409138 106264 409144 106276
rect 183520 106236 409144 106264
rect 183520 106224 183526 106236
rect 409138 106224 409144 106236
rect 409196 106224 409202 106276
rect 346394 105544 346400 105596
rect 346452 105584 346458 105596
rect 349522 105584 349528 105596
rect 346452 105556 349528 105584
rect 346452 105544 346458 105556
rect 349522 105544 349528 105556
rect 349580 105544 349586 105596
rect 109770 104796 109776 104848
rect 109828 104836 109834 104848
rect 111150 104836 111156 104848
rect 109828 104808 111156 104836
rect 109828 104796 109834 104808
rect 111150 104796 111156 104808
rect 111208 104796 111214 104848
rect 183462 104796 183468 104848
rect 183520 104836 183526 104848
rect 407758 104836 407764 104848
rect 183520 104808 407764 104836
rect 183520 104796 183526 104808
rect 407758 104796 407764 104808
rect 407816 104796 407822 104848
rect 183462 103436 183468 103488
rect 183520 103476 183526 103488
rect 406378 103476 406384 103488
rect 183520 103448 406384 103476
rect 183520 103436 183526 103448
rect 406378 103436 406384 103448
rect 406436 103436 406442 103488
rect 343634 102144 343640 102196
rect 343692 102184 343698 102196
rect 346394 102184 346400 102196
rect 343692 102156 346400 102184
rect 343692 102144 343698 102156
rect 346394 102144 346400 102156
rect 346452 102144 346458 102196
rect 182910 102076 182916 102128
rect 182968 102116 182974 102128
rect 404998 102116 405004 102128
rect 182968 102088 405004 102116
rect 182968 102076 182974 102088
rect 404998 102076 405004 102088
rect 405056 102076 405062 102128
rect 93118 101396 93124 101448
rect 93176 101436 93182 101448
rect 102134 101436 102140 101448
rect 93176 101408 102140 101436
rect 93176 101396 93182 101408
rect 102134 101396 102140 101408
rect 102192 101396 102198 101448
rect 182910 100648 182916 100700
rect 182968 100688 182974 100700
rect 403618 100688 403624 100700
rect 182968 100660 403624 100688
rect 182968 100648 182974 100660
rect 403618 100648 403624 100660
rect 403676 100648 403682 100700
rect 117958 99356 117964 99408
rect 118016 99396 118022 99408
rect 120902 99396 120908 99408
rect 118016 99368 120908 99396
rect 118016 99356 118022 99368
rect 120902 99356 120908 99368
rect 120960 99356 120966 99408
rect 180334 99356 180340 99408
rect 180392 99396 180398 99408
rect 580166 99396 580172 99408
rect 180392 99368 580172 99396
rect 180392 99356 180398 99368
rect 580166 99356 580172 99368
rect 580224 99356 580230 99408
rect 102134 99288 102140 99340
rect 102192 99328 102198 99340
rect 105538 99328 105544 99340
rect 102192 99300 105544 99328
rect 102192 99288 102198 99300
rect 105538 99288 105544 99300
rect 105596 99288 105602 99340
rect 183094 99288 183100 99340
rect 183152 99328 183158 99340
rect 400858 99328 400864 99340
rect 183152 99300 400864 99328
rect 183152 99288 183158 99300
rect 400858 99288 400864 99300
rect 400916 99288 400922 99340
rect 111150 97928 111156 97980
rect 111208 97968 111214 97980
rect 112438 97968 112444 97980
rect 111208 97940 112444 97968
rect 111208 97928 111214 97940
rect 112438 97928 112444 97940
rect 112496 97928 112502 97980
rect 183462 97928 183468 97980
rect 183520 97968 183526 97980
rect 399478 97968 399484 97980
rect 183520 97940 399484 97968
rect 183520 97928 183526 97940
rect 399478 97928 399484 97940
rect 399536 97928 399542 97980
rect 183186 96568 183192 96620
rect 183244 96608 183250 96620
rect 421558 96608 421564 96620
rect 183244 96580 421564 96608
rect 183244 96568 183250 96580
rect 421558 96568 421564 96580
rect 421616 96568 421622 96620
rect 183278 95140 183284 95192
rect 183336 95180 183342 95192
rect 418798 95180 418804 95192
rect 183336 95152 418804 95180
rect 183336 95140 183342 95152
rect 418798 95140 418804 95152
rect 418856 95140 418862 95192
rect 339218 94936 339224 94988
rect 339276 94976 339282 94988
rect 343634 94976 343640 94988
rect 339276 94948 343640 94976
rect 339276 94936 339282 94948
rect 343634 94936 343640 94948
rect 343692 94936 343698 94988
rect 183278 93780 183284 93832
rect 183336 93820 183342 93832
rect 417418 93820 417424 93832
rect 183336 93792 417424 93820
rect 183336 93780 183342 93792
rect 417418 93780 417424 93792
rect 417476 93780 417482 93832
rect 183462 92420 183468 92472
rect 183520 92460 183526 92472
rect 414658 92460 414664 92472
rect 183520 92432 414664 92460
rect 183520 92420 183526 92432
rect 414658 92420 414664 92432
rect 414716 92420 414722 92472
rect 112438 92216 112444 92268
rect 112496 92256 112502 92268
rect 113910 92256 113916 92268
rect 112496 92228 113916 92256
rect 112496 92216 112502 92228
rect 113910 92216 113916 92228
rect 113968 92216 113974 92268
rect 329098 91740 329104 91792
rect 329156 91780 329162 91792
rect 339218 91780 339224 91792
rect 329156 91752 339224 91780
rect 329156 91740 329162 91752
rect 339218 91740 339224 91752
rect 339276 91740 339282 91792
rect 182174 89632 182180 89684
rect 182232 89672 182238 89684
rect 188338 89672 188344 89684
rect 182232 89644 188344 89672
rect 182232 89632 182238 89644
rect 188338 89632 188344 89644
rect 188396 89632 188402 89684
rect 180978 88272 180984 88324
rect 181036 88312 181042 88324
rect 226978 88312 226984 88324
rect 181036 88284 226984 88312
rect 181036 88272 181042 88284
rect 226978 88272 226984 88284
rect 227036 88272 227042 88324
rect 113910 86912 113916 86964
rect 113968 86952 113974 86964
rect 116670 86952 116676 86964
rect 113968 86924 116676 86952
rect 113968 86912 113974 86924
rect 116670 86912 116676 86924
rect 116728 86912 116734 86964
rect 182174 86708 182180 86760
rect 182232 86748 182238 86760
rect 184198 86748 184204 86760
rect 182232 86720 184204 86748
rect 182232 86708 182238 86720
rect 184198 86708 184204 86720
rect 184256 86708 184262 86760
rect 105538 86232 105544 86284
rect 105596 86272 105602 86284
rect 120718 86272 120724 86284
rect 105596 86244 120724 86272
rect 105596 86232 105602 86244
rect 120718 86232 120724 86244
rect 120776 86232 120782 86284
rect 182634 85552 182640 85604
rect 182692 85592 182698 85604
rect 580166 85592 580172 85604
rect 182692 85564 580172 85592
rect 182692 85552 182698 85564
rect 580166 85552 580172 85564
rect 580224 85552 580230 85604
rect 3142 84804 3148 84856
rect 3200 84844 3206 84856
rect 3326 84844 3332 84856
rect 3200 84816 3332 84844
rect 3200 84804 3206 84816
rect 3326 84804 3332 84816
rect 3384 84804 3390 84856
rect 3418 84804 3424 84856
rect 3476 84844 3482 84856
rect 3602 84844 3608 84856
rect 3476 84816 3608 84844
rect 3476 84804 3482 84816
rect 3602 84804 3608 84816
rect 3660 84804 3666 84856
rect 3970 84736 3976 84788
rect 4028 84736 4034 84788
rect 3602 84668 3608 84720
rect 3660 84708 3666 84720
rect 3786 84708 3792 84720
rect 3660 84680 3792 84708
rect 3660 84668 3666 84680
rect 3786 84668 3792 84680
rect 3844 84668 3850 84720
rect 3786 84532 3792 84584
rect 3844 84572 3850 84584
rect 3988 84572 4016 84736
rect 3844 84544 4016 84572
rect 3844 84532 3850 84544
rect 3970 84192 3976 84244
rect 4028 84232 4034 84244
rect 120442 84232 120448 84244
rect 4028 84204 120448 84232
rect 4028 84192 4034 84204
rect 120442 84192 120448 84204
rect 120500 84192 120506 84244
rect 116670 82356 116676 82408
rect 116728 82396 116734 82408
rect 119982 82396 119988 82408
rect 116728 82368 119988 82396
rect 116728 82356 116734 82368
rect 119982 82356 119988 82368
rect 120040 82356 120046 82408
rect 182450 81404 182456 81456
rect 182508 81444 182514 81456
rect 555418 81444 555424 81456
rect 182508 81416 555424 81444
rect 182508 81404 182514 81416
rect 555418 81404 555424 81416
rect 555476 81404 555482 81456
rect 119430 80724 119436 80776
rect 119488 80764 119494 80776
rect 396810 80764 396816 80776
rect 119488 80736 158024 80764
rect 119488 80724 119494 80736
rect 5258 80656 5264 80708
rect 5316 80696 5322 80708
rect 5316 80668 151814 80696
rect 5316 80656 5322 80668
rect 151786 80560 151814 80668
rect 140746 80532 146938 80560
rect 151786 80532 154344 80560
rect 140746 80424 140774 80532
rect 139366 80396 140774 80424
rect 119982 80044 119988 80096
rect 120040 80084 120046 80096
rect 120040 80056 122834 80084
rect 120040 80044 120046 80056
rect 122806 80016 122834 80056
rect 124122 80016 124128 80028
rect 122806 79988 124128 80016
rect 124122 79976 124128 79988
rect 124180 79976 124186 80028
rect 139366 80016 139394 80396
rect 125704 79988 126054 80016
rect 125704 79756 125732 79988
rect 126026 79960 126054 79988
rect 129752 79988 130654 80016
rect 125824 79908 125830 79960
rect 125882 79908 125888 79960
rect 125916 79908 125922 79960
rect 125974 79908 125980 79960
rect 126008 79908 126014 79960
rect 126066 79908 126072 79960
rect 126376 79908 126382 79960
rect 126434 79908 126440 79960
rect 126560 79908 126566 79960
rect 126618 79908 126624 79960
rect 127756 79948 127762 79960
rect 127406 79920 127762 79948
rect 125842 79824 125870 79908
rect 125934 79880 125962 79908
rect 125934 79852 126008 79880
rect 125842 79784 125876 79824
rect 125870 79772 125876 79784
rect 125928 79772 125934 79824
rect 125686 79704 125692 79756
rect 125744 79704 125750 79756
rect 125980 79620 126008 79852
rect 5166 79568 5172 79620
rect 5224 79608 5230 79620
rect 5224 79580 115934 79608
rect 5224 79568 5230 79580
rect 115906 79404 115934 79580
rect 125962 79568 125968 79620
rect 126020 79568 126026 79620
rect 126146 79568 126152 79620
rect 126204 79608 126210 79620
rect 126394 79608 126422 79908
rect 126468 79840 126474 79892
rect 126526 79840 126532 79892
rect 126204 79580 126422 79608
rect 126204 79568 126210 79580
rect 126486 79552 126514 79840
rect 126578 79756 126606 79908
rect 126928 79880 126934 79892
rect 126900 79840 126934 79880
rect 126986 79880 126992 79892
rect 126986 79852 127033 79880
rect 126986 79840 126992 79852
rect 127112 79840 127118 79892
rect 127170 79880 127176 79892
rect 127296 79880 127302 79892
rect 127170 79840 127204 79880
rect 126578 79716 126612 79756
rect 126606 79704 126612 79716
rect 126664 79704 126670 79756
rect 126900 79552 126928 79840
rect 127176 79756 127204 79840
rect 127268 79840 127302 79880
rect 127354 79840 127360 79892
rect 127268 79756 127296 79840
rect 127158 79704 127164 79756
rect 127216 79704 127222 79756
rect 127250 79704 127256 79756
rect 127308 79704 127314 79756
rect 127406 79552 127434 79920
rect 127756 79908 127762 79920
rect 127814 79908 127820 79960
rect 128032 79908 128038 79960
rect 128090 79948 128096 79960
rect 128090 79920 128170 79948
rect 128090 79908 128096 79920
rect 127848 79840 127854 79892
rect 127906 79840 127912 79892
rect 127940 79840 127946 79892
rect 127998 79880 128004 79892
rect 127998 79840 128032 79880
rect 127866 79756 127894 79840
rect 128004 79756 128032 79840
rect 128142 79824 128170 79920
rect 128216 79908 128222 79960
rect 128274 79908 128280 79960
rect 128860 79908 128866 79960
rect 128918 79908 128924 79960
rect 128952 79908 128958 79960
rect 129010 79908 129016 79960
rect 128078 79772 128084 79824
rect 128136 79784 128170 79824
rect 128136 79772 128142 79784
rect 127866 79716 127900 79756
rect 127894 79704 127900 79716
rect 127952 79704 127958 79756
rect 127986 79704 127992 79756
rect 128044 79704 128050 79756
rect 128234 79688 128262 79908
rect 128400 79840 128406 79892
rect 128458 79840 128464 79892
rect 128584 79840 128590 79892
rect 128642 79840 128648 79892
rect 128418 79744 128446 79840
rect 128372 79716 128446 79744
rect 128234 79648 128268 79688
rect 128262 79636 128268 79648
rect 128320 79636 128326 79688
rect 128372 79620 128400 79716
rect 128602 79676 128630 79840
rect 128676 79772 128682 79824
rect 128734 79772 128740 79824
rect 128464 79648 128630 79676
rect 128694 79688 128722 79772
rect 128878 79756 128906 79908
rect 128814 79704 128820 79756
rect 128872 79716 128906 79756
rect 128872 79704 128878 79716
rect 128694 79648 128728 79688
rect 128464 79620 128492 79648
rect 128722 79636 128728 79648
rect 128780 79636 128786 79688
rect 128354 79568 128360 79620
rect 128412 79568 128418 79620
rect 128446 79568 128452 79620
rect 128504 79568 128510 79620
rect 128630 79568 128636 79620
rect 128688 79608 128694 79620
rect 128970 79608 128998 79908
rect 129596 79840 129602 79892
rect 129654 79840 129660 79892
rect 129614 79620 129642 79840
rect 129752 79620 129780 79988
rect 130626 79960 130654 79988
rect 131086 79988 133046 80016
rect 130056 79908 130062 79960
rect 130114 79908 130120 79960
rect 130332 79908 130338 79960
rect 130390 79948 130396 79960
rect 130390 79920 130562 79948
rect 130390 79908 130396 79920
rect 129872 79772 129878 79824
rect 129930 79772 129936 79824
rect 129890 79688 129918 79772
rect 130074 79756 130102 79908
rect 130240 79840 130246 79892
rect 130298 79880 130304 79892
rect 130298 79840 130332 79880
rect 130424 79840 130430 79892
rect 130482 79840 130488 79892
rect 130148 79772 130154 79824
rect 130206 79772 130212 79824
rect 130010 79704 130016 79756
rect 130068 79716 130102 79756
rect 130068 79704 130074 79716
rect 130166 79688 130194 79772
rect 130304 79756 130332 79840
rect 130442 79756 130470 79840
rect 130286 79704 130292 79756
rect 130344 79704 130350 79756
rect 130378 79704 130384 79756
rect 130436 79716 130470 79756
rect 130436 79704 130442 79716
rect 130534 79688 130562 79920
rect 130608 79908 130614 79960
rect 130666 79908 130672 79960
rect 130700 79908 130706 79960
rect 130758 79908 130764 79960
rect 130792 79908 130798 79960
rect 130850 79908 130856 79960
rect 130976 79908 130982 79960
rect 131034 79908 131040 79960
rect 130718 79688 130746 79908
rect 129826 79636 129832 79688
rect 129884 79648 129918 79688
rect 129884 79636 129890 79648
rect 130102 79636 130108 79688
rect 130160 79648 130194 79688
rect 130160 79636 130166 79648
rect 130470 79636 130476 79688
rect 130528 79648 130562 79688
rect 130528 79636 130534 79648
rect 130654 79636 130660 79688
rect 130712 79648 130746 79688
rect 130712 79636 130718 79648
rect 130810 79620 130838 79908
rect 128688 79580 128998 79608
rect 128688 79568 128694 79580
rect 129550 79568 129556 79620
rect 129608 79580 129642 79620
rect 129608 79568 129614 79580
rect 129734 79568 129740 79620
rect 129792 79568 129798 79620
rect 130746 79568 130752 79620
rect 130804 79580 130838 79620
rect 130804 79568 130810 79580
rect 130994 79552 131022 79908
rect 126422 79500 126428 79552
rect 126480 79512 126514 79552
rect 126480 79500 126486 79512
rect 126882 79500 126888 79552
rect 126940 79500 126946 79552
rect 127342 79500 127348 79552
rect 127400 79512 127434 79552
rect 127820 79512 128032 79540
rect 127400 79500 127406 79512
rect 116578 79432 116584 79484
rect 116636 79472 116642 79484
rect 127820 79472 127848 79512
rect 116636 79444 127848 79472
rect 116636 79432 116642 79444
rect 127894 79432 127900 79484
rect 127952 79432 127958 79484
rect 128004 79472 128032 79512
rect 130930 79500 130936 79552
rect 130988 79512 131022 79552
rect 130988 79500 130994 79512
rect 128004 79444 129412 79472
rect 115906 79376 118832 79404
rect 3326 79296 3332 79348
rect 3384 79336 3390 79348
rect 118804 79336 118832 79376
rect 127434 79364 127440 79416
rect 127492 79404 127498 79416
rect 127912 79404 127940 79432
rect 127492 79376 127940 79404
rect 127492 79364 127498 79376
rect 3384 79308 118694 79336
rect 118804 79308 125594 79336
rect 3384 79296 3390 79308
rect 118666 79132 118694 79308
rect 125566 79268 125594 79308
rect 127618 79296 127624 79348
rect 127676 79336 127682 79348
rect 127894 79336 127900 79348
rect 127676 79308 127900 79336
rect 127676 79296 127682 79308
rect 127894 79296 127900 79308
rect 127952 79296 127958 79348
rect 129384 79336 129412 79444
rect 129458 79432 129464 79484
rect 129516 79472 129522 79484
rect 131086 79472 131114 79988
rect 133018 79960 133046 79988
rect 133110 79988 133506 80016
rect 131344 79908 131350 79960
rect 131402 79908 131408 79960
rect 131528 79908 131534 79960
rect 131586 79908 131592 79960
rect 132632 79908 132638 79960
rect 132690 79908 132696 79960
rect 133000 79908 133006 79960
rect 133058 79908 133064 79960
rect 131160 79840 131166 79892
rect 131218 79840 131224 79892
rect 131252 79840 131258 79892
rect 131310 79840 131316 79892
rect 131178 79552 131206 79840
rect 131270 79620 131298 79840
rect 131362 79824 131390 79908
rect 131344 79772 131350 79824
rect 131402 79772 131408 79824
rect 131270 79580 131304 79620
rect 131298 79568 131304 79580
rect 131356 79568 131362 79620
rect 131546 79552 131574 79908
rect 131988 79840 131994 79892
rect 132046 79840 132052 79892
rect 132650 79880 132678 79908
rect 132650 79852 132724 79880
rect 131804 79772 131810 79824
rect 131862 79772 131868 79824
rect 131822 79688 131850 79772
rect 132006 79756 132034 79840
rect 132172 79772 132178 79824
rect 132230 79772 132236 79824
rect 132448 79772 132454 79824
rect 132506 79772 132512 79824
rect 131942 79704 131948 79756
rect 132000 79716 132034 79756
rect 132190 79744 132218 79772
rect 132144 79716 132218 79744
rect 132000 79704 132006 79716
rect 131822 79648 131856 79688
rect 131850 79636 131856 79648
rect 131908 79636 131914 79688
rect 132144 79620 132172 79716
rect 132126 79568 132132 79620
rect 132184 79568 132190 79620
rect 132466 79552 132494 79772
rect 132696 79756 132724 79852
rect 132678 79704 132684 79756
rect 132736 79704 132742 79756
rect 132954 79704 132960 79756
rect 133012 79704 133018 79756
rect 132586 79636 132592 79688
rect 132644 79676 132650 79688
rect 132972 79676 133000 79704
rect 132644 79648 133000 79676
rect 132644 79636 132650 79648
rect 133110 79608 133138 79988
rect 133478 79960 133506 79988
rect 136882 79988 137508 80016
rect 133460 79908 133466 79960
rect 133518 79908 133524 79960
rect 133828 79908 133834 79960
rect 133886 79908 133892 79960
rect 134104 79908 134110 79960
rect 134162 79908 134168 79960
rect 134196 79908 134202 79960
rect 134254 79908 134260 79960
rect 134564 79948 134570 79960
rect 134490 79920 134570 79948
rect 133276 79840 133282 79892
rect 133334 79880 133340 79892
rect 133846 79880 133874 79908
rect 133334 79840 133368 79880
rect 133184 79772 133190 79824
rect 133242 79812 133248 79824
rect 133242 79772 133276 79812
rect 133248 79620 133276 79772
rect 131178 79512 131212 79552
rect 131206 79500 131212 79512
rect 131264 79500 131270 79552
rect 131482 79500 131488 79552
rect 131540 79512 131574 79552
rect 131540 79500 131546 79512
rect 132402 79500 132408 79552
rect 132460 79512 132494 79552
rect 132972 79580 133138 79608
rect 132460 79500 132466 79512
rect 129516 79444 131114 79472
rect 132972 79472 133000 79580
rect 133230 79568 133236 79620
rect 133288 79568 133294 79620
rect 133046 79500 133052 79552
rect 133104 79540 133110 79552
rect 133340 79540 133368 79840
rect 133800 79852 133874 79880
rect 133552 79812 133558 79824
rect 133478 79784 133558 79812
rect 133478 79608 133506 79784
rect 133552 79772 133558 79784
rect 133610 79772 133616 79824
rect 133644 79772 133650 79824
rect 133702 79772 133708 79824
rect 133662 79688 133690 79772
rect 133800 79756 133828 79852
rect 133920 79840 133926 79892
rect 133978 79840 133984 79892
rect 133938 79812 133966 79840
rect 133892 79784 133966 79812
rect 133892 79756 133920 79784
rect 133782 79704 133788 79756
rect 133840 79704 133846 79756
rect 133874 79704 133880 79756
rect 133932 79704 133938 79756
rect 133966 79704 133972 79756
rect 134024 79744 134030 79756
rect 134122 79744 134150 79908
rect 134214 79824 134242 79908
rect 134380 79840 134386 79892
rect 134438 79840 134444 79892
rect 134214 79784 134248 79824
rect 134242 79772 134248 79784
rect 134300 79772 134306 79824
rect 134024 79716 134150 79744
rect 134024 79704 134030 79716
rect 133598 79636 133604 79688
rect 133656 79648 133690 79688
rect 133656 79636 133662 79648
rect 134398 79620 134426 79840
rect 133432 79580 133506 79608
rect 133432 79552 133460 79580
rect 134334 79568 134340 79620
rect 134392 79580 134426 79620
rect 134392 79568 134398 79580
rect 133104 79512 133368 79540
rect 133104 79500 133110 79512
rect 133414 79500 133420 79552
rect 133472 79500 133478 79552
rect 134058 79500 134064 79552
rect 134116 79540 134122 79552
rect 134490 79540 134518 79920
rect 134564 79908 134570 79920
rect 134622 79908 134628 79960
rect 134840 79908 134846 79960
rect 134898 79908 134904 79960
rect 135024 79908 135030 79960
rect 135082 79908 135088 79960
rect 135116 79908 135122 79960
rect 135174 79908 135180 79960
rect 135576 79948 135582 79960
rect 135548 79908 135582 79948
rect 135634 79908 135640 79960
rect 135668 79908 135674 79960
rect 135726 79908 135732 79960
rect 136036 79908 136042 79960
rect 136094 79908 136100 79960
rect 136128 79908 136134 79960
rect 136186 79908 136192 79960
rect 136220 79908 136226 79960
rect 136278 79908 136284 79960
rect 136312 79908 136318 79960
rect 136370 79908 136376 79960
rect 136496 79908 136502 79960
rect 136554 79908 136560 79960
rect 136772 79948 136778 79960
rect 136652 79920 136778 79948
rect 134656 79880 134662 79892
rect 134628 79840 134662 79880
rect 134714 79840 134720 79892
rect 134748 79840 134754 79892
rect 134806 79840 134812 79892
rect 134628 79756 134656 79840
rect 134766 79812 134794 79840
rect 134720 79784 134794 79812
rect 134720 79756 134748 79784
rect 134858 79756 134886 79908
rect 134610 79704 134616 79756
rect 134668 79704 134674 79756
rect 134702 79704 134708 79756
rect 134760 79704 134766 79756
rect 134794 79704 134800 79756
rect 134852 79716 134886 79756
rect 135042 79744 135070 79908
rect 134996 79716 135070 79744
rect 134852 79704 134858 79716
rect 134996 79688 135024 79716
rect 135134 79688 135162 79908
rect 135548 79688 135576 79908
rect 135686 79880 135714 79908
rect 135944 79880 135950 79892
rect 135640 79852 135714 79880
rect 134978 79636 134984 79688
rect 135036 79636 135042 79688
rect 135070 79636 135076 79688
rect 135128 79648 135162 79688
rect 135128 79636 135134 79648
rect 135530 79636 135536 79688
rect 135588 79636 135594 79688
rect 134116 79512 134518 79540
rect 134116 79500 134122 79512
rect 133230 79472 133236 79484
rect 132972 79444 133236 79472
rect 129516 79432 129522 79444
rect 133230 79432 133236 79444
rect 133288 79432 133294 79484
rect 135640 79472 135668 79852
rect 135916 79840 135950 79880
rect 136002 79840 136008 79892
rect 135760 79772 135766 79824
rect 135818 79772 135824 79824
rect 135778 79688 135806 79772
rect 135714 79636 135720 79688
rect 135772 79648 135806 79688
rect 135772 79636 135778 79648
rect 135916 79620 135944 79840
rect 136054 79812 136082 79908
rect 136008 79784 136082 79812
rect 136008 79756 136036 79784
rect 136146 79756 136174 79908
rect 135990 79704 135996 79756
rect 136048 79704 136054 79756
rect 136082 79704 136088 79756
rect 136140 79716 136174 79756
rect 136140 79704 136146 79716
rect 135898 79568 135904 79620
rect 135956 79568 135962 79620
rect 135806 79500 135812 79552
rect 135864 79540 135870 79552
rect 136238 79540 136266 79908
rect 136330 79620 136358 79908
rect 136514 79824 136542 79908
rect 136450 79772 136456 79824
rect 136508 79784 136542 79824
rect 136508 79772 136514 79784
rect 136652 79620 136680 79920
rect 136772 79908 136778 79920
rect 136830 79908 136836 79960
rect 136882 79892 136910 79988
rect 137140 79908 137146 79960
rect 137198 79908 137204 79960
rect 137232 79908 137238 79960
rect 137290 79908 137296 79960
rect 136864 79840 136870 79892
rect 136922 79840 136928 79892
rect 137158 79824 137186 79908
rect 136956 79772 136962 79824
rect 137014 79772 137020 79824
rect 137094 79772 137100 79824
rect 137152 79784 137186 79824
rect 137152 79772 137158 79784
rect 136974 79744 137002 79772
rect 136928 79716 137002 79744
rect 136928 79688 136956 79716
rect 136910 79636 136916 79688
rect 136968 79636 136974 79688
rect 137002 79636 137008 79688
rect 137060 79676 137066 79688
rect 137250 79676 137278 79908
rect 137324 79840 137330 79892
rect 137382 79880 137388 79892
rect 137382 79840 137416 79880
rect 137060 79648 137278 79676
rect 137060 79636 137066 79648
rect 137388 79620 137416 79840
rect 137480 79620 137508 79988
rect 139044 79988 139394 80016
rect 140378 79988 142154 80016
rect 138060 79908 138066 79960
rect 138118 79908 138124 79960
rect 138152 79908 138158 79960
rect 138210 79908 138216 79960
rect 138428 79908 138434 79960
rect 138486 79908 138492 79960
rect 138704 79908 138710 79960
rect 138762 79908 138768 79960
rect 138796 79908 138802 79960
rect 138854 79908 138860 79960
rect 138888 79908 138894 79960
rect 138946 79948 138952 79960
rect 138946 79908 138980 79948
rect 137600 79840 137606 79892
rect 137658 79840 137664 79892
rect 137968 79880 137974 79892
rect 137802 79852 137974 79880
rect 136330 79580 136364 79620
rect 136358 79568 136364 79580
rect 136416 79568 136422 79620
rect 136634 79568 136640 79620
rect 136692 79568 136698 79620
rect 137370 79568 137376 79620
rect 137428 79568 137434 79620
rect 137462 79568 137468 79620
rect 137520 79568 137526 79620
rect 137618 79540 137646 79840
rect 135864 79512 136266 79540
rect 136744 79512 137646 79540
rect 135864 79500 135870 79512
rect 136744 79484 136772 79512
rect 137802 79484 137830 79852
rect 137968 79840 137974 79852
rect 138026 79840 138032 79892
rect 137876 79772 137882 79824
rect 137934 79772 137940 79824
rect 137894 79552 137922 79772
rect 138078 79552 138106 79908
rect 138170 79608 138198 79908
rect 138336 79840 138342 79892
rect 138394 79840 138400 79892
rect 138354 79812 138382 79840
rect 138308 79784 138382 79812
rect 138308 79676 138336 79784
rect 138446 79756 138474 79908
rect 138382 79704 138388 79756
rect 138440 79716 138474 79756
rect 138440 79704 138446 79716
rect 138308 79648 138428 79676
rect 138290 79608 138296 79620
rect 138170 79580 138296 79608
rect 138290 79568 138296 79580
rect 138348 79568 138354 79620
rect 137894 79512 137928 79552
rect 137922 79500 137928 79512
rect 137980 79500 137986 79552
rect 138014 79500 138020 79552
rect 138072 79512 138106 79552
rect 138072 79500 138078 79512
rect 134950 79444 135668 79472
rect 134950 79416 134978 79444
rect 136726 79432 136732 79484
rect 136784 79432 136790 79484
rect 137278 79432 137284 79484
rect 137336 79472 137342 79484
rect 137646 79472 137652 79484
rect 137336 79444 137652 79472
rect 137336 79432 137342 79444
rect 137646 79432 137652 79444
rect 137704 79432 137710 79484
rect 137802 79444 137836 79484
rect 137830 79432 137836 79444
rect 137888 79432 137894 79484
rect 138106 79432 138112 79484
rect 138164 79472 138170 79484
rect 138400 79472 138428 79648
rect 138566 79636 138572 79688
rect 138624 79676 138630 79688
rect 138722 79676 138750 79908
rect 138624 79648 138750 79676
rect 138624 79636 138630 79648
rect 138814 79620 138842 79908
rect 138814 79580 138848 79620
rect 138842 79568 138848 79580
rect 138900 79568 138906 79620
rect 138658 79500 138664 79552
rect 138716 79540 138722 79552
rect 138952 79540 138980 79908
rect 139044 79688 139072 79988
rect 140378 79960 140406 79988
rect 139164 79948 139170 79960
rect 139136 79908 139170 79948
rect 139222 79908 139228 79960
rect 139256 79908 139262 79960
rect 139314 79908 139320 79960
rect 139808 79948 139814 79960
rect 139596 79920 139814 79948
rect 139136 79688 139164 79908
rect 139274 79824 139302 79908
rect 139440 79840 139446 79892
rect 139498 79840 139504 79892
rect 139210 79772 139216 79824
rect 139268 79784 139302 79824
rect 139268 79772 139274 79784
rect 139026 79636 139032 79688
rect 139084 79636 139090 79688
rect 139118 79636 139124 79688
rect 139176 79636 139182 79688
rect 139458 79620 139486 79840
rect 139394 79568 139400 79620
rect 139452 79580 139486 79620
rect 139452 79568 139458 79580
rect 139596 79552 139624 79920
rect 139808 79908 139814 79920
rect 139866 79908 139872 79960
rect 140176 79908 140182 79960
rect 140234 79908 140240 79960
rect 140268 79908 140274 79960
rect 140326 79908 140332 79960
rect 140360 79908 140366 79960
rect 140418 79908 140424 79960
rect 140820 79948 140826 79960
rect 140792 79908 140826 79948
rect 140878 79908 140884 79960
rect 140912 79908 140918 79960
rect 140970 79908 140976 79960
rect 141372 79908 141378 79960
rect 141430 79908 141436 79960
rect 141464 79908 141470 79960
rect 141522 79908 141528 79960
rect 141556 79908 141562 79960
rect 141614 79908 141620 79960
rect 141924 79948 141930 79960
rect 141896 79908 141930 79948
rect 141982 79908 141988 79960
rect 139900 79880 139906 79892
rect 139872 79840 139906 79880
rect 139958 79840 139964 79892
rect 139872 79756 139900 79840
rect 139992 79812 139998 79824
rect 139964 79772 139998 79812
rect 140050 79772 140056 79824
rect 139854 79704 139860 79756
rect 139912 79704 139918 79756
rect 139964 79688 139992 79772
rect 139946 79636 139952 79688
rect 140004 79636 140010 79688
rect 140194 79608 140222 79908
rect 140286 79676 140314 79908
rect 140636 79840 140642 79892
rect 140694 79840 140700 79892
rect 140654 79744 140682 79840
rect 140516 79716 140682 79744
rect 140406 79676 140412 79688
rect 140286 79648 140412 79676
rect 140406 79636 140412 79648
rect 140464 79636 140470 79688
rect 140194 79580 140268 79608
rect 138716 79512 138980 79540
rect 138716 79500 138722 79512
rect 139578 79500 139584 79552
rect 139636 79500 139642 79552
rect 138164 79444 138428 79472
rect 140240 79472 140268 79580
rect 140314 79568 140320 79620
rect 140372 79608 140378 79620
rect 140516 79608 140544 79716
rect 140682 79636 140688 79688
rect 140740 79676 140746 79688
rect 140792 79676 140820 79908
rect 140930 79688 140958 79908
rect 141188 79840 141194 79892
rect 141246 79840 141252 79892
rect 141096 79772 141102 79824
rect 141154 79772 141160 79824
rect 141114 79688 141142 79772
rect 140740 79648 140820 79676
rect 140740 79636 140746 79648
rect 140866 79636 140872 79688
rect 140924 79648 140958 79688
rect 140924 79636 140930 79648
rect 141050 79636 141056 79688
rect 141108 79648 141142 79688
rect 141108 79636 141114 79648
rect 140372 79580 140544 79608
rect 140372 79568 140378 79580
rect 140774 79568 140780 79620
rect 140832 79608 140838 79620
rect 141206 79608 141234 79840
rect 141390 79688 141418 79908
rect 141326 79636 141332 79688
rect 141384 79648 141418 79688
rect 141384 79636 141390 79648
rect 140832 79580 141234 79608
rect 141482 79620 141510 79908
rect 141574 79688 141602 79908
rect 141740 79840 141746 79892
rect 141798 79880 141804 79892
rect 141798 79840 141832 79880
rect 141804 79756 141832 79840
rect 141786 79704 141792 79756
rect 141844 79704 141850 79756
rect 141574 79648 141608 79688
rect 141602 79636 141608 79648
rect 141660 79636 141666 79688
rect 141896 79620 141924 79908
rect 142016 79840 142022 79892
rect 142074 79840 142080 79892
rect 141482 79580 141516 79620
rect 140832 79568 140838 79580
rect 141510 79568 141516 79580
rect 141568 79568 141574 79620
rect 141878 79568 141884 79620
rect 141936 79568 141942 79620
rect 140314 79472 140320 79484
rect 140240 79444 140320 79472
rect 138164 79432 138170 79444
rect 140314 79432 140320 79444
rect 140372 79432 140378 79484
rect 131114 79364 131120 79416
rect 131172 79404 131178 79416
rect 131172 79376 131804 79404
rect 131172 79364 131178 79376
rect 131776 79336 131804 79376
rect 132862 79364 132868 79416
rect 132920 79404 132926 79416
rect 133138 79404 133144 79416
rect 132920 79376 133144 79404
rect 132920 79364 132926 79376
rect 133138 79364 133144 79376
rect 133196 79364 133202 79416
rect 134886 79364 134892 79416
rect 134944 79376 134978 79416
rect 140498 79404 140504 79416
rect 135226 79376 140504 79404
rect 134944 79364 134950 79376
rect 135226 79336 135254 79376
rect 140498 79364 140504 79376
rect 140556 79364 140562 79416
rect 129384 79308 131252 79336
rect 131776 79308 135254 79336
rect 131114 79268 131120 79280
rect 125566 79240 131120 79268
rect 131114 79228 131120 79240
rect 131172 79228 131178 79280
rect 131224 79268 131252 79308
rect 141326 79296 141332 79348
rect 141384 79336 141390 79348
rect 141694 79336 141700 79348
rect 141384 79308 141700 79336
rect 141384 79296 141390 79308
rect 141694 79296 141700 79308
rect 141752 79296 141758 79348
rect 142034 79336 142062 79840
rect 142126 79540 142154 79988
rect 142218 79988 146202 80016
rect 142218 79960 142246 79988
rect 142200 79908 142206 79960
rect 142258 79908 142264 79960
rect 142292 79908 142298 79960
rect 142350 79908 142356 79960
rect 142476 79908 142482 79960
rect 142534 79908 142540 79960
rect 143212 79908 143218 79960
rect 143270 79908 143276 79960
rect 143304 79908 143310 79960
rect 143362 79908 143368 79960
rect 143488 79908 143494 79960
rect 143546 79908 143552 79960
rect 143580 79908 143586 79960
rect 143638 79908 143644 79960
rect 144224 79908 144230 79960
rect 144282 79908 144288 79960
rect 144500 79908 144506 79960
rect 144558 79908 144564 79960
rect 144592 79908 144598 79960
rect 144650 79948 144656 79960
rect 145328 79948 145334 79960
rect 144650 79908 144684 79948
rect 142310 79756 142338 79908
rect 142246 79704 142252 79756
rect 142304 79716 142338 79756
rect 142304 79704 142310 79716
rect 142494 79688 142522 79908
rect 142660 79840 142666 79892
rect 142718 79840 142724 79892
rect 142844 79840 142850 79892
rect 142902 79840 142908 79892
rect 142430 79636 142436 79688
rect 142488 79648 142522 79688
rect 142488 79636 142494 79648
rect 142678 79608 142706 79840
rect 142862 79688 142890 79840
rect 142936 79772 142942 79824
rect 142994 79772 143000 79824
rect 142954 79744 142982 79772
rect 142954 79716 143028 79744
rect 142862 79648 142896 79688
rect 142890 79636 142896 79648
rect 142948 79636 142954 79688
rect 142798 79608 142804 79620
rect 142678 79580 142804 79608
rect 142798 79568 142804 79580
rect 142856 79568 142862 79620
rect 143000 79552 143028 79716
rect 143230 79688 143258 79908
rect 143322 79824 143350 79908
rect 143322 79784 143356 79824
rect 143350 79772 143356 79784
rect 143408 79772 143414 79824
rect 143506 79812 143534 79908
rect 143460 79784 143534 79812
rect 143460 79744 143488 79784
rect 143368 79716 143488 79744
rect 143230 79648 143264 79688
rect 143258 79636 143264 79648
rect 143316 79636 143322 79688
rect 143368 79608 143396 79716
rect 143442 79636 143448 79688
rect 143500 79676 143506 79688
rect 143598 79676 143626 79908
rect 143672 79840 143678 79892
rect 143730 79840 143736 79892
rect 143500 79648 143626 79676
rect 143500 79636 143506 79648
rect 143534 79608 143540 79620
rect 143368 79580 143540 79608
rect 143534 79568 143540 79580
rect 143592 79568 143598 79620
rect 142126 79512 142936 79540
rect 142908 79472 142936 79512
rect 142982 79500 142988 79552
rect 143040 79500 143046 79552
rect 143690 79540 143718 79840
rect 143948 79772 143954 79824
rect 144006 79772 144012 79824
rect 143966 79744 143994 79772
rect 143828 79716 143994 79744
rect 143690 79512 143764 79540
rect 143626 79472 143632 79484
rect 142908 79444 143632 79472
rect 143626 79432 143632 79444
rect 143684 79432 143690 79484
rect 142154 79336 142160 79348
rect 142034 79308 142160 79336
rect 142154 79296 142160 79308
rect 142212 79296 142218 79348
rect 143736 79336 143764 79512
rect 143828 79484 143856 79716
rect 143902 79636 143908 79688
rect 143960 79636 143966 79688
rect 143920 79608 143948 79636
rect 144242 79620 144270 79908
rect 144408 79840 144414 79892
rect 144466 79840 144472 79892
rect 144426 79688 144454 79840
rect 144518 79744 144546 79908
rect 144518 79716 144592 79744
rect 144564 79688 144592 79716
rect 144426 79648 144460 79688
rect 144454 79636 144460 79648
rect 144512 79636 144518 79688
rect 144546 79636 144552 79688
rect 144604 79636 144610 79688
rect 143920 79580 144132 79608
rect 144242 79580 144276 79620
rect 144104 79552 144132 79580
rect 144270 79568 144276 79580
rect 144328 79568 144334 79620
rect 144086 79500 144092 79552
rect 144144 79500 144150 79552
rect 143810 79432 143816 79484
rect 143868 79432 143874 79484
rect 144656 79472 144684 79908
rect 144748 79920 145334 79948
rect 144748 79552 144776 79920
rect 145328 79908 145334 79920
rect 145386 79908 145392 79960
rect 145604 79908 145610 79960
rect 145662 79908 145668 79960
rect 144960 79840 144966 79892
rect 145018 79840 145024 79892
rect 145144 79840 145150 79892
rect 145202 79840 145208 79892
rect 144978 79756 145006 79840
rect 144914 79704 144920 79756
rect 144972 79716 145006 79756
rect 145162 79744 145190 79840
rect 145116 79716 145190 79744
rect 144972 79704 144978 79716
rect 145116 79688 145144 79716
rect 145098 79636 145104 79688
rect 145156 79636 145162 79688
rect 144730 79500 144736 79552
rect 144788 79500 144794 79552
rect 145282 79500 145288 79552
rect 145340 79540 145346 79552
rect 145622 79540 145650 79908
rect 146174 79620 146202 79988
rect 146248 79908 146254 79960
rect 146306 79908 146312 79960
rect 146432 79948 146438 79960
rect 146358 79920 146438 79948
rect 146266 79688 146294 79908
rect 146358 79756 146386 79920
rect 146432 79908 146438 79920
rect 146490 79908 146496 79960
rect 146616 79908 146622 79960
rect 146674 79908 146680 79960
rect 146524 79880 146530 79892
rect 146496 79840 146530 79880
rect 146582 79840 146588 79892
rect 146496 79756 146524 79840
rect 146358 79716 146392 79756
rect 146386 79704 146392 79716
rect 146444 79704 146450 79756
rect 146478 79704 146484 79756
rect 146536 79704 146542 79756
rect 146266 79648 146300 79688
rect 146294 79636 146300 79648
rect 146352 79636 146358 79688
rect 146174 79580 146208 79620
rect 146202 79568 146208 79580
rect 146260 79568 146266 79620
rect 145340 79512 145650 79540
rect 146634 79552 146662 79908
rect 146800 79840 146806 79892
rect 146858 79840 146864 79892
rect 146634 79512 146668 79552
rect 145340 79500 145346 79512
rect 146662 79500 146668 79512
rect 146720 79500 146726 79552
rect 146202 79472 146208 79484
rect 144656 79444 146208 79472
rect 146202 79432 146208 79444
rect 146260 79432 146266 79484
rect 146386 79432 146392 79484
rect 146444 79472 146450 79484
rect 146818 79472 146846 79840
rect 146910 79552 146938 80532
rect 149118 80464 151814 80492
rect 149118 79960 149146 80464
rect 151786 80424 151814 80464
rect 151786 80396 152366 80424
rect 150866 79988 151400 80016
rect 150866 79960 150894 79988
rect 147260 79948 147266 79960
rect 147232 79908 147266 79948
rect 147318 79908 147324 79960
rect 147444 79908 147450 79960
rect 147502 79908 147508 79960
rect 147536 79908 147542 79960
rect 147594 79908 147600 79960
rect 147628 79908 147634 79960
rect 147686 79908 147692 79960
rect 147720 79908 147726 79960
rect 147778 79908 147784 79960
rect 147904 79908 147910 79960
rect 147962 79908 147968 79960
rect 147996 79908 148002 79960
rect 148054 79908 148060 79960
rect 148088 79908 148094 79960
rect 148146 79908 148152 79960
rect 148364 79908 148370 79960
rect 148422 79908 148428 79960
rect 148456 79908 148462 79960
rect 148514 79908 148520 79960
rect 148732 79908 148738 79960
rect 148790 79948 148796 79960
rect 148790 79908 148824 79948
rect 149100 79908 149106 79960
rect 149158 79908 149164 79960
rect 149468 79948 149474 79960
rect 149210 79920 149474 79948
rect 146984 79840 146990 79892
rect 147042 79840 147048 79892
rect 147002 79620 147030 79840
rect 147002 79580 147036 79620
rect 147030 79568 147036 79580
rect 147088 79568 147094 79620
rect 147232 79608 147260 79908
rect 147352 79880 147358 79892
rect 147324 79840 147358 79880
rect 147410 79840 147416 79892
rect 147324 79756 147352 79840
rect 147462 79812 147490 79908
rect 147416 79784 147490 79812
rect 147416 79756 147444 79784
rect 147306 79704 147312 79756
rect 147364 79704 147370 79756
rect 147398 79704 147404 79756
rect 147456 79704 147462 79756
rect 147554 79688 147582 79908
rect 147490 79636 147496 79688
rect 147548 79648 147582 79688
rect 147548 79636 147554 79648
rect 147646 79620 147674 79908
rect 147232 79580 147352 79608
rect 146910 79512 146944 79552
rect 146938 79500 146944 79512
rect 146996 79500 147002 79552
rect 146444 79444 146846 79472
rect 146444 79432 146450 79444
rect 147122 79432 147128 79484
rect 147180 79472 147186 79484
rect 147324 79472 147352 79580
rect 147582 79568 147588 79620
rect 147640 79580 147674 79620
rect 147640 79568 147646 79580
rect 147738 79540 147766 79908
rect 147922 79880 147950 79908
rect 147876 79852 147950 79880
rect 147876 79756 147904 79852
rect 148014 79812 148042 79908
rect 147968 79784 148042 79812
rect 147968 79756 147996 79784
rect 148106 79756 148134 79908
rect 147858 79704 147864 79756
rect 147916 79704 147922 79756
rect 147950 79704 147956 79756
rect 148008 79704 148014 79756
rect 148042 79704 148048 79756
rect 148100 79716 148134 79756
rect 148100 79704 148106 79716
rect 148382 79620 148410 79908
rect 148318 79568 148324 79620
rect 148376 79580 148410 79620
rect 148474 79608 148502 79908
rect 148796 79620 148824 79908
rect 149210 79812 149238 79920
rect 149468 79908 149474 79920
rect 149526 79908 149532 79960
rect 149652 79908 149658 79960
rect 149710 79908 149716 79960
rect 149744 79908 149750 79960
rect 149802 79908 149808 79960
rect 150020 79948 150026 79960
rect 149854 79920 150026 79948
rect 149284 79840 149290 79892
rect 149342 79880 149348 79892
rect 149670 79880 149698 79908
rect 149342 79852 149468 79880
rect 149342 79840 149348 79852
rect 149210 79784 149376 79812
rect 149348 79688 149376 79784
rect 149330 79636 149336 79688
rect 149388 79636 149394 79688
rect 149440 79620 149468 79852
rect 149624 79852 149698 79880
rect 149624 79688 149652 79852
rect 149762 79824 149790 79908
rect 149698 79772 149704 79824
rect 149756 79784 149790 79824
rect 149756 79772 149762 79784
rect 149606 79636 149612 79688
rect 149664 79636 149670 79688
rect 148594 79608 148600 79620
rect 148474 79580 148600 79608
rect 148376 79568 148382 79580
rect 148594 79568 148600 79580
rect 148652 79568 148658 79620
rect 148778 79568 148784 79620
rect 148836 79568 148842 79620
rect 149422 79568 149428 79620
rect 149480 79568 149486 79620
rect 149854 79608 149882 79920
rect 150020 79908 150026 79920
rect 150078 79908 150084 79960
rect 150848 79908 150854 79960
rect 150906 79908 150912 79960
rect 151032 79908 151038 79960
rect 151090 79908 151096 79960
rect 149928 79840 149934 79892
rect 149986 79840 149992 79892
rect 150388 79840 150394 79892
rect 150446 79880 150452 79892
rect 150446 79852 150572 79880
rect 150446 79840 150452 79852
rect 149946 79676 149974 79840
rect 150342 79676 150348 79688
rect 149946 79648 150348 79676
rect 150342 79636 150348 79648
rect 150400 79636 150406 79688
rect 150544 79620 150572 79852
rect 150710 79636 150716 79688
rect 150768 79676 150774 79688
rect 151050 79676 151078 79908
rect 151216 79840 151222 79892
rect 151274 79840 151280 79892
rect 151234 79688 151262 79840
rect 150768 79648 151078 79676
rect 150768 79636 150774 79648
rect 151170 79636 151176 79688
rect 151228 79648 151262 79688
rect 151228 79636 151234 79648
rect 151372 79620 151400 79988
rect 151584 79908 151590 79960
rect 151642 79908 151648 79960
rect 152228 79948 152234 79960
rect 151832 79920 152234 79948
rect 151492 79840 151498 79892
rect 151550 79840 151556 79892
rect 149974 79608 149980 79620
rect 149854 79580 149980 79608
rect 149974 79568 149980 79580
rect 150032 79568 150038 79620
rect 150526 79568 150532 79620
rect 150584 79568 150590 79620
rect 151354 79568 151360 79620
rect 151412 79568 151418 79620
rect 150066 79540 150072 79552
rect 147738 79512 150072 79540
rect 150066 79500 150072 79512
rect 150124 79500 150130 79552
rect 147180 79444 147352 79472
rect 147180 79432 147186 79444
rect 147674 79432 147680 79484
rect 147732 79472 147738 79484
rect 151510 79472 151538 79840
rect 151602 79552 151630 79908
rect 151676 79840 151682 79892
rect 151734 79880 151740 79892
rect 151734 79840 151768 79880
rect 151740 79620 151768 79840
rect 151832 79620 151860 79920
rect 152228 79908 152234 79920
rect 152286 79908 152292 79960
rect 152044 79840 152050 79892
rect 152102 79840 152108 79892
rect 151722 79568 151728 79620
rect 151780 79568 151786 79620
rect 151814 79568 151820 79620
rect 151872 79568 151878 79620
rect 152062 79608 152090 79840
rect 152338 79744 152366 80396
rect 152688 79908 152694 79960
rect 152746 79908 152752 79960
rect 152872 79948 152878 79960
rect 152844 79908 152878 79948
rect 152930 79908 152936 79960
rect 152964 79908 152970 79960
rect 153022 79908 153028 79960
rect 153056 79908 153062 79960
rect 153114 79908 153120 79960
rect 153240 79908 153246 79960
rect 153298 79908 153304 79960
rect 152706 79824 152734 79908
rect 152642 79772 152648 79824
rect 152700 79784 152734 79824
rect 152700 79772 152706 79784
rect 152734 79744 152740 79756
rect 152338 79716 152740 79744
rect 152734 79704 152740 79716
rect 152792 79704 152798 79756
rect 152844 79688 152872 79908
rect 152982 79880 153010 79908
rect 152936 79852 153010 79880
rect 152936 79744 152964 79852
rect 153074 79824 153102 79908
rect 153010 79772 153016 79824
rect 153068 79784 153102 79824
rect 153068 79772 153074 79784
rect 152936 79716 153056 79744
rect 152826 79636 152832 79688
rect 152884 79636 152890 79688
rect 152918 79608 152924 79620
rect 152062 79580 152924 79608
rect 152918 79568 152924 79580
rect 152976 79568 152982 79620
rect 151602 79512 151636 79552
rect 151630 79500 151636 79512
rect 151688 79500 151694 79552
rect 147732 79444 151538 79472
rect 153028 79472 153056 79716
rect 153258 79608 153286 79908
rect 153608 79840 153614 79892
rect 153666 79880 153672 79892
rect 153666 79852 154022 79880
rect 153666 79840 153672 79852
rect 153562 79608 153568 79620
rect 153258 79580 153568 79608
rect 153562 79568 153568 79580
rect 153620 79568 153626 79620
rect 153994 79608 154022 79852
rect 153994 79580 154068 79608
rect 154040 79540 154068 79580
rect 154114 79540 154120 79552
rect 154040 79512 154120 79540
rect 154114 79500 154120 79512
rect 154172 79500 154178 79552
rect 153378 79472 153384 79484
rect 153028 79444 153384 79472
rect 147732 79432 147738 79444
rect 153378 79432 153384 79444
rect 153436 79432 153442 79484
rect 154316 79472 154344 80532
rect 154804 79908 154810 79960
rect 154862 79948 154868 79960
rect 156184 79948 156190 79960
rect 154862 79920 155724 79948
rect 154862 79908 154868 79920
rect 155356 79840 155362 79892
rect 155414 79840 155420 79892
rect 155218 79472 155224 79484
rect 154316 79444 155224 79472
rect 155218 79432 155224 79444
rect 155276 79432 155282 79484
rect 155374 79472 155402 79840
rect 155696 79540 155724 79920
rect 155926 79920 156190 79948
rect 155816 79840 155822 79892
rect 155874 79840 155880 79892
rect 155834 79756 155862 79840
rect 155770 79704 155776 79756
rect 155828 79716 155862 79756
rect 155828 79704 155834 79716
rect 155926 79676 155954 79920
rect 156184 79908 156190 79920
rect 156242 79908 156248 79960
rect 156368 79908 156374 79960
rect 156426 79908 156432 79960
rect 156460 79908 156466 79960
rect 156518 79908 156524 79960
rect 156828 79908 156834 79960
rect 156886 79908 156892 79960
rect 156000 79840 156006 79892
rect 156058 79880 156064 79892
rect 156058 79852 156138 79880
rect 156058 79840 156064 79852
rect 156110 79812 156138 79852
rect 156276 79840 156282 79892
rect 156334 79840 156340 79892
rect 156110 79784 156184 79812
rect 156156 79688 156184 79784
rect 156294 79688 156322 79840
rect 156386 79824 156414 79908
rect 156368 79772 156374 79824
rect 156426 79772 156432 79824
rect 156478 79744 156506 79908
rect 156736 79840 156742 79892
rect 156794 79840 156800 79892
rect 156846 79880 156874 79908
rect 156846 79852 157196 79880
rect 156644 79772 156650 79824
rect 156702 79772 156708 79824
rect 156046 79676 156052 79688
rect 155926 79648 156052 79676
rect 156046 79636 156052 79648
rect 156104 79636 156110 79688
rect 156138 79636 156144 79688
rect 156196 79636 156202 79688
rect 156230 79636 156236 79688
rect 156288 79648 156322 79688
rect 156386 79716 156506 79744
rect 156288 79636 156294 79648
rect 156386 79608 156414 79716
rect 156662 79688 156690 79772
rect 156598 79636 156604 79688
rect 156656 79648 156690 79688
rect 156656 79636 156662 79648
rect 156386 79580 156460 79608
rect 156322 79540 156328 79552
rect 155696 79512 156328 79540
rect 156322 79500 156328 79512
rect 156380 79500 156386 79552
rect 156432 79540 156460 79580
rect 156506 79568 156512 79620
rect 156564 79608 156570 79620
rect 156754 79608 156782 79840
rect 156920 79772 156926 79824
rect 156978 79812 156984 79824
rect 156978 79784 157104 79812
rect 156978 79772 156984 79784
rect 156564 79580 156782 79608
rect 156564 79568 156570 79580
rect 156966 79540 156972 79552
rect 156432 79512 156972 79540
rect 156966 79500 156972 79512
rect 157024 79500 157030 79552
rect 155862 79472 155868 79484
rect 155374 79444 155868 79472
rect 155862 79432 155868 79444
rect 155920 79432 155926 79484
rect 157076 79472 157104 79784
rect 157168 79688 157196 79852
rect 157380 79840 157386 79892
rect 157438 79840 157444 79892
rect 157840 79840 157846 79892
rect 157898 79840 157904 79892
rect 157288 79812 157294 79824
rect 157260 79772 157294 79812
rect 157346 79772 157352 79824
rect 157260 79688 157288 79772
rect 157398 79688 157426 79840
rect 157472 79772 157478 79824
rect 157530 79772 157536 79824
rect 157150 79636 157156 79688
rect 157208 79636 157214 79688
rect 157242 79636 157248 79688
rect 157300 79636 157306 79688
rect 157334 79636 157340 79688
rect 157392 79648 157426 79688
rect 157392 79636 157398 79648
rect 157490 79620 157518 79772
rect 157426 79568 157432 79620
rect 157484 79580 157518 79620
rect 157484 79568 157490 79580
rect 157610 79500 157616 79552
rect 157668 79540 157674 79552
rect 157858 79540 157886 79840
rect 157996 79620 158024 80736
rect 158456 80736 172514 80764
rect 158116 79840 158122 79892
rect 158174 79840 158180 79892
rect 157978 79568 157984 79620
rect 158036 79568 158042 79620
rect 158134 79608 158162 79840
rect 158346 79608 158352 79620
rect 158134 79580 158352 79608
rect 158346 79568 158352 79580
rect 158404 79568 158410 79620
rect 157668 79512 157886 79540
rect 157668 79500 157674 79512
rect 157886 79472 157892 79484
rect 157076 79444 157892 79472
rect 157886 79432 157892 79444
rect 157944 79432 157950 79484
rect 146266 79376 155264 79404
rect 143902 79336 143908 79348
rect 143736 79308 143908 79336
rect 143902 79296 143908 79308
rect 143960 79296 143966 79348
rect 144362 79296 144368 79348
rect 144420 79336 144426 79348
rect 146266 79336 146294 79376
rect 144420 79308 146294 79336
rect 144420 79296 144426 79308
rect 148410 79296 148416 79348
rect 148468 79336 148474 79348
rect 155034 79336 155040 79348
rect 148468 79308 155040 79336
rect 148468 79296 148474 79308
rect 155034 79296 155040 79308
rect 155092 79296 155098 79348
rect 131224 79240 139394 79268
rect 120442 79160 120448 79212
rect 120500 79200 120506 79212
rect 139026 79200 139032 79212
rect 120500 79172 139032 79200
rect 120500 79160 120506 79172
rect 139026 79160 139032 79172
rect 139084 79160 139090 79212
rect 139366 79200 139394 79240
rect 141970 79228 141976 79280
rect 142028 79268 142034 79280
rect 145466 79268 145472 79280
rect 142028 79240 145472 79268
rect 142028 79228 142034 79240
rect 145466 79228 145472 79240
rect 145524 79228 145530 79280
rect 155236 79268 155264 79376
rect 156690 79364 156696 79416
rect 156748 79404 156754 79416
rect 158456 79404 158484 80736
rect 172486 80696 172514 80736
rect 174924 80736 396816 80764
rect 174924 80708 174952 80736
rect 396810 80724 396816 80736
rect 396868 80724 396874 80776
rect 174814 80696 174820 80708
rect 159100 80668 164234 80696
rect 172486 80668 174820 80696
rect 158668 79908 158674 79960
rect 158726 79908 158732 79960
rect 158760 79908 158766 79960
rect 158818 79908 158824 79960
rect 158686 79620 158714 79908
rect 158622 79568 158628 79620
rect 158680 79580 158714 79620
rect 158680 79568 158686 79580
rect 156748 79376 158484 79404
rect 156748 79364 156754 79376
rect 158778 79336 158806 79908
rect 158898 79568 158904 79620
rect 158956 79608 158962 79620
rect 159100 79608 159128 80668
rect 164206 80628 164234 80668
rect 174814 80656 174820 80668
rect 174872 80656 174878 80708
rect 174906 80656 174912 80708
rect 174964 80656 174970 80708
rect 580350 80696 580356 80708
rect 182146 80668 580356 80696
rect 175918 80628 175924 80640
rect 164206 80600 169754 80628
rect 169726 80560 169754 80600
rect 172486 80600 175924 80628
rect 162826 80532 164234 80560
rect 169726 80532 171134 80560
rect 162826 80220 162854 80532
rect 164206 80356 164234 80532
rect 171106 80492 171134 80532
rect 172486 80492 172514 80600
rect 175918 80588 175924 80600
rect 175976 80588 175982 80640
rect 182146 80560 182174 80668
rect 580350 80656 580356 80668
rect 580408 80656 580414 80708
rect 393958 80628 393964 80640
rect 171106 80464 172514 80492
rect 173866 80532 182174 80560
rect 186286 80600 393964 80628
rect 173866 80356 173894 80532
rect 174722 80452 174728 80504
rect 174780 80492 174786 80504
rect 186286 80492 186314 80600
rect 393958 80588 393964 80600
rect 394016 80588 394022 80640
rect 174780 80464 186314 80492
rect 174780 80452 174786 80464
rect 175090 80384 175096 80436
rect 175148 80424 175154 80436
rect 180242 80424 180248 80436
rect 175148 80396 180248 80424
rect 175148 80384 175154 80396
rect 180242 80384 180248 80396
rect 180300 80384 180306 80436
rect 164206 80328 169754 80356
rect 169726 80288 169754 80328
rect 172026 80328 173894 80356
rect 169726 80260 171134 80288
rect 159928 80192 162854 80220
rect 159588 79948 159594 79960
rect 159330 79920 159594 79948
rect 159220 79840 159226 79892
rect 159278 79840 159284 79892
rect 159238 79744 159266 79840
rect 159192 79716 159266 79744
rect 159192 79688 159220 79716
rect 159174 79636 159180 79688
rect 159232 79636 159238 79688
rect 158956 79580 159128 79608
rect 158956 79568 158962 79580
rect 159330 79404 159358 79920
rect 159588 79908 159594 79920
rect 159646 79908 159652 79960
rect 159772 79908 159778 79960
rect 159830 79908 159836 79960
rect 159404 79840 159410 79892
rect 159462 79840 159468 79892
rect 159790 79880 159818 79908
rect 159744 79852 159818 79880
rect 159422 79472 159450 79840
rect 159744 79620 159772 79852
rect 159928 79620 159956 80192
rect 161446 80124 169708 80152
rect 161446 80016 161474 80124
rect 160250 79988 161474 80016
rect 162136 80056 169064 80084
rect 159726 79568 159732 79620
rect 159784 79568 159790 79620
rect 159910 79568 159916 79620
rect 159968 79568 159974 79620
rect 160002 79568 160008 79620
rect 160060 79608 160066 79620
rect 160250 79608 160278 79988
rect 160600 79908 160606 79960
rect 160658 79908 160664 79960
rect 161336 79908 161342 79960
rect 161394 79948 161400 79960
rect 161394 79908 161428 79948
rect 161888 79908 161894 79960
rect 161946 79908 161952 79960
rect 161980 79908 161986 79960
rect 162038 79908 162044 79960
rect 160324 79840 160330 79892
rect 160382 79840 160388 79892
rect 160618 79880 160646 79908
rect 160618 79852 161336 79880
rect 160342 79812 160370 79840
rect 160646 79812 160652 79824
rect 160342 79784 160652 79812
rect 160646 79772 160652 79784
rect 160704 79772 160710 79824
rect 160784 79772 160790 79824
rect 160842 79772 160848 79824
rect 161060 79772 161066 79824
rect 161118 79772 161124 79824
rect 160802 79688 160830 79772
rect 161078 79744 161106 79772
rect 160940 79716 161106 79744
rect 160802 79648 160836 79688
rect 160830 79636 160836 79648
rect 160888 79636 160894 79688
rect 160370 79608 160376 79620
rect 160060 79568 160094 79608
rect 160250 79580 160376 79608
rect 160370 79568 160376 79580
rect 160428 79568 160434 79620
rect 159910 79472 159916 79484
rect 159422 79444 159916 79472
rect 159910 79432 159916 79444
rect 159968 79432 159974 79484
rect 160066 79416 160094 79568
rect 160278 79500 160284 79552
rect 160336 79540 160342 79552
rect 160940 79540 160968 79716
rect 161308 79688 161336 79852
rect 161290 79636 161296 79688
rect 161348 79636 161354 79688
rect 161106 79568 161112 79620
rect 161164 79608 161170 79620
rect 161400 79608 161428 79908
rect 161906 79880 161934 79908
rect 161492 79852 161934 79880
rect 161998 79880 162026 79908
rect 161998 79852 162072 79880
rect 161492 79620 161520 79852
rect 161164 79580 161428 79608
rect 161164 79568 161170 79580
rect 161474 79568 161480 79620
rect 161532 79568 161538 79620
rect 161842 79568 161848 79620
rect 161900 79608 161906 79620
rect 162044 79608 162072 79852
rect 161900 79580 162072 79608
rect 161900 79568 161906 79580
rect 160336 79512 160968 79540
rect 160336 79500 160342 79512
rect 161014 79500 161020 79552
rect 161072 79540 161078 79552
rect 162136 79540 162164 80056
rect 169036 80016 169064 80056
rect 163010 79988 163544 80016
rect 163010 79960 163038 79988
rect 162716 79948 162722 79960
rect 162458 79920 162722 79948
rect 162256 79840 162262 79892
rect 162314 79840 162320 79892
rect 162274 79744 162302 79840
rect 162458 79812 162486 79920
rect 162716 79908 162722 79920
rect 162774 79908 162780 79960
rect 162992 79908 162998 79960
rect 163050 79908 163056 79960
rect 162532 79840 162538 79892
rect 162590 79880 162596 79892
rect 162590 79852 162900 79880
rect 162590 79840 162596 79852
rect 162458 79784 162716 79812
rect 162486 79744 162492 79756
rect 162274 79716 162492 79744
rect 162486 79704 162492 79716
rect 162544 79704 162550 79756
rect 162688 79688 162716 79784
rect 162670 79636 162676 79688
rect 162728 79636 162734 79688
rect 162872 79620 162900 79852
rect 163360 79840 163366 79892
rect 163418 79840 163424 79892
rect 162854 79568 162860 79620
rect 162912 79568 162918 79620
rect 163130 79568 163136 79620
rect 163188 79608 163194 79620
rect 163378 79608 163406 79840
rect 163516 79620 163544 79988
rect 163654 79988 166626 80016
rect 163654 79960 163682 79988
rect 163636 79908 163642 79960
rect 163694 79908 163700 79960
rect 164740 79948 164746 79960
rect 164252 79920 164746 79948
rect 163820 79840 163826 79892
rect 163878 79840 163884 79892
rect 163188 79580 163406 79608
rect 163188 79568 163194 79580
rect 163498 79568 163504 79620
rect 163556 79568 163562 79620
rect 163682 79568 163688 79620
rect 163740 79608 163746 79620
rect 163838 79608 163866 79840
rect 164252 79620 164280 79920
rect 164740 79908 164746 79920
rect 164798 79908 164804 79960
rect 166028 79948 166034 79960
rect 166000 79908 166034 79948
rect 166086 79908 166092 79960
rect 166120 79908 166126 79960
rect 166178 79908 166184 79960
rect 166212 79908 166218 79960
rect 166270 79908 166276 79960
rect 164372 79840 164378 79892
rect 164430 79840 164436 79892
rect 165752 79840 165758 79892
rect 165810 79840 165816 79892
rect 164390 79676 164418 79840
rect 165200 79772 165206 79824
rect 165258 79772 165264 79824
rect 164602 79676 164608 79688
rect 164390 79648 164608 79676
rect 164602 79636 164608 79648
rect 164660 79636 164666 79688
rect 163740 79580 163866 79608
rect 163740 79568 163746 79580
rect 164234 79568 164240 79620
rect 164292 79568 164298 79620
rect 165218 79608 165246 79772
rect 165770 79676 165798 79840
rect 166000 79824 166028 79908
rect 165982 79772 165988 79824
rect 166040 79772 166046 79824
rect 166138 79756 166166 79908
rect 166074 79704 166080 79756
rect 166132 79716 166166 79756
rect 166132 79704 166138 79716
rect 165890 79676 165896 79688
rect 165770 79648 165896 79676
rect 165890 79636 165896 79648
rect 165948 79636 165954 79688
rect 165338 79608 165344 79620
rect 165218 79580 165344 79608
rect 165338 79568 165344 79580
rect 165396 79568 165402 79620
rect 165614 79568 165620 79620
rect 165672 79608 165678 79620
rect 166230 79608 166258 79908
rect 166304 79840 166310 79892
rect 166362 79840 166368 79892
rect 165672 79580 166258 79608
rect 165672 79568 165678 79580
rect 161072 79512 162164 79540
rect 161072 79500 161078 79512
rect 162946 79500 162952 79552
rect 163004 79540 163010 79552
rect 163406 79540 163412 79552
rect 163004 79512 163412 79540
rect 163004 79500 163010 79512
rect 163406 79500 163412 79512
rect 163464 79500 163470 79552
rect 165798 79500 165804 79552
rect 165856 79540 165862 79552
rect 166322 79540 166350 79840
rect 165856 79512 166350 79540
rect 166598 79540 166626 79988
rect 167012 79988 167730 80016
rect 169036 79988 169110 80016
rect 166672 79908 166678 79960
rect 166730 79908 166736 79960
rect 166690 79608 166718 79908
rect 167012 79620 167040 79988
rect 167702 79960 167730 79988
rect 167592 79948 167598 79960
rect 167426 79920 167598 79948
rect 167426 79676 167454 79920
rect 167592 79908 167598 79920
rect 167650 79908 167656 79960
rect 167684 79908 167690 79960
rect 167742 79908 167748 79960
rect 167776 79908 167782 79960
rect 167834 79908 167840 79960
rect 167868 79908 167874 79960
rect 167926 79908 167932 79960
rect 168144 79908 168150 79960
rect 168202 79908 168208 79960
rect 168328 79948 168334 79960
rect 168300 79908 168334 79948
rect 168386 79908 168392 79960
rect 168788 79948 168794 79960
rect 168760 79908 168794 79948
rect 168846 79908 168852 79960
rect 168972 79908 168978 79960
rect 169030 79908 169036 79960
rect 169082 79948 169110 79988
rect 169082 79920 169432 79948
rect 167794 79880 167822 79908
rect 167656 79852 167822 79880
rect 167886 79880 167914 79908
rect 167886 79852 168098 79880
rect 167546 79676 167552 79688
rect 167426 79648 167552 79676
rect 167546 79636 167552 79648
rect 167604 79636 167610 79688
rect 166902 79608 166908 79620
rect 166690 79580 166908 79608
rect 166902 79568 166908 79580
rect 166960 79568 166966 79620
rect 166994 79568 167000 79620
rect 167052 79568 167058 79620
rect 167454 79568 167460 79620
rect 167512 79608 167518 79620
rect 167656 79608 167684 79852
rect 167730 79636 167736 79688
rect 167788 79676 167794 79688
rect 168070 79676 168098 79852
rect 167788 79648 168098 79676
rect 168162 79688 168190 79908
rect 168162 79648 168196 79688
rect 167788 79636 167794 79648
rect 168190 79636 168196 79648
rect 168248 79636 168254 79688
rect 167512 79580 167684 79608
rect 167512 79568 167518 79580
rect 168300 79552 168328 79908
rect 168512 79840 168518 79892
rect 168570 79840 168576 79892
rect 168604 79840 168610 79892
rect 168662 79840 168668 79892
rect 168374 79704 168380 79756
rect 168432 79744 168438 79756
rect 168530 79744 168558 79840
rect 168432 79716 168558 79744
rect 168432 79704 168438 79716
rect 168466 79636 168472 79688
rect 168524 79676 168530 79688
rect 168622 79676 168650 79840
rect 168760 79688 168788 79908
rect 168880 79880 168886 79892
rect 168852 79840 168886 79880
rect 168938 79840 168944 79892
rect 168524 79648 168650 79676
rect 168524 79636 168530 79648
rect 168742 79636 168748 79688
rect 168800 79636 168806 79688
rect 168852 79620 168880 79840
rect 168990 79812 169018 79908
rect 169064 79840 169070 79892
rect 169122 79840 169128 79892
rect 169156 79840 169162 79892
rect 169214 79840 169220 79892
rect 168944 79784 169018 79812
rect 168944 79756 168972 79784
rect 169082 79756 169110 79840
rect 168926 79704 168932 79756
rect 168984 79704 168990 79756
rect 169018 79704 169024 79756
rect 169076 79716 169110 79756
rect 169076 79704 169082 79716
rect 169174 79688 169202 79840
rect 169110 79636 169116 79688
rect 169168 79648 169202 79688
rect 169168 79636 169174 79648
rect 168834 79568 168840 79620
rect 168892 79568 168898 79620
rect 167822 79540 167828 79552
rect 166598 79512 167828 79540
rect 165856 79500 165862 79512
rect 167822 79500 167828 79512
rect 167880 79500 167886 79552
rect 168282 79500 168288 79552
rect 168340 79500 168346 79552
rect 169404 79484 169432 79920
rect 169524 79840 169530 79892
rect 169582 79840 169588 79892
rect 169542 79688 169570 79840
rect 169478 79636 169484 79688
rect 169536 79648 169570 79688
rect 169536 79636 169542 79648
rect 169680 79620 169708 80124
rect 171106 80016 171134 80260
rect 171106 79988 171962 80016
rect 169800 79908 169806 79960
rect 169858 79908 169864 79960
rect 170168 79948 170174 79960
rect 170048 79920 170174 79948
rect 169662 79568 169668 79620
rect 169720 79568 169726 79620
rect 169818 79540 169846 79908
rect 170048 79688 170076 79920
rect 170168 79908 170174 79920
rect 170226 79908 170232 79960
rect 170352 79908 170358 79960
rect 170410 79908 170416 79960
rect 170444 79908 170450 79960
rect 170502 79908 170508 79960
rect 170628 79908 170634 79960
rect 170686 79908 170692 79960
rect 170720 79908 170726 79960
rect 170778 79948 170784 79960
rect 170778 79920 171548 79948
rect 170778 79908 170784 79920
rect 170370 79880 170398 79908
rect 170232 79852 170398 79880
rect 170030 79636 170036 79688
rect 170088 79636 170094 79688
rect 170232 79608 170260 79852
rect 170462 79812 170490 79908
rect 170536 79840 170542 79892
rect 170594 79840 170600 79892
rect 170324 79784 170490 79812
rect 170324 79688 170352 79784
rect 170398 79704 170404 79756
rect 170456 79744 170462 79756
rect 170554 79744 170582 79840
rect 170456 79716 170582 79744
rect 170646 79744 170674 79908
rect 170904 79840 170910 79892
rect 170962 79840 170968 79892
rect 170996 79840 171002 79892
rect 171054 79840 171060 79892
rect 171180 79880 171186 79892
rect 171152 79840 171186 79880
rect 171238 79840 171244 79892
rect 170766 79772 170772 79824
rect 170824 79812 170830 79824
rect 170922 79812 170950 79840
rect 170824 79784 170950 79812
rect 170824 79772 170830 79784
rect 170858 79744 170864 79756
rect 170646 79716 170864 79744
rect 170456 79704 170462 79716
rect 170858 79704 170864 79716
rect 170916 79704 170922 79756
rect 170306 79636 170312 79688
rect 170364 79636 170370 79688
rect 171014 79620 171042 79840
rect 171152 79688 171180 79840
rect 171520 79744 171548 79920
rect 171824 79840 171830 79892
rect 171882 79840 171888 79892
rect 171934 79880 171962 79988
rect 172026 79960 172054 80328
rect 174446 80248 174452 80300
rect 174504 80288 174510 80300
rect 182174 80288 182180 80300
rect 174504 80260 182180 80288
rect 174504 80248 174510 80260
rect 182174 80248 182180 80260
rect 182232 80248 182238 80300
rect 200114 80220 200120 80232
rect 175844 80192 200120 80220
rect 175734 80152 175740 80164
rect 172578 80124 175740 80152
rect 172008 79908 172014 79960
rect 172066 79908 172072 79960
rect 172284 79908 172290 79960
rect 172342 79948 172348 79960
rect 172578 79948 172606 80124
rect 175734 80112 175740 80124
rect 175792 80112 175798 80164
rect 175844 80084 175872 80192
rect 200114 80180 200120 80192
rect 200172 80180 200178 80232
rect 177022 80112 177028 80164
rect 177080 80152 177086 80164
rect 231854 80152 231860 80164
rect 177080 80124 231860 80152
rect 177080 80112 177086 80124
rect 231854 80112 231860 80124
rect 231912 80112 231918 80164
rect 173268 80056 175872 80084
rect 172928 79948 172934 79960
rect 172342 79920 172606 79948
rect 172854 79920 172934 79948
rect 172342 79908 172348 79920
rect 172854 79880 172882 79920
rect 172928 79908 172934 79920
rect 172986 79908 172992 79960
rect 171934 79852 172882 79880
rect 171842 79812 171870 79840
rect 171962 79812 171968 79824
rect 171842 79784 171968 79812
rect 171962 79772 171968 79784
rect 172020 79772 172026 79824
rect 171520 79716 171640 79744
rect 171612 79688 171640 79716
rect 171870 79704 171876 79756
rect 171928 79744 171934 79756
rect 173268 79744 173296 80056
rect 175918 80044 175924 80096
rect 175976 80084 175982 80096
rect 252554 80084 252560 80096
rect 175976 80056 252560 80084
rect 175976 80044 175982 80056
rect 252554 80044 252560 80056
rect 252612 80044 252618 80096
rect 174814 80016 174820 80028
rect 173958 79988 174820 80016
rect 173958 79960 173986 79988
rect 174814 79976 174820 79988
rect 174872 79976 174878 80028
rect 173480 79908 173486 79960
rect 173538 79908 173544 79960
rect 173848 79908 173854 79960
rect 173906 79908 173912 79960
rect 173940 79908 173946 79960
rect 173998 79908 174004 79960
rect 174032 79908 174038 79960
rect 174090 79908 174096 79960
rect 174124 79908 174130 79960
rect 174182 79908 174188 79960
rect 173388 79840 173394 79892
rect 173446 79840 173452 79892
rect 171928 79716 173296 79744
rect 171928 79704 171934 79716
rect 171134 79636 171140 79688
rect 171192 79636 171198 79688
rect 171364 79636 171370 79688
rect 171422 79636 171428 79688
rect 171594 79636 171600 79688
rect 171652 79636 171658 79688
rect 173250 79636 173256 79688
rect 173308 79676 173314 79688
rect 173406 79676 173434 79840
rect 173308 79648 173434 79676
rect 173498 79676 173526 79908
rect 173756 79840 173762 79892
rect 173814 79840 173820 79892
rect 173774 79756 173802 79840
rect 173866 79824 173894 79908
rect 174050 79824 174078 79908
rect 174142 79880 174170 79908
rect 174142 79852 174216 79880
rect 174188 79824 174216 79852
rect 173866 79784 173900 79824
rect 173894 79772 173900 79784
rect 173952 79772 173958 79824
rect 173986 79772 173992 79824
rect 174044 79784 174078 79824
rect 174044 79772 174050 79784
rect 174170 79772 174176 79824
rect 174228 79772 174234 79824
rect 173774 79716 173808 79756
rect 173802 79704 173808 79716
rect 173860 79704 173866 79756
rect 173618 79676 173624 79688
rect 173498 79648 173624 79676
rect 173308 79636 173314 79648
rect 173618 79636 173624 79648
rect 173676 79636 173682 79688
rect 170490 79608 170496 79620
rect 170232 79580 170496 79608
rect 170490 79568 170496 79580
rect 170548 79568 170554 79620
rect 170950 79568 170956 79620
rect 171008 79580 171042 79620
rect 171382 79608 171410 79636
rect 174722 79608 174728 79620
rect 171382 79580 174728 79608
rect 171008 79568 171014 79580
rect 174722 79568 174728 79580
rect 174780 79568 174786 79620
rect 170398 79540 170404 79552
rect 169818 79512 170404 79540
rect 170398 79500 170404 79512
rect 170456 79500 170462 79552
rect 174170 79540 174176 79552
rect 170508 79512 174176 79540
rect 163222 79432 163228 79484
rect 163280 79472 163286 79484
rect 166442 79472 166448 79484
rect 163280 79444 166448 79472
rect 163280 79432 163286 79444
rect 166442 79432 166448 79444
rect 166500 79432 166506 79484
rect 169386 79432 169392 79484
rect 169444 79432 169450 79484
rect 159450 79404 159456 79416
rect 159330 79376 159456 79404
rect 159450 79364 159456 79376
rect 159508 79364 159514 79416
rect 160002 79364 160008 79416
rect 160060 79376 160094 79416
rect 160060 79364 160066 79376
rect 164326 79364 164332 79416
rect 164384 79404 164390 79416
rect 167638 79404 167644 79416
rect 164384 79376 167644 79404
rect 164384 79364 164390 79376
rect 167638 79364 167644 79376
rect 167696 79364 167702 79416
rect 163222 79336 163228 79348
rect 158778 79308 163228 79336
rect 163222 79296 163228 79308
rect 163280 79296 163286 79348
rect 163406 79296 163412 79348
rect 163464 79336 163470 79348
rect 170508 79336 170536 79512
rect 174170 79500 174176 79512
rect 174228 79500 174234 79552
rect 170674 79432 170680 79484
rect 170732 79472 170738 79484
rect 171870 79472 171876 79484
rect 170732 79444 171876 79472
rect 170732 79432 170738 79444
rect 171870 79432 171876 79444
rect 171928 79432 171934 79484
rect 173066 79432 173072 79484
rect 173124 79472 173130 79484
rect 173124 79444 180794 79472
rect 173124 79432 173130 79444
rect 171226 79364 171232 79416
rect 171284 79404 171290 79416
rect 171284 79376 178034 79404
rect 171284 79364 171290 79376
rect 163464 79308 170536 79336
rect 163464 79296 163470 79308
rect 171502 79296 171508 79348
rect 171560 79336 171566 79348
rect 174906 79336 174912 79348
rect 171560 79308 174912 79336
rect 171560 79296 171566 79308
rect 174906 79296 174912 79308
rect 174964 79296 174970 79348
rect 178006 79336 178034 79376
rect 180058 79336 180064 79348
rect 178006 79308 180064 79336
rect 180058 79296 180064 79308
rect 180116 79296 180122 79348
rect 180766 79336 180794 79444
rect 580534 79336 580540 79348
rect 180766 79308 580540 79336
rect 580534 79296 580540 79308
rect 580592 79296 580598 79348
rect 149026 79240 150434 79268
rect 155236 79240 160094 79268
rect 149026 79200 149054 79240
rect 139366 79172 149054 79200
rect 148410 79132 148416 79144
rect 118666 79104 148416 79132
rect 148410 79092 148416 79104
rect 148468 79092 148474 79144
rect 127526 79024 127532 79076
rect 127584 79064 127590 79076
rect 127710 79064 127716 79076
rect 127584 79036 127716 79064
rect 127584 79024 127590 79036
rect 127710 79024 127716 79036
rect 127768 79024 127774 79076
rect 141142 79024 141148 79076
rect 141200 79064 141206 79076
rect 141694 79064 141700 79076
rect 141200 79036 141700 79064
rect 141200 79024 141206 79036
rect 141694 79024 141700 79036
rect 141752 79024 141758 79076
rect 150406 79064 150434 79240
rect 155218 79160 155224 79212
rect 155276 79200 155282 79212
rect 156690 79200 156696 79212
rect 155276 79172 156696 79200
rect 155276 79160 155282 79172
rect 156690 79160 156696 79172
rect 156748 79160 156754 79212
rect 157978 79160 157984 79212
rect 158036 79200 158042 79212
rect 158990 79200 158996 79212
rect 158036 79172 158996 79200
rect 158036 79160 158042 79172
rect 158990 79160 158996 79172
rect 159048 79160 159054 79212
rect 160066 79200 160094 79240
rect 164142 79228 164148 79280
rect 164200 79268 164206 79280
rect 178126 79268 178132 79280
rect 164200 79240 178132 79268
rect 164200 79228 164206 79240
rect 178126 79228 178132 79240
rect 178184 79228 178190 79280
rect 173894 79200 173900 79212
rect 160066 79172 173900 79200
rect 173894 79160 173900 79172
rect 173952 79160 173958 79212
rect 164326 79092 164332 79144
rect 164384 79132 164390 79144
rect 195974 79132 195980 79144
rect 164384 79104 195980 79132
rect 164384 79092 164390 79104
rect 195974 79092 195980 79104
rect 196032 79092 196038 79144
rect 164786 79064 164792 79076
rect 150406 79036 164792 79064
rect 164786 79024 164792 79036
rect 164844 79024 164850 79076
rect 165154 79024 165160 79076
rect 165212 79064 165218 79076
rect 249794 79064 249800 79076
rect 165212 79036 249800 79064
rect 165212 79024 165218 79036
rect 249794 79024 249800 79036
rect 249852 79024 249858 79076
rect 118666 78968 144914 78996
rect 5074 78820 5080 78872
rect 5132 78860 5138 78872
rect 118666 78860 118694 78968
rect 140498 78888 140504 78940
rect 140556 78928 140562 78940
rect 144362 78928 144368 78940
rect 140556 78900 144368 78928
rect 140556 78888 140562 78900
rect 144362 78888 144368 78900
rect 144420 78888 144426 78940
rect 5132 78832 118694 78860
rect 144886 78860 144914 78968
rect 164050 78956 164056 79008
rect 164108 78996 164114 79008
rect 213914 78996 213920 79008
rect 164108 78968 213920 78996
rect 164108 78956 164114 78968
rect 213914 78956 213920 78968
rect 213972 78956 213978 79008
rect 147766 78888 147772 78940
rect 147824 78928 147830 78940
rect 267734 78928 267740 78940
rect 147824 78900 267740 78928
rect 147824 78888 147830 78900
rect 267734 78888 267740 78900
rect 267792 78888 267798 78940
rect 144886 78832 150434 78860
rect 5132 78820 5138 78832
rect 127710 78684 127716 78736
rect 127768 78724 127774 78736
rect 128998 78724 129004 78736
rect 127768 78696 129004 78724
rect 127768 78684 127774 78696
rect 128998 78684 129004 78696
rect 129056 78684 129062 78736
rect 150406 78724 150434 78832
rect 155218 78820 155224 78872
rect 155276 78860 155282 78872
rect 161014 78860 161020 78872
rect 155276 78832 161020 78860
rect 155276 78820 155282 78832
rect 161014 78820 161020 78832
rect 161072 78820 161078 78872
rect 173710 78860 173716 78872
rect 164896 78832 173716 78860
rect 164896 78724 164924 78832
rect 173710 78820 173716 78832
rect 173768 78820 173774 78872
rect 176654 78820 176660 78872
rect 176712 78860 176718 78872
rect 329098 78860 329104 78872
rect 176712 78832 329104 78860
rect 176712 78820 176718 78832
rect 329098 78820 329104 78832
rect 329156 78820 329162 78872
rect 166350 78752 166356 78804
rect 166408 78792 166414 78804
rect 444374 78792 444380 78804
rect 166408 78764 444380 78792
rect 166408 78752 166414 78764
rect 444374 78752 444380 78764
rect 444432 78752 444438 78804
rect 150406 78696 164924 78724
rect 168650 78684 168656 78736
rect 168708 78724 168714 78736
rect 554774 78724 554780 78736
rect 168708 78696 554780 78724
rect 168708 78684 168714 78696
rect 554774 78684 554780 78696
rect 554832 78684 554838 78736
rect 126054 78616 126060 78668
rect 126112 78656 126118 78668
rect 126330 78656 126336 78668
rect 126112 78628 126336 78656
rect 126112 78616 126118 78628
rect 126330 78616 126336 78628
rect 126388 78616 126394 78668
rect 128722 78616 128728 78668
rect 128780 78656 128786 78668
rect 129366 78656 129372 78668
rect 128780 78628 129372 78656
rect 128780 78616 128786 78628
rect 129366 78616 129372 78628
rect 129424 78616 129430 78668
rect 137186 78616 137192 78668
rect 137244 78656 137250 78668
rect 137462 78656 137468 78668
rect 137244 78628 137468 78656
rect 137244 78616 137250 78628
rect 137462 78616 137468 78628
rect 137520 78616 137526 78668
rect 145190 78616 145196 78668
rect 145248 78656 145254 78668
rect 158898 78656 158904 78668
rect 145248 78628 158904 78656
rect 145248 78616 145254 78628
rect 158898 78616 158904 78628
rect 158956 78616 158962 78668
rect 163222 78616 163228 78668
rect 163280 78656 163286 78668
rect 171686 78656 171692 78668
rect 163280 78628 171692 78656
rect 163280 78616 163286 78628
rect 171686 78616 171692 78628
rect 171744 78616 171750 78668
rect 171778 78616 171784 78668
rect 171836 78656 171842 78668
rect 178586 78656 178592 78668
rect 171836 78628 178592 78656
rect 171836 78616 171842 78628
rect 178586 78616 178592 78628
rect 178644 78616 178650 78668
rect 139210 78548 139216 78600
rect 139268 78588 139274 78600
rect 140498 78588 140504 78600
rect 139268 78560 140504 78588
rect 139268 78548 139274 78560
rect 140498 78548 140504 78560
rect 140556 78548 140562 78600
rect 144914 78548 144920 78600
rect 144972 78588 144978 78600
rect 165154 78588 165160 78600
rect 144972 78560 165160 78588
rect 144972 78548 144978 78560
rect 165154 78548 165160 78560
rect 165212 78548 165218 78600
rect 166442 78548 166448 78600
rect 166500 78588 166506 78600
rect 171502 78588 171508 78600
rect 166500 78560 171508 78588
rect 166500 78548 166506 78560
rect 171502 78548 171508 78560
rect 171560 78548 171566 78600
rect 172330 78548 172336 78600
rect 172388 78588 172394 78600
rect 176562 78588 176568 78600
rect 172388 78560 176568 78588
rect 172388 78548 172394 78560
rect 176562 78548 176568 78560
rect 176620 78548 176626 78600
rect 126330 78480 126336 78532
rect 126388 78520 126394 78532
rect 130562 78520 130568 78532
rect 126388 78492 130568 78520
rect 126388 78480 126394 78492
rect 130562 78480 130568 78492
rect 130620 78480 130626 78532
rect 140682 78480 140688 78532
rect 140740 78520 140746 78532
rect 164326 78520 164332 78532
rect 140740 78492 164332 78520
rect 140740 78480 140746 78492
rect 164326 78480 164332 78492
rect 164384 78480 164390 78532
rect 170122 78480 170128 78532
rect 170180 78520 170186 78532
rect 170582 78520 170588 78532
rect 170180 78492 170588 78520
rect 170180 78480 170186 78492
rect 170582 78480 170588 78492
rect 170640 78480 170646 78532
rect 141050 78412 141056 78464
rect 141108 78452 141114 78464
rect 155218 78452 155224 78464
rect 141108 78424 155224 78452
rect 141108 78412 141114 78424
rect 155218 78412 155224 78424
rect 155276 78412 155282 78464
rect 161198 78412 161204 78464
rect 161256 78452 161262 78464
rect 161256 78424 164740 78452
rect 161256 78412 161262 78424
rect 146754 78344 146760 78396
rect 146812 78384 146818 78396
rect 164050 78384 164056 78396
rect 146812 78356 164056 78384
rect 146812 78344 146818 78356
rect 164050 78344 164056 78356
rect 164108 78344 164114 78396
rect 132402 78316 132408 78328
rect 125566 78288 132408 78316
rect 125042 78208 125048 78260
rect 125100 78248 125106 78260
rect 125566 78248 125594 78288
rect 132402 78276 132408 78288
rect 132460 78276 132466 78328
rect 154298 78276 154304 78328
rect 154356 78316 154362 78328
rect 162394 78316 162400 78328
rect 154356 78288 162400 78316
rect 154356 78276 154362 78288
rect 162394 78276 162400 78288
rect 162452 78276 162458 78328
rect 164712 78316 164740 78424
rect 164786 78412 164792 78464
rect 164844 78452 164850 78464
rect 173802 78452 173808 78464
rect 164844 78424 173808 78452
rect 164844 78412 164850 78424
rect 173802 78412 173808 78424
rect 173860 78412 173866 78464
rect 165706 78344 165712 78396
rect 165764 78384 165770 78396
rect 171870 78384 171876 78396
rect 165764 78356 171876 78384
rect 165764 78344 165770 78356
rect 171870 78344 171876 78356
rect 171928 78344 171934 78396
rect 173986 78344 173992 78396
rect 174044 78384 174050 78396
rect 174538 78384 174544 78396
rect 174044 78356 174544 78384
rect 174044 78344 174050 78356
rect 174538 78344 174544 78356
rect 174596 78344 174602 78396
rect 247678 78316 247684 78328
rect 164712 78288 247684 78316
rect 247678 78276 247684 78288
rect 247736 78276 247742 78328
rect 125100 78220 125594 78248
rect 125100 78208 125106 78220
rect 133506 78208 133512 78260
rect 133564 78248 133570 78260
rect 136910 78248 136916 78260
rect 133564 78220 136916 78248
rect 133564 78208 133570 78220
rect 136910 78208 136916 78220
rect 136968 78208 136974 78260
rect 146386 78208 146392 78260
rect 146444 78248 146450 78260
rect 147030 78248 147036 78260
rect 146444 78220 147036 78248
rect 146444 78208 146450 78220
rect 147030 78208 147036 78220
rect 147088 78208 147094 78260
rect 161658 78208 161664 78260
rect 161716 78248 161722 78260
rect 253198 78248 253204 78260
rect 161716 78220 253204 78248
rect 161716 78208 161722 78220
rect 253198 78208 253204 78220
rect 253256 78208 253262 78260
rect 89714 78140 89720 78192
rect 89772 78180 89778 78192
rect 132494 78180 132500 78192
rect 89772 78152 132500 78180
rect 89772 78140 89778 78152
rect 132494 78140 132500 78152
rect 132552 78140 132558 78192
rect 148134 78140 148140 78192
rect 148192 78180 148198 78192
rect 148318 78180 148324 78192
rect 148192 78152 148324 78180
rect 148192 78140 148198 78152
rect 148318 78140 148324 78152
rect 148376 78140 148382 78192
rect 153102 78140 153108 78192
rect 153160 78180 153166 78192
rect 161014 78180 161020 78192
rect 153160 78152 161020 78180
rect 153160 78140 153166 78152
rect 161014 78140 161020 78152
rect 161072 78140 161078 78192
rect 171594 78140 171600 78192
rect 171652 78180 171658 78192
rect 322198 78180 322204 78192
rect 171652 78152 322204 78180
rect 171652 78140 171658 78152
rect 322198 78140 322204 78152
rect 322256 78140 322262 78192
rect 46198 78072 46204 78124
rect 46256 78112 46262 78124
rect 126698 78112 126704 78124
rect 46256 78084 126704 78112
rect 46256 78072 46262 78084
rect 126698 78072 126704 78084
rect 126756 78072 126762 78124
rect 136818 78072 136824 78124
rect 136876 78112 136882 78124
rect 137462 78112 137468 78124
rect 136876 78084 137468 78112
rect 136876 78072 136882 78084
rect 137462 78072 137468 78084
rect 137520 78072 137526 78124
rect 140866 78072 140872 78124
rect 140924 78112 140930 78124
rect 150158 78112 150164 78124
rect 140924 78084 150164 78112
rect 140924 78072 140930 78084
rect 150158 78072 150164 78084
rect 150216 78072 150222 78124
rect 158898 78072 158904 78124
rect 158956 78112 158962 78124
rect 159542 78112 159548 78124
rect 158956 78084 159548 78112
rect 158956 78072 158962 78084
rect 159542 78072 159548 78084
rect 159600 78072 159606 78124
rect 162486 78072 162492 78124
rect 162544 78112 162550 78124
rect 471974 78112 471980 78124
rect 162544 78084 471980 78112
rect 162544 78072 162550 78084
rect 471974 78072 471980 78084
rect 472032 78072 472038 78124
rect 57238 78004 57244 78056
rect 57296 78044 57302 78056
rect 127618 78044 127624 78056
rect 57296 78016 127624 78044
rect 57296 78004 57302 78016
rect 127618 78004 127624 78016
rect 127676 78004 127682 78056
rect 149238 78004 149244 78056
rect 149296 78044 149302 78056
rect 149790 78044 149796 78056
rect 149296 78016 149796 78044
rect 149296 78004 149302 78016
rect 149790 78004 149796 78016
rect 149848 78004 149854 78056
rect 163958 78004 163964 78056
rect 164016 78044 164022 78056
rect 480254 78044 480260 78056
rect 164016 78016 480260 78044
rect 164016 78004 164022 78016
rect 480254 78004 480260 78016
rect 480312 78004 480318 78056
rect 22738 77936 22744 77988
rect 22796 77976 22802 77988
rect 125686 77976 125692 77988
rect 22796 77948 125692 77976
rect 22796 77936 22802 77948
rect 125686 77936 125692 77948
rect 125744 77936 125750 77988
rect 134518 77936 134524 77988
rect 134576 77976 134582 77988
rect 135254 77976 135260 77988
rect 134576 77948 135260 77976
rect 134576 77936 134582 77948
rect 135254 77936 135260 77948
rect 135312 77936 135318 77988
rect 147858 77936 147864 77988
rect 147916 77976 147922 77988
rect 148134 77976 148140 77988
rect 147916 77948 148140 77976
rect 147916 77936 147922 77948
rect 148134 77936 148140 77948
rect 148192 77936 148198 77988
rect 150066 77936 150072 77988
rect 150124 77976 150130 77988
rect 157058 77976 157064 77988
rect 150124 77948 157064 77976
rect 150124 77936 150130 77948
rect 157058 77936 157064 77948
rect 157116 77936 157122 77988
rect 167638 77936 167644 77988
rect 167696 77976 167702 77988
rect 498194 77976 498200 77988
rect 167696 77948 498200 77976
rect 167696 77936 167702 77948
rect 498194 77936 498200 77948
rect 498252 77936 498258 77988
rect 125318 77868 125324 77920
rect 125376 77908 125382 77920
rect 133414 77908 133420 77920
rect 125376 77880 133420 77908
rect 125376 77868 125382 77880
rect 133414 77868 133420 77880
rect 133472 77868 133478 77920
rect 152458 77868 152464 77920
rect 152516 77908 152522 77920
rect 159634 77908 159640 77920
rect 152516 77880 159640 77908
rect 152516 77868 152522 77880
rect 159634 77868 159640 77880
rect 159692 77868 159698 77920
rect 161290 77868 161296 77920
rect 161348 77908 161354 77920
rect 180058 77908 180064 77920
rect 161348 77880 180064 77908
rect 161348 77868 161354 77880
rect 180058 77868 180064 77880
rect 180116 77868 180122 77920
rect 125226 77800 125232 77852
rect 125284 77840 125290 77852
rect 129458 77840 129464 77852
rect 125284 77812 129464 77840
rect 125284 77800 125290 77812
rect 129458 77800 129464 77812
rect 129516 77800 129522 77852
rect 159174 77800 159180 77852
rect 159232 77840 159238 77852
rect 170214 77840 170220 77852
rect 159232 77812 170220 77840
rect 159232 77800 159238 77812
rect 170214 77800 170220 77812
rect 170272 77800 170278 77852
rect 123570 77732 123576 77784
rect 123628 77772 123634 77784
rect 132770 77772 132776 77784
rect 123628 77744 132776 77772
rect 123628 77732 123634 77744
rect 132770 77732 132776 77744
rect 132828 77732 132834 77784
rect 158622 77732 158628 77784
rect 158680 77772 158686 77784
rect 174538 77772 174544 77784
rect 158680 77744 174544 77772
rect 158680 77732 158686 77744
rect 174538 77732 174544 77744
rect 174596 77732 174602 77784
rect 120810 77664 120816 77716
rect 120868 77704 120874 77716
rect 128998 77704 129004 77716
rect 120868 77676 129004 77704
rect 120868 77664 120874 77676
rect 128998 77664 129004 77676
rect 129056 77664 129062 77716
rect 129090 77664 129096 77716
rect 129148 77704 129154 77716
rect 130286 77704 130292 77716
rect 129148 77676 130292 77704
rect 129148 77664 129154 77676
rect 130286 77664 130292 77676
rect 130344 77664 130350 77716
rect 141694 77664 141700 77716
rect 141752 77704 141758 77716
rect 141752 77676 150434 77704
rect 141752 77664 141758 77676
rect 120626 77596 120632 77648
rect 120684 77636 120690 77648
rect 128446 77636 128452 77648
rect 120684 77608 128452 77636
rect 120684 77596 120690 77608
rect 128446 77596 128452 77608
rect 128504 77596 128510 77648
rect 122282 77528 122288 77580
rect 122340 77568 122346 77580
rect 128078 77568 128084 77580
rect 122340 77540 128084 77568
rect 122340 77528 122346 77540
rect 128078 77528 128084 77540
rect 128136 77528 128142 77580
rect 128998 77528 129004 77580
rect 129056 77568 129062 77580
rect 131390 77568 131396 77580
rect 129056 77540 131396 77568
rect 129056 77528 129062 77540
rect 131390 77528 131396 77540
rect 131448 77528 131454 77580
rect 143442 77528 143448 77580
rect 143500 77568 143506 77580
rect 150406 77568 150434 77676
rect 158346 77664 158352 77716
rect 158404 77704 158410 77716
rect 172422 77704 172428 77716
rect 158404 77676 172428 77704
rect 158404 77664 158410 77676
rect 172422 77664 172428 77676
rect 172480 77664 172486 77716
rect 157518 77596 157524 77648
rect 157576 77636 157582 77648
rect 171410 77636 171416 77648
rect 157576 77608 171416 77636
rect 157576 77596 157582 77608
rect 171410 77596 171416 77608
rect 171468 77596 171474 77648
rect 174446 77636 174452 77648
rect 171612 77608 174452 77636
rect 171612 77568 171640 77608
rect 174446 77596 174452 77608
rect 174504 77596 174510 77648
rect 143500 77540 149054 77568
rect 150406 77540 171640 77568
rect 143500 77528 143506 77540
rect 122098 77460 122104 77512
rect 122156 77500 122162 77512
rect 125870 77500 125876 77512
rect 122156 77472 125876 77500
rect 122156 77460 122162 77472
rect 125870 77460 125876 77472
rect 125928 77460 125934 77512
rect 127618 77392 127624 77444
rect 127676 77432 127682 77444
rect 129182 77432 129188 77444
rect 127676 77404 129188 77432
rect 127676 77392 127682 77404
rect 129182 77392 129188 77404
rect 129240 77392 129246 77444
rect 149026 77432 149054 77540
rect 172054 77528 172060 77580
rect 172112 77568 172118 77580
rect 580718 77568 580724 77580
rect 172112 77540 580724 77568
rect 172112 77528 172118 77540
rect 580718 77528 580724 77540
rect 580776 77528 580782 77580
rect 155218 77460 155224 77512
rect 155276 77500 155282 77512
rect 164142 77500 164148 77512
rect 155276 77472 164148 77500
rect 155276 77460 155282 77472
rect 164142 77460 164148 77472
rect 164200 77460 164206 77512
rect 164510 77460 164516 77512
rect 164568 77500 164574 77512
rect 166442 77500 166448 77512
rect 164568 77472 166448 77500
rect 164568 77460 164574 77472
rect 166442 77460 166448 77472
rect 166500 77460 166506 77512
rect 170214 77460 170220 77512
rect 170272 77500 170278 77512
rect 175918 77500 175924 77512
rect 170272 77472 175924 77500
rect 170272 77460 170278 77472
rect 175918 77460 175924 77472
rect 175976 77460 175982 77512
rect 177022 77432 177028 77444
rect 149026 77404 177028 77432
rect 177022 77392 177028 77404
rect 177080 77392 177086 77444
rect 124950 77324 124956 77376
rect 125008 77364 125014 77376
rect 126514 77364 126520 77376
rect 125008 77336 126520 77364
rect 125008 77324 125014 77336
rect 126514 77324 126520 77336
rect 126572 77324 126578 77376
rect 129826 77324 129832 77376
rect 129884 77364 129890 77376
rect 134886 77364 134892 77376
rect 129884 77336 134892 77364
rect 129884 77324 129890 77336
rect 134886 77324 134892 77336
rect 134944 77324 134950 77376
rect 139394 77324 139400 77376
rect 139452 77364 139458 77376
rect 155218 77364 155224 77376
rect 139452 77336 155224 77364
rect 139452 77324 139458 77336
rect 155218 77324 155224 77336
rect 155276 77324 155282 77376
rect 164786 77364 164792 77376
rect 156248 77336 164792 77364
rect 120718 77256 120724 77308
rect 120776 77296 120782 77308
rect 120776 77268 124260 77296
rect 120776 77256 120782 77268
rect 124232 77228 124260 77268
rect 125134 77256 125140 77308
rect 125192 77296 125198 77308
rect 126974 77296 126980 77308
rect 125192 77268 126980 77296
rect 125192 77256 125198 77268
rect 126974 77256 126980 77268
rect 127032 77256 127038 77308
rect 132494 77256 132500 77308
rect 132552 77296 132558 77308
rect 133874 77296 133880 77308
rect 132552 77268 133880 77296
rect 132552 77256 132558 77268
rect 133874 77256 133880 77268
rect 133932 77256 133938 77308
rect 153562 77256 153568 77308
rect 153620 77296 153626 77308
rect 156248 77296 156276 77336
rect 164786 77324 164792 77336
rect 164844 77324 164850 77376
rect 168282 77324 168288 77376
rect 168340 77364 168346 77376
rect 169386 77364 169392 77376
rect 168340 77336 169392 77364
rect 168340 77324 168346 77336
rect 169386 77324 169392 77336
rect 169444 77324 169450 77376
rect 153620 77268 156276 77296
rect 153620 77256 153626 77268
rect 156322 77256 156328 77308
rect 156380 77296 156386 77308
rect 165154 77296 165160 77308
rect 156380 77268 165160 77296
rect 156380 77256 156386 77268
rect 165154 77256 165160 77268
rect 165212 77256 165218 77308
rect 167086 77256 167092 77308
rect 167144 77296 167150 77308
rect 173158 77296 173164 77308
rect 167144 77268 173164 77296
rect 167144 77256 167150 77268
rect 173158 77256 173164 77268
rect 173216 77256 173222 77308
rect 124232 77200 128354 77228
rect 128326 77160 128354 77200
rect 153194 77188 153200 77240
rect 153252 77228 153258 77240
rect 153470 77228 153476 77240
rect 153252 77200 153476 77228
rect 153252 77188 153258 77200
rect 153470 77188 153476 77200
rect 153528 77188 153534 77240
rect 156138 77188 156144 77240
rect 156196 77228 156202 77240
rect 156966 77228 156972 77240
rect 156196 77200 156972 77228
rect 156196 77188 156202 77200
rect 156966 77188 156972 77200
rect 157024 77188 157030 77240
rect 162210 77188 162216 77240
rect 162268 77228 162274 77240
rect 167914 77228 167920 77240
rect 162268 77200 167920 77228
rect 162268 77188 162274 77200
rect 167914 77188 167920 77200
rect 167972 77188 167978 77240
rect 168282 77188 168288 77240
rect 168340 77228 168346 77240
rect 168834 77228 168840 77240
rect 168340 77200 168840 77228
rect 168340 77188 168346 77200
rect 168834 77188 168840 77200
rect 168892 77188 168898 77240
rect 175734 77188 175740 77240
rect 175792 77228 175798 77240
rect 527174 77228 527180 77240
rect 175792 77200 527180 77228
rect 175792 77188 175798 77200
rect 527174 77188 527180 77200
rect 527232 77188 527238 77240
rect 172606 77160 172612 77172
rect 128326 77132 172612 77160
rect 172606 77120 172612 77132
rect 172664 77120 172670 77172
rect 145098 77052 145104 77104
rect 145156 77092 145162 77104
rect 147398 77092 147404 77104
rect 145156 77064 147404 77092
rect 145156 77052 145162 77064
rect 147398 77052 147404 77064
rect 147456 77052 147462 77104
rect 150158 77052 150164 77104
rect 150216 77092 150222 77104
rect 197354 77092 197360 77104
rect 150216 77064 197360 77092
rect 150216 77052 150222 77064
rect 197354 77052 197360 77064
rect 197412 77052 197418 77104
rect 124858 76984 124864 77036
rect 124916 77024 124922 77036
rect 134794 77024 134800 77036
rect 124916 76996 134800 77024
rect 124916 76984 124922 76996
rect 134794 76984 134800 76996
rect 134852 76984 134858 77036
rect 152182 76984 152188 77036
rect 152240 77024 152246 77036
rect 152458 77024 152464 77036
rect 152240 76996 152464 77024
rect 152240 76984 152246 76996
rect 152458 76984 152464 76996
rect 152516 76984 152522 77036
rect 153470 76984 153476 77036
rect 153528 77024 153534 77036
rect 154114 77024 154120 77036
rect 153528 76996 154120 77024
rect 153528 76984 153534 76996
rect 154114 76984 154120 76996
rect 154172 76984 154178 77036
rect 157426 76984 157432 77036
rect 157484 77024 157490 77036
rect 158622 77024 158628 77036
rect 157484 76996 158628 77024
rect 157484 76984 157490 76996
rect 158622 76984 158628 76996
rect 158680 76984 158686 77036
rect 162762 76984 162768 77036
rect 162820 77024 162826 77036
rect 211798 77024 211804 77036
rect 162820 76996 211804 77024
rect 162820 76984 162826 76996
rect 211798 76984 211804 76996
rect 211856 76984 211862 77036
rect 133414 76916 133420 76968
rect 133472 76956 133478 76968
rect 135530 76956 135536 76968
rect 133472 76928 135536 76956
rect 133472 76916 133478 76928
rect 135530 76916 135536 76928
rect 135588 76916 135594 76968
rect 143166 76916 143172 76968
rect 143224 76956 143230 76968
rect 226334 76956 226340 76968
rect 143224 76928 226340 76956
rect 143224 76916 143230 76928
rect 226334 76916 226340 76928
rect 226392 76916 226398 76968
rect 122834 76848 122840 76900
rect 122892 76888 122898 76900
rect 135070 76888 135076 76900
rect 122892 76860 135076 76888
rect 122892 76848 122898 76860
rect 135070 76848 135076 76860
rect 135128 76848 135134 76900
rect 144270 76848 144276 76900
rect 144328 76888 144334 76900
rect 240134 76888 240140 76900
rect 144328 76860 240140 76888
rect 144328 76848 144334 76860
rect 240134 76848 240140 76860
rect 240192 76848 240198 76900
rect 102134 76780 102140 76832
rect 102192 76820 102198 76832
rect 102192 76792 128354 76820
rect 102192 76780 102198 76792
rect 86954 76712 86960 76764
rect 87012 76752 87018 76764
rect 123478 76752 123484 76764
rect 87012 76724 123484 76752
rect 87012 76712 87018 76724
rect 123478 76712 123484 76724
rect 123536 76712 123542 76764
rect 128326 76752 128354 76792
rect 131390 76780 131396 76832
rect 131448 76820 131454 76832
rect 131758 76820 131764 76832
rect 131448 76792 131764 76820
rect 131448 76780 131454 76792
rect 131758 76780 131764 76792
rect 131816 76780 131822 76832
rect 134242 76780 134248 76832
rect 134300 76820 134306 76832
rect 134610 76820 134616 76832
rect 134300 76792 134616 76820
rect 134300 76780 134306 76792
rect 134610 76780 134616 76792
rect 134668 76780 134674 76832
rect 145926 76780 145932 76832
rect 145984 76820 145990 76832
rect 260834 76820 260840 76832
rect 145984 76792 260840 76820
rect 145984 76780 145990 76792
rect 260834 76780 260840 76792
rect 260892 76780 260898 76832
rect 133230 76752 133236 76764
rect 128326 76724 133236 76752
rect 133230 76712 133236 76724
rect 133288 76712 133294 76764
rect 133874 76712 133880 76764
rect 133932 76752 133938 76764
rect 135898 76752 135904 76764
rect 133932 76724 135904 76752
rect 133932 76712 133938 76724
rect 135898 76712 135904 76724
rect 135956 76712 135962 76764
rect 140222 76712 140228 76764
rect 140280 76752 140286 76764
rect 140406 76752 140412 76764
rect 140280 76724 140412 76752
rect 140280 76712 140286 76724
rect 140406 76712 140412 76724
rect 140464 76712 140470 76764
rect 147950 76712 147956 76764
rect 148008 76752 148014 76764
rect 288434 76752 288440 76764
rect 148008 76724 288440 76752
rect 148008 76712 148014 76724
rect 288434 76712 288440 76724
rect 288492 76712 288498 76764
rect 69014 76644 69020 76696
rect 69072 76684 69078 76696
rect 130930 76684 130936 76696
rect 69072 76656 130936 76684
rect 69072 76644 69078 76656
rect 130930 76644 130936 76656
rect 130988 76644 130994 76696
rect 133046 76644 133052 76696
rect 133104 76684 133110 76696
rect 133782 76684 133788 76696
rect 133104 76656 133788 76684
rect 133104 76644 133110 76656
rect 133782 76644 133788 76656
rect 133840 76644 133846 76696
rect 148870 76644 148876 76696
rect 148928 76684 148934 76696
rect 296714 76684 296720 76696
rect 148928 76656 296720 76684
rect 148928 76644 148934 76656
rect 296714 76644 296720 76656
rect 296772 76644 296778 76696
rect 44174 76576 44180 76628
rect 44232 76616 44238 76628
rect 128814 76616 128820 76628
rect 44232 76588 128820 76616
rect 44232 76576 44238 76588
rect 128814 76576 128820 76588
rect 128872 76576 128878 76628
rect 134426 76576 134432 76628
rect 134484 76616 134490 76628
rect 135162 76616 135168 76628
rect 134484 76588 135168 76616
rect 134484 76576 134490 76588
rect 135162 76576 135168 76588
rect 135220 76576 135226 76628
rect 135898 76576 135904 76628
rect 135956 76616 135962 76628
rect 136450 76616 136456 76628
rect 135956 76588 136456 76616
rect 135956 76576 135962 76588
rect 136450 76576 136456 76588
rect 136508 76576 136514 76628
rect 136634 76576 136640 76628
rect 136692 76616 136698 76628
rect 136818 76616 136824 76628
rect 136692 76588 136824 76616
rect 136692 76576 136698 76588
rect 136818 76576 136824 76588
rect 136876 76576 136882 76628
rect 137094 76576 137100 76628
rect 137152 76616 137158 76628
rect 137738 76616 137744 76628
rect 137152 76588 137744 76616
rect 137152 76576 137158 76588
rect 137738 76576 137744 76588
rect 137796 76576 137802 76628
rect 150894 76576 150900 76628
rect 150952 76616 150958 76628
rect 151078 76616 151084 76628
rect 150952 76588 151084 76616
rect 150952 76576 150958 76588
rect 151078 76576 151084 76588
rect 151136 76576 151142 76628
rect 152182 76576 152188 76628
rect 152240 76616 152246 76628
rect 152550 76616 152556 76628
rect 152240 76588 152556 76616
rect 152240 76576 152246 76588
rect 152550 76576 152556 76588
rect 152608 76576 152614 76628
rect 153286 76576 153292 76628
rect 153344 76616 153350 76628
rect 153562 76616 153568 76628
rect 153344 76588 153568 76616
rect 153344 76576 153350 76588
rect 153562 76576 153568 76588
rect 153620 76576 153626 76628
rect 154758 76576 154764 76628
rect 154816 76616 154822 76628
rect 155218 76616 155224 76628
rect 154816 76588 155224 76616
rect 154816 76576 154822 76588
rect 155218 76576 155224 76588
rect 155276 76576 155282 76628
rect 156138 76576 156144 76628
rect 156196 76616 156202 76628
rect 156598 76616 156604 76628
rect 156196 76588 156604 76616
rect 156196 76576 156202 76588
rect 156598 76576 156604 76588
rect 156656 76576 156662 76628
rect 156690 76576 156696 76628
rect 156748 76616 156754 76628
rect 157150 76616 157156 76628
rect 156748 76588 157156 76616
rect 156748 76576 156754 76588
rect 157150 76576 157156 76588
rect 157208 76576 157214 76628
rect 157702 76576 157708 76628
rect 157760 76616 157766 76628
rect 157886 76616 157892 76628
rect 157760 76588 157892 76616
rect 157760 76576 157766 76588
rect 157886 76576 157892 76588
rect 157944 76576 157950 76628
rect 159634 76576 159640 76628
rect 159692 76616 159698 76628
rect 324406 76616 324412 76628
rect 159692 76588 324412 76616
rect 159692 76576 159698 76588
rect 324406 76576 324412 76588
rect 324464 76576 324470 76628
rect 30374 76508 30380 76560
rect 30432 76548 30438 76560
rect 127986 76548 127992 76560
rect 30432 76520 127992 76548
rect 30432 76508 30438 76520
rect 127986 76508 127992 76520
rect 128044 76508 128050 76560
rect 128096 76520 138014 76548
rect 124214 76440 124220 76492
rect 124272 76480 124278 76492
rect 128096 76480 128124 76520
rect 132218 76480 132224 76492
rect 124272 76452 128124 76480
rect 128188 76452 132224 76480
rect 124272 76440 124278 76452
rect 123478 76372 123484 76424
rect 123536 76412 123542 76424
rect 128188 76412 128216 76452
rect 132218 76440 132224 76452
rect 132276 76440 132282 76492
rect 137986 76480 138014 76520
rect 151906 76508 151912 76560
rect 151964 76548 151970 76560
rect 152366 76548 152372 76560
rect 151964 76520 152372 76548
rect 151964 76508 151970 76520
rect 152366 76508 152372 76520
rect 152424 76508 152430 76560
rect 158714 76508 158720 76560
rect 158772 76548 158778 76560
rect 159266 76548 159272 76560
rect 158772 76520 159272 76548
rect 158772 76508 158778 76520
rect 159266 76508 159272 76520
rect 159324 76508 159330 76560
rect 160278 76508 160284 76560
rect 160336 76548 160342 76560
rect 160554 76548 160560 76560
rect 160336 76520 160560 76548
rect 160336 76508 160342 76520
rect 160554 76508 160560 76520
rect 160612 76508 160618 76560
rect 161566 76508 161572 76560
rect 161624 76548 161630 76560
rect 162210 76548 162216 76560
rect 161624 76520 162216 76548
rect 161624 76508 161630 76520
rect 162210 76508 162216 76520
rect 162268 76508 162274 76560
rect 163038 76508 163044 76560
rect 163096 76548 163102 76560
rect 163406 76548 163412 76560
rect 163096 76520 163412 76548
rect 163096 76508 163102 76520
rect 163406 76508 163412 76520
rect 163464 76508 163470 76560
rect 164326 76508 164332 76560
rect 164384 76548 164390 76560
rect 164694 76548 164700 76560
rect 164384 76520 164700 76548
rect 164384 76508 164390 76520
rect 164694 76508 164700 76520
rect 164752 76508 164758 76560
rect 165706 76508 165712 76560
rect 165764 76548 165770 76560
rect 166718 76548 166724 76560
rect 165764 76520 166724 76548
rect 165764 76508 165770 76520
rect 166718 76508 166724 76520
rect 166776 76508 166782 76560
rect 167546 76508 167552 76560
rect 167604 76548 167610 76560
rect 167730 76548 167736 76560
rect 167604 76520 167736 76548
rect 167604 76508 167610 76520
rect 167730 76508 167736 76520
rect 167788 76508 167794 76560
rect 167914 76508 167920 76560
rect 167972 76548 167978 76560
rect 454034 76548 454040 76560
rect 167972 76520 454040 76548
rect 167972 76508 167978 76520
rect 454034 76508 454040 76520
rect 454092 76508 454098 76560
rect 172882 76480 172888 76492
rect 137986 76452 172888 76480
rect 172882 76440 172888 76452
rect 172940 76440 172946 76492
rect 172790 76412 172796 76424
rect 123536 76384 128216 76412
rect 128326 76384 172796 76412
rect 123536 76372 123542 76384
rect 120902 76304 120908 76356
rect 120960 76344 120966 76356
rect 128326 76344 128354 76384
rect 172790 76372 172796 76384
rect 172848 76372 172854 76424
rect 120960 76316 128354 76344
rect 120960 76304 120966 76316
rect 131666 76304 131672 76356
rect 131724 76344 131730 76356
rect 132126 76344 132132 76356
rect 131724 76316 132132 76344
rect 131724 76304 131730 76316
rect 132126 76304 132132 76316
rect 132184 76304 132190 76356
rect 151906 76304 151912 76356
rect 151964 76344 151970 76356
rect 152274 76344 152280 76356
rect 151964 76316 152280 76344
rect 151964 76304 151970 76316
rect 152274 76304 152280 76316
rect 152332 76304 152338 76356
rect 154758 76304 154764 76356
rect 154816 76344 154822 76356
rect 155126 76344 155132 76356
rect 154816 76316 155132 76344
rect 154816 76304 154822 76316
rect 155126 76304 155132 76316
rect 155184 76304 155190 76356
rect 163222 76304 163228 76356
rect 163280 76344 163286 76356
rect 163866 76344 163872 76356
rect 163280 76316 163872 76344
rect 163280 76304 163286 76316
rect 163866 76304 163872 76316
rect 163924 76304 163930 76356
rect 164510 76304 164516 76356
rect 164568 76344 164574 76356
rect 165338 76344 165344 76356
rect 164568 76316 165344 76344
rect 164568 76304 164574 76316
rect 165338 76304 165344 76316
rect 165396 76304 165402 76356
rect 168374 76304 168380 76356
rect 168432 76344 168438 76356
rect 168742 76344 168748 76356
rect 168432 76316 168748 76344
rect 168432 76304 168438 76316
rect 168742 76304 168748 76316
rect 168800 76304 168806 76356
rect 169662 76304 169668 76356
rect 169720 76344 169726 76356
rect 172238 76344 172244 76356
rect 169720 76316 172244 76344
rect 169720 76304 169726 76316
rect 172238 76304 172244 76316
rect 172296 76304 172302 76356
rect 144730 76236 144736 76288
rect 144788 76276 144794 76288
rect 145190 76276 145196 76288
rect 144788 76248 145196 76276
rect 144788 76236 144794 76248
rect 145190 76236 145196 76248
rect 145248 76236 145254 76288
rect 154574 76236 154580 76288
rect 154632 76276 154638 76288
rect 162762 76276 162768 76288
rect 154632 76248 162768 76276
rect 154632 76236 154638 76248
rect 162762 76236 162768 76248
rect 162820 76236 162826 76288
rect 163038 76236 163044 76288
rect 163096 76276 163102 76288
rect 163682 76276 163688 76288
rect 163096 76248 163688 76276
rect 163096 76236 163102 76248
rect 163682 76236 163688 76248
rect 163740 76236 163746 76288
rect 164786 76236 164792 76288
rect 164844 76276 164850 76288
rect 172054 76276 172060 76288
rect 164844 76248 172060 76276
rect 164844 76236 164850 76248
rect 172054 76236 172060 76248
rect 172112 76236 172118 76288
rect 135346 76168 135352 76220
rect 135404 76208 135410 76220
rect 135990 76208 135996 76220
rect 135404 76180 135996 76208
rect 135404 76168 135410 76180
rect 135990 76168 135996 76180
rect 136048 76168 136054 76220
rect 143626 76168 143632 76220
rect 143684 76208 143690 76220
rect 148686 76208 148692 76220
rect 143684 76180 148692 76208
rect 143684 76168 143690 76180
rect 148686 76168 148692 76180
rect 148744 76168 148750 76220
rect 151998 76168 152004 76220
rect 152056 76208 152062 76220
rect 152274 76208 152280 76220
rect 152056 76180 152280 76208
rect 152056 76168 152062 76180
rect 152274 76168 152280 76180
rect 152332 76168 152338 76220
rect 154666 76168 154672 76220
rect 154724 76208 154730 76220
rect 155126 76208 155132 76220
rect 154724 76180 155132 76208
rect 154724 76168 154730 76180
rect 155126 76168 155132 76180
rect 155184 76168 155190 76220
rect 160554 76168 160560 76220
rect 160612 76208 160618 76220
rect 160922 76208 160928 76220
rect 160612 76180 160928 76208
rect 160612 76168 160618 76180
rect 160922 76168 160928 76180
rect 160980 76168 160986 76220
rect 142338 76100 142344 76152
rect 142396 76140 142402 76152
rect 145834 76140 145840 76152
rect 142396 76112 145840 76140
rect 142396 76100 142402 76112
rect 145834 76100 145840 76112
rect 145892 76100 145898 76152
rect 150526 76100 150532 76152
rect 150584 76140 150590 76152
rect 158438 76140 158444 76152
rect 150584 76112 158444 76140
rect 150584 76100 150590 76112
rect 158438 76100 158444 76112
rect 158496 76100 158502 76152
rect 160370 76100 160376 76152
rect 160428 76140 160434 76152
rect 160738 76140 160744 76152
rect 160428 76112 160744 76140
rect 160428 76100 160434 76112
rect 160738 76100 160744 76112
rect 160796 76100 160802 76152
rect 142430 76032 142436 76084
rect 142488 76072 142494 76084
rect 142614 76072 142620 76084
rect 142488 76044 142620 76072
rect 142488 76032 142494 76044
rect 142614 76032 142620 76044
rect 142672 76032 142678 76084
rect 143718 76032 143724 76084
rect 143776 76072 143782 76084
rect 144270 76072 144276 76084
rect 143776 76044 144276 76072
rect 143776 76032 143782 76044
rect 144270 76032 144276 76044
rect 144328 76032 144334 76084
rect 145098 76032 145104 76084
rect 145156 76072 145162 76084
rect 145374 76072 145380 76084
rect 145156 76044 145380 76072
rect 145156 76032 145162 76044
rect 145374 76032 145380 76044
rect 145432 76032 145438 76084
rect 137646 75964 137652 76016
rect 137704 76004 137710 76016
rect 144638 76004 144644 76016
rect 137704 75976 144644 76004
rect 137704 75964 137710 75976
rect 144638 75964 144644 75976
rect 144696 75964 144702 76016
rect 144914 75964 144920 76016
rect 144972 76004 144978 76016
rect 145742 76004 145748 76016
rect 144972 75976 145748 76004
rect 144972 75964 144978 75976
rect 145742 75964 145748 75976
rect 145800 75964 145806 76016
rect 139394 75896 139400 75948
rect 139452 75936 139458 75948
rect 139578 75936 139584 75948
rect 139452 75908 139584 75936
rect 139452 75896 139458 75908
rect 139578 75896 139584 75908
rect 139636 75896 139642 75948
rect 139946 75896 139952 75948
rect 140004 75936 140010 75948
rect 140222 75936 140228 75948
rect 140004 75908 140228 75936
rect 140004 75896 140010 75908
rect 140222 75896 140228 75908
rect 140280 75896 140286 75948
rect 141142 75896 141148 75948
rect 141200 75936 141206 75948
rect 141602 75936 141608 75948
rect 141200 75908 141608 75936
rect 141200 75896 141206 75908
rect 141602 75896 141608 75908
rect 141660 75896 141666 75948
rect 143626 75896 143632 75948
rect 143684 75936 143690 75948
rect 143994 75936 144000 75948
rect 143684 75908 144000 75936
rect 143684 75896 143690 75908
rect 143994 75896 144000 75908
rect 144052 75896 144058 75948
rect 145374 75896 145380 75948
rect 145432 75936 145438 75948
rect 145650 75936 145656 75948
rect 145432 75908 145656 75936
rect 145432 75896 145438 75908
rect 145650 75896 145656 75908
rect 145708 75896 145714 75948
rect 157610 75896 157616 75948
rect 157668 75936 157674 75948
rect 158070 75936 158076 75948
rect 157668 75908 158076 75936
rect 157668 75896 157674 75908
rect 158070 75896 158076 75908
rect 158128 75896 158134 75948
rect 161566 75896 161572 75948
rect 161624 75936 161630 75948
rect 162026 75936 162032 75948
rect 161624 75908 162032 75936
rect 161624 75896 161630 75908
rect 162026 75896 162032 75908
rect 162084 75896 162090 75948
rect 169018 75896 169024 75948
rect 169076 75936 169082 75948
rect 170674 75936 170680 75948
rect 169076 75908 170680 75936
rect 169076 75896 169082 75908
rect 170674 75896 170680 75908
rect 170732 75896 170738 75948
rect 125686 75828 125692 75880
rect 125744 75868 125750 75880
rect 126238 75868 126244 75880
rect 125744 75840 126244 75868
rect 125744 75828 125750 75840
rect 126238 75828 126244 75840
rect 126296 75828 126302 75880
rect 140958 75828 140964 75880
rect 141016 75868 141022 75880
rect 141510 75868 141516 75880
rect 141016 75840 141516 75868
rect 141016 75828 141022 75840
rect 141510 75828 141516 75840
rect 141568 75828 141574 75880
rect 142154 75828 142160 75880
rect 142212 75868 142218 75880
rect 142798 75868 142804 75880
rect 142212 75840 142804 75868
rect 142212 75828 142218 75840
rect 142798 75828 142804 75840
rect 142856 75828 142862 75880
rect 143718 75828 143724 75880
rect 143776 75868 143782 75880
rect 144454 75868 144460 75880
rect 143776 75840 144460 75868
rect 143776 75828 143782 75840
rect 144454 75828 144460 75840
rect 144512 75828 144518 75880
rect 147766 75828 147772 75880
rect 147824 75868 147830 75880
rect 148410 75868 148416 75880
rect 147824 75840 148416 75868
rect 147824 75828 147830 75840
rect 148410 75828 148416 75840
rect 148468 75828 148474 75880
rect 155770 75828 155776 75880
rect 155828 75868 155834 75880
rect 156966 75868 156972 75880
rect 155828 75840 156972 75868
rect 155828 75828 155834 75840
rect 156966 75828 156972 75840
rect 157024 75828 157030 75880
rect 169846 75828 169852 75880
rect 169904 75868 169910 75880
rect 170490 75868 170496 75880
rect 169904 75840 170496 75868
rect 169904 75828 169910 75840
rect 170490 75828 170496 75840
rect 170548 75828 170554 75880
rect 139670 75760 139676 75812
rect 139728 75800 139734 75812
rect 140314 75800 140320 75812
rect 139728 75772 140320 75800
rect 139728 75760 139734 75772
rect 140314 75760 140320 75772
rect 140372 75760 140378 75812
rect 142522 75760 142528 75812
rect 142580 75800 142586 75812
rect 142706 75800 142712 75812
rect 142580 75772 142712 75800
rect 142580 75760 142586 75772
rect 142706 75760 142712 75772
rect 142764 75760 142770 75812
rect 143994 75760 144000 75812
rect 144052 75800 144058 75812
rect 144546 75800 144552 75812
rect 144052 75772 144552 75800
rect 144052 75760 144058 75772
rect 144546 75760 144552 75772
rect 144604 75760 144610 75812
rect 148042 75760 148048 75812
rect 148100 75800 148106 75812
rect 148594 75800 148600 75812
rect 148100 75772 148600 75800
rect 148100 75760 148106 75772
rect 148594 75760 148600 75772
rect 148652 75760 148658 75812
rect 126974 75692 126980 75744
rect 127032 75732 127038 75744
rect 134978 75732 134984 75744
rect 127032 75704 134984 75732
rect 127032 75692 127038 75704
rect 134978 75692 134984 75704
rect 135036 75692 135042 75744
rect 135990 75692 135996 75744
rect 136048 75732 136054 75744
rect 136542 75732 136548 75744
rect 136048 75704 136548 75732
rect 136048 75692 136054 75704
rect 136542 75692 136548 75704
rect 136600 75692 136606 75744
rect 139578 75692 139584 75744
rect 139636 75732 139642 75744
rect 140130 75732 140136 75744
rect 139636 75704 140136 75732
rect 139636 75692 139642 75704
rect 140130 75692 140136 75704
rect 140188 75692 140194 75744
rect 158990 75692 158996 75744
rect 159048 75732 159054 75744
rect 164786 75732 164792 75744
rect 159048 75704 164792 75732
rect 159048 75692 159054 75704
rect 164786 75692 164792 75704
rect 164844 75692 164850 75744
rect 130010 75624 130016 75676
rect 130068 75664 130074 75676
rect 130654 75664 130660 75676
rect 130068 75636 130660 75664
rect 130068 75624 130074 75636
rect 130654 75624 130660 75636
rect 130712 75624 130718 75676
rect 132678 75624 132684 75676
rect 132736 75664 132742 75676
rect 133598 75664 133604 75676
rect 132736 75636 133604 75664
rect 132736 75624 132742 75636
rect 133598 75624 133604 75636
rect 133656 75624 133662 75676
rect 158254 75624 158260 75676
rect 158312 75664 158318 75676
rect 158312 75636 169754 75664
rect 158312 75624 158318 75636
rect 122190 75556 122196 75608
rect 122248 75596 122254 75608
rect 130470 75596 130476 75608
rect 122248 75568 130476 75596
rect 122248 75556 122254 75568
rect 130470 75556 130476 75568
rect 130528 75556 130534 75608
rect 159542 75556 159548 75608
rect 159600 75596 159606 75608
rect 169726 75596 169754 75636
rect 396074 75596 396080 75608
rect 159600 75568 160094 75596
rect 169726 75568 396080 75596
rect 159600 75556 159606 75568
rect 121454 75420 121460 75472
rect 121512 75460 121518 75472
rect 126974 75460 126980 75472
rect 121512 75432 126980 75460
rect 121512 75420 121518 75432
rect 126974 75420 126980 75432
rect 127032 75420 127038 75472
rect 160066 75460 160094 75568
rect 396074 75556 396080 75568
rect 396132 75556 396138 75608
rect 164786 75488 164792 75540
rect 164844 75528 164850 75540
rect 431954 75528 431960 75540
rect 164844 75500 431960 75528
rect 164844 75488 164850 75500
rect 431954 75488 431960 75500
rect 432012 75488 432018 75540
rect 438854 75460 438860 75472
rect 160066 75432 438860 75460
rect 438854 75420 438860 75432
rect 438912 75420 438918 75472
rect 51074 75352 51080 75404
rect 51132 75392 51138 75404
rect 128722 75392 128728 75404
rect 51132 75364 128728 75392
rect 51132 75352 51138 75364
rect 128722 75352 128728 75364
rect 128780 75352 128786 75404
rect 138014 75352 138020 75404
rect 138072 75392 138078 75404
rect 138566 75392 138572 75404
rect 138072 75364 138572 75392
rect 138072 75352 138078 75364
rect 138566 75352 138572 75364
rect 138624 75352 138630 75404
rect 146754 75352 146760 75404
rect 146812 75392 146818 75404
rect 147214 75392 147220 75404
rect 146812 75364 147220 75392
rect 146812 75352 146818 75364
rect 147214 75352 147220 75364
rect 147272 75352 147278 75404
rect 161842 75352 161848 75404
rect 161900 75392 161906 75404
rect 467834 75392 467840 75404
rect 161900 75364 467840 75392
rect 161900 75352 161906 75364
rect 467834 75352 467840 75364
rect 467892 75352 467898 75404
rect 107654 75284 107660 75336
rect 107712 75324 107718 75336
rect 132494 75324 132500 75336
rect 107712 75296 132500 75324
rect 107712 75284 107718 75296
rect 132494 75284 132500 75296
rect 132552 75284 132558 75336
rect 157334 75284 157340 75336
rect 157392 75324 157398 75336
rect 157978 75324 157984 75336
rect 157392 75296 157984 75324
rect 157392 75284 157398 75296
rect 157978 75284 157984 75296
rect 158036 75284 158042 75336
rect 167822 75284 167828 75336
rect 167880 75324 167886 75336
rect 490006 75324 490012 75336
rect 167880 75296 490012 75324
rect 167880 75284 167886 75296
rect 490006 75284 490012 75296
rect 490064 75284 490070 75336
rect 42794 75216 42800 75268
rect 42852 75256 42858 75268
rect 42852 75228 128354 75256
rect 42852 75216 42858 75228
rect 6914 75148 6920 75200
rect 6972 75188 6978 75200
rect 125686 75188 125692 75200
rect 6972 75160 125692 75188
rect 6972 75148 6978 75160
rect 125686 75148 125692 75160
rect 125744 75148 125750 75200
rect 125962 75148 125968 75200
rect 126020 75188 126026 75200
rect 126238 75188 126244 75200
rect 126020 75160 126244 75188
rect 126020 75148 126026 75160
rect 126238 75148 126244 75160
rect 126296 75148 126302 75200
rect 127250 75148 127256 75200
rect 127308 75188 127314 75200
rect 128170 75188 128176 75200
rect 127308 75160 128176 75188
rect 127308 75148 127314 75160
rect 128170 75148 128176 75160
rect 128228 75148 128234 75200
rect 128326 75188 128354 75228
rect 128538 75216 128544 75268
rect 128596 75256 128602 75268
rect 129274 75256 129280 75268
rect 128596 75228 129280 75256
rect 128596 75216 128602 75228
rect 129274 75216 129280 75228
rect 129332 75216 129338 75268
rect 130286 75216 130292 75268
rect 130344 75256 130350 75268
rect 131022 75256 131028 75268
rect 130344 75228 131028 75256
rect 130344 75216 130350 75228
rect 131022 75216 131028 75228
rect 131080 75216 131086 75268
rect 138382 75216 138388 75268
rect 138440 75256 138446 75268
rect 138566 75256 138572 75268
rect 138440 75228 138572 75256
rect 138440 75216 138446 75228
rect 138566 75216 138572 75228
rect 138624 75216 138630 75268
rect 140866 75216 140872 75268
rect 140924 75256 140930 75268
rect 141786 75256 141792 75268
rect 140924 75228 141792 75256
rect 140924 75216 140930 75228
rect 141786 75216 141792 75228
rect 141844 75216 141850 75268
rect 146478 75216 146484 75268
rect 146536 75256 146542 75268
rect 146754 75256 146760 75268
rect 146536 75228 146760 75256
rect 146536 75216 146542 75228
rect 146754 75216 146760 75228
rect 146812 75216 146818 75268
rect 149330 75216 149336 75268
rect 149388 75256 149394 75268
rect 149698 75256 149704 75268
rect 149388 75228 149704 75256
rect 149388 75216 149394 75228
rect 149698 75216 149704 75228
rect 149756 75216 149762 75268
rect 166442 75216 166448 75268
rect 166500 75256 166506 75268
rect 499574 75256 499580 75268
rect 166500 75228 499580 75256
rect 166500 75216 166506 75228
rect 499574 75216 499580 75228
rect 499632 75216 499638 75268
rect 128906 75188 128912 75200
rect 128326 75160 128912 75188
rect 128906 75148 128912 75160
rect 128964 75148 128970 75200
rect 131298 75148 131304 75200
rect 131356 75188 131362 75200
rect 132034 75188 132040 75200
rect 131356 75160 132040 75188
rect 131356 75148 131362 75160
rect 132034 75148 132040 75160
rect 132092 75148 132098 75200
rect 146570 75148 146576 75200
rect 146628 75188 146634 75200
rect 146846 75188 146852 75200
rect 146628 75160 146852 75188
rect 146628 75148 146634 75160
rect 146846 75148 146852 75160
rect 146904 75148 146910 75200
rect 160186 75148 160192 75200
rect 160244 75188 160250 75200
rect 160830 75188 160836 75200
rect 160244 75160 160836 75188
rect 160244 75148 160250 75160
rect 160830 75148 160836 75160
rect 160888 75148 160894 75200
rect 169294 75148 169300 75200
rect 169352 75188 169358 75200
rect 564434 75188 564440 75200
rect 169352 75160 564440 75188
rect 169352 75148 169358 75160
rect 564434 75148 564440 75160
rect 564492 75148 564498 75200
rect 125870 75080 125876 75132
rect 125928 75120 125934 75132
rect 126606 75120 126612 75132
rect 125928 75092 126612 75120
rect 125928 75080 125934 75092
rect 126606 75080 126612 75092
rect 126664 75080 126670 75132
rect 127342 75080 127348 75132
rect 127400 75120 127406 75132
rect 128262 75120 128268 75132
rect 127400 75092 128268 75120
rect 127400 75080 127406 75092
rect 128262 75080 128268 75092
rect 128320 75080 128326 75132
rect 128722 75080 128728 75132
rect 128780 75120 128786 75132
rect 129642 75120 129648 75132
rect 128780 75092 129648 75120
rect 128780 75080 128786 75092
rect 129642 75080 129648 75092
rect 129700 75080 129706 75132
rect 138198 75080 138204 75132
rect 138256 75120 138262 75132
rect 138382 75120 138388 75132
rect 138256 75092 138388 75120
rect 138256 75080 138262 75092
rect 138382 75080 138388 75092
rect 138440 75080 138446 75132
rect 142522 75080 142528 75132
rect 142580 75120 142586 75132
rect 142890 75120 142896 75132
rect 142580 75092 142896 75120
rect 142580 75080 142586 75092
rect 142890 75080 142896 75092
rect 142948 75080 142954 75132
rect 170214 75080 170220 75132
rect 170272 75120 170278 75132
rect 170766 75120 170772 75132
rect 170272 75092 170772 75120
rect 170272 75080 170278 75092
rect 170766 75080 170772 75092
rect 170824 75080 170830 75132
rect 125962 75012 125968 75064
rect 126020 75052 126026 75064
rect 126882 75052 126888 75064
rect 126020 75024 126888 75052
rect 126020 75012 126026 75024
rect 126882 75012 126888 75024
rect 126940 75012 126946 75064
rect 128354 75012 128360 75064
rect 128412 75052 128418 75064
rect 133414 75052 133420 75064
rect 128412 75024 133420 75052
rect 128412 75012 128418 75024
rect 133414 75012 133420 75024
rect 133472 75012 133478 75064
rect 125686 74944 125692 74996
rect 125744 74984 125750 74996
rect 126790 74984 126796 74996
rect 125744 74956 126796 74984
rect 125744 74944 125750 74956
rect 126790 74944 126796 74956
rect 126848 74944 126854 74996
rect 128446 74944 128452 74996
rect 128504 74984 128510 74996
rect 129550 74984 129556 74996
rect 128504 74956 129556 74984
rect 128504 74944 128510 74956
rect 129550 74944 129556 74956
rect 129608 74944 129614 74996
rect 138198 74944 138204 74996
rect 138256 74984 138262 74996
rect 138658 74984 138664 74996
rect 138256 74956 138664 74984
rect 138256 74944 138262 74956
rect 138658 74944 138664 74956
rect 138716 74944 138722 74996
rect 164694 74944 164700 74996
rect 164752 74984 164758 74996
rect 164970 74984 164976 74996
rect 164752 74956 164976 74984
rect 164752 74944 164758 74956
rect 164970 74944 164976 74956
rect 165028 74944 165034 74996
rect 146478 74876 146484 74928
rect 146536 74916 146542 74928
rect 147122 74916 147128 74928
rect 146536 74888 147128 74916
rect 146536 74876 146542 74888
rect 147122 74876 147128 74888
rect 147180 74876 147186 74928
rect 155862 74808 155868 74860
rect 155920 74848 155926 74860
rect 159634 74848 159640 74860
rect 155920 74820 159640 74848
rect 155920 74808 155926 74820
rect 159634 74808 159640 74820
rect 159692 74808 159698 74860
rect 146294 74740 146300 74792
rect 146352 74780 146358 74792
rect 147306 74780 147312 74792
rect 146352 74752 147312 74780
rect 146352 74740 146358 74752
rect 147306 74740 147312 74752
rect 147364 74740 147370 74792
rect 161842 74740 161848 74792
rect 161900 74780 161906 74792
rect 162302 74780 162308 74792
rect 161900 74752 162308 74780
rect 161900 74740 161906 74752
rect 162302 74740 162308 74752
rect 162360 74740 162366 74792
rect 147674 74604 147680 74656
rect 147732 74644 147738 74656
rect 148502 74644 148508 74656
rect 147732 74616 148508 74644
rect 147732 74604 147738 74616
rect 148502 74604 148508 74616
rect 148560 74604 148566 74656
rect 154574 74536 154580 74588
rect 154632 74576 154638 74588
rect 155494 74576 155500 74588
rect 154632 74548 155500 74576
rect 154632 74536 154638 74548
rect 155494 74536 155500 74548
rect 155552 74536 155558 74588
rect 168558 74468 168564 74520
rect 168616 74508 168622 74520
rect 173342 74508 173348 74520
rect 168616 74480 173348 74508
rect 168616 74468 168622 74480
rect 173342 74468 173348 74480
rect 173400 74468 173406 74520
rect 153286 74400 153292 74452
rect 153344 74440 153350 74452
rect 153838 74440 153844 74452
rect 153344 74412 153844 74440
rect 153344 74400 153350 74412
rect 153838 74400 153844 74412
rect 153896 74400 153902 74452
rect 150434 74332 150440 74384
rect 150492 74372 150498 74384
rect 156874 74372 156880 74384
rect 150492 74344 156880 74372
rect 150492 74332 150498 74344
rect 156874 74332 156880 74344
rect 156932 74332 156938 74384
rect 145466 74196 145472 74248
rect 145524 74236 145530 74248
rect 209774 74236 209780 74248
rect 145524 74208 209780 74236
rect 145524 74196 145530 74208
rect 209774 74196 209780 74208
rect 209832 74196 209838 74248
rect 145834 74128 145840 74180
rect 145892 74168 145898 74180
rect 216674 74168 216680 74180
rect 145892 74140 216680 74168
rect 145892 74128 145898 74140
rect 216674 74128 216680 74140
rect 216732 74128 216738 74180
rect 118694 74060 118700 74112
rect 118752 74100 118758 74112
rect 134702 74100 134708 74112
rect 118752 74072 134708 74100
rect 118752 74060 118758 74072
rect 134702 74060 134708 74072
rect 134760 74060 134766 74112
rect 142982 74060 142988 74112
rect 143040 74100 143046 74112
rect 223574 74100 223580 74112
rect 143040 74072 223580 74100
rect 143040 74060 143046 74072
rect 223574 74060 223580 74072
rect 223632 74060 223638 74112
rect 93946 73992 93952 74044
rect 94004 74032 94010 74044
rect 133138 74032 133144 74044
rect 94004 74004 133144 74032
rect 94004 73992 94010 74004
rect 133138 73992 133144 74004
rect 133196 73992 133202 74044
rect 145006 73992 145012 74044
rect 145064 74032 145070 74044
rect 145466 74032 145472 74044
rect 145064 74004 145472 74032
rect 145064 73992 145070 74004
rect 145466 73992 145472 74004
rect 145524 73992 145530 74044
rect 147398 73992 147404 74044
rect 147456 74032 147462 74044
rect 251174 74032 251180 74044
rect 147456 74004 251180 74032
rect 147456 73992 147462 74004
rect 251174 73992 251180 74004
rect 251232 73992 251238 74044
rect 64874 73924 64880 73976
rect 64932 73964 64938 73976
rect 129734 73964 129740 73976
rect 64932 73936 129740 73964
rect 64932 73924 64938 73936
rect 129734 73924 129740 73936
rect 129792 73924 129798 73976
rect 142246 73924 142252 73976
rect 142304 73964 142310 73976
rect 143074 73964 143080 73976
rect 142304 73936 143080 73964
rect 142304 73924 142310 73936
rect 143074 73924 143080 73936
rect 143132 73924 143138 73976
rect 157702 73924 157708 73976
rect 157760 73964 157766 73976
rect 158162 73964 158168 73976
rect 157760 73936 158168 73964
rect 157760 73924 157766 73936
rect 158162 73924 158168 73936
rect 158220 73924 158226 73976
rect 158438 73924 158444 73976
rect 158496 73964 158502 73976
rect 318794 73964 318800 73976
rect 158496 73936 318800 73964
rect 158496 73924 158502 73936
rect 318794 73924 318800 73936
rect 318852 73924 318858 73976
rect 27614 73856 27620 73908
rect 27672 73896 27678 73908
rect 127802 73896 127808 73908
rect 27672 73868 127808 73896
rect 27672 73856 27678 73868
rect 127802 73856 127808 73868
rect 127860 73856 127866 73908
rect 135714 73856 135720 73908
rect 135772 73896 135778 73908
rect 136358 73896 136364 73908
rect 135772 73868 136364 73896
rect 135772 73856 135778 73868
rect 136358 73856 136364 73868
rect 136416 73856 136422 73908
rect 145006 73856 145012 73908
rect 145064 73896 145070 73908
rect 146018 73896 146024 73908
rect 145064 73868 146024 73896
rect 145064 73856 145070 73868
rect 146018 73856 146024 73868
rect 146076 73856 146082 73908
rect 151998 73856 152004 73908
rect 152056 73896 152062 73908
rect 152642 73896 152648 73908
rect 152056 73868 152648 73896
rect 152056 73856 152062 73868
rect 152642 73856 152648 73868
rect 152700 73856 152706 73908
rect 153102 73856 153108 73908
rect 153160 73896 153166 73908
rect 354674 73896 354680 73908
rect 153160 73868 354680 73896
rect 153160 73856 153166 73868
rect 354674 73856 354680 73868
rect 354732 73856 354738 73908
rect 26234 73788 26240 73840
rect 26292 73828 26298 73840
rect 127894 73828 127900 73840
rect 26292 73800 127900 73828
rect 26292 73788 26298 73800
rect 127894 73788 127900 73800
rect 127952 73788 127958 73840
rect 143534 73788 143540 73840
rect 143592 73828 143598 73840
rect 144362 73828 144368 73840
rect 143592 73800 144368 73828
rect 143592 73788 143598 73800
rect 144362 73788 144368 73800
rect 144420 73788 144426 73840
rect 164786 73788 164792 73840
rect 164844 73828 164850 73840
rect 165062 73828 165068 73840
rect 164844 73800 165068 73828
rect 164844 73788 164850 73800
rect 165062 73788 165068 73800
rect 165120 73788 165126 73840
rect 165154 73788 165160 73840
rect 165212 73828 165218 73840
rect 375374 73828 375380 73840
rect 165212 73800 375380 73828
rect 165212 73788 165218 73800
rect 375374 73788 375380 73800
rect 375432 73788 375438 73840
rect 150526 73720 150532 73772
rect 150584 73760 150590 73772
rect 151262 73760 151268 73772
rect 150584 73732 151268 73760
rect 150584 73720 150590 73732
rect 151262 73720 151268 73732
rect 151320 73720 151326 73772
rect 158990 73720 158996 73772
rect 159048 73760 159054 73772
rect 159818 73760 159824 73772
rect 159048 73732 159824 73760
rect 159048 73720 159054 73732
rect 159818 73720 159824 73732
rect 159876 73720 159882 73772
rect 161658 73584 161664 73636
rect 161716 73624 161722 73636
rect 162118 73624 162124 73636
rect 161716 73596 162124 73624
rect 161716 73584 161722 73596
rect 162118 73584 162124 73596
rect 162176 73584 162182 73636
rect 137462 73448 137468 73500
rect 137520 73488 137526 73500
rect 138934 73488 138940 73500
rect 137520 73460 138940 73488
rect 137520 73448 137526 73460
rect 138934 73448 138940 73460
rect 138992 73448 138998 73500
rect 155954 73448 155960 73500
rect 156012 73488 156018 73500
rect 156506 73488 156512 73500
rect 156012 73460 156512 73488
rect 156012 73448 156018 73460
rect 156506 73448 156512 73460
rect 156564 73448 156570 73500
rect 154758 73244 154764 73296
rect 154816 73284 154822 73296
rect 155402 73284 155408 73296
rect 154816 73256 155408 73284
rect 154816 73244 154822 73256
rect 155402 73244 155408 73256
rect 155460 73244 155466 73296
rect 137370 73176 137376 73228
rect 137428 73216 137434 73228
rect 142982 73216 142988 73228
rect 137428 73188 142988 73216
rect 137428 73176 137434 73188
rect 142982 73176 142988 73188
rect 143040 73176 143046 73228
rect 177298 73108 177304 73160
rect 177356 73148 177362 73160
rect 580166 73148 580172 73160
rect 177356 73120 580172 73148
rect 177356 73108 177362 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 158714 72904 158720 72956
rect 158772 72944 158778 72956
rect 158990 72944 158996 72956
rect 158772 72916 158996 72944
rect 158772 72904 158778 72916
rect 158990 72904 158996 72916
rect 159048 72904 159054 72956
rect 148318 72632 148324 72684
rect 148376 72672 148382 72684
rect 291194 72672 291200 72684
rect 148376 72644 291200 72672
rect 148376 72632 148382 72644
rect 291194 72632 291200 72644
rect 291252 72632 291258 72684
rect 149882 72564 149888 72616
rect 149940 72604 149946 72616
rect 311894 72604 311900 72616
rect 149940 72576 311900 72604
rect 149940 72564 149946 72576
rect 311894 72564 311900 72576
rect 311952 72564 311958 72616
rect 152734 72496 152740 72548
rect 152792 72536 152798 72548
rect 340874 72536 340880 72548
rect 152792 72508 340880 72536
rect 152792 72496 152798 72508
rect 340874 72496 340880 72508
rect 340932 72496 340938 72548
rect 153194 72428 153200 72480
rect 153252 72468 153258 72480
rect 357434 72468 357440 72480
rect 153252 72440 357440 72468
rect 153252 72428 153258 72440
rect 357434 72428 357440 72440
rect 357492 72428 357498 72480
rect 165246 72360 165252 72412
rect 165304 72400 165310 72412
rect 171870 72400 171876 72412
rect 165304 72372 171876 72400
rect 165304 72360 165310 72372
rect 171870 72360 171876 72372
rect 171928 72360 171934 72412
rect 168558 72292 168564 72344
rect 168616 72332 168622 72344
rect 169110 72332 169116 72344
rect 168616 72304 169116 72332
rect 168616 72292 168622 72304
rect 169110 72292 169116 72304
rect 169168 72292 169174 72344
rect 167086 72088 167092 72140
rect 167144 72128 167150 72140
rect 168006 72128 168012 72140
rect 167144 72100 168012 72128
rect 167144 72088 167150 72100
rect 168006 72088 168012 72100
rect 168064 72088 168070 72140
rect 3418 71680 3424 71732
rect 3476 71720 3482 71732
rect 179598 71720 179604 71732
rect 3476 71692 179604 71720
rect 3476 71680 3482 71692
rect 179598 71680 179604 71692
rect 179656 71680 179662 71732
rect 78674 71000 78680 71052
rect 78732 71040 78738 71052
rect 131758 71040 131764 71052
rect 78732 71012 131764 71040
rect 78732 71000 78738 71012
rect 131758 71000 131764 71012
rect 131816 71000 131822 71052
rect 138842 71000 138848 71052
rect 138900 71040 138906 71052
rect 152550 71040 152556 71052
rect 138900 71012 152556 71040
rect 138900 71000 138906 71012
rect 152550 71000 152556 71012
rect 152608 71000 152614 71052
rect 157334 71000 157340 71052
rect 157392 71040 157398 71052
rect 284386 71040 284392 71052
rect 157392 71012 284392 71040
rect 157392 71000 157398 71012
rect 284386 71000 284392 71012
rect 284444 71000 284450 71052
rect 138658 70320 138664 70372
rect 138716 70360 138722 70372
rect 142798 70360 142804 70372
rect 138716 70332 142804 70360
rect 138716 70320 138722 70332
rect 142798 70320 142804 70332
rect 142856 70320 142862 70372
rect 141510 70048 141516 70100
rect 141568 70088 141574 70100
rect 209866 70088 209872 70100
rect 141568 70060 209872 70088
rect 141568 70048 141574 70060
rect 209866 70048 209872 70060
rect 209924 70048 209930 70100
rect 155310 69980 155316 70032
rect 155368 70020 155374 70032
rect 382274 70020 382280 70032
rect 155368 69992 382280 70020
rect 155368 69980 155374 69992
rect 382274 69980 382280 69992
rect 382332 69980 382338 70032
rect 156782 69912 156788 69964
rect 156840 69952 156846 69964
rect 390554 69952 390560 69964
rect 156840 69924 390560 69952
rect 156840 69912 156846 69924
rect 390554 69912 390560 69924
rect 390612 69912 390618 69964
rect 171686 69844 171692 69896
rect 171744 69884 171750 69896
rect 426434 69884 426440 69896
rect 171744 69856 426440 69884
rect 171744 69844 171750 69856
rect 426434 69844 426440 69856
rect 426492 69844 426498 69896
rect 164878 69776 164884 69828
rect 164936 69816 164942 69828
rect 505094 69816 505100 69828
rect 164936 69788 505100 69816
rect 164936 69776 164942 69788
rect 505094 69776 505100 69788
rect 505152 69776 505158 69828
rect 166626 69708 166632 69760
rect 166684 69748 166690 69760
rect 518894 69748 518900 69760
rect 166684 69720 518900 69748
rect 166684 69708 166690 69720
rect 518894 69708 518900 69720
rect 518952 69708 518958 69760
rect 170306 69640 170312 69692
rect 170364 69680 170370 69692
rect 568574 69680 568580 69692
rect 170364 69652 568580 69680
rect 170364 69640 170370 69652
rect 568574 69640 568580 69652
rect 568632 69640 568638 69692
rect 170214 68960 170220 69012
rect 170272 69000 170278 69012
rect 171686 69000 171692 69012
rect 170272 68972 171692 69000
rect 170272 68960 170278 68972
rect 171686 68960 171692 68972
rect 171744 68960 171750 69012
rect 140038 68620 140044 68672
rect 140096 68660 140102 68672
rect 184934 68660 184940 68672
rect 140096 68632 184940 68660
rect 140096 68620 140102 68632
rect 184934 68620 184940 68632
rect 184992 68620 184998 68672
rect 142706 68552 142712 68604
rect 142764 68592 142770 68604
rect 218054 68592 218060 68604
rect 142764 68564 218060 68592
rect 142764 68552 142770 68564
rect 218054 68552 218060 68564
rect 218112 68552 218118 68604
rect 156874 68484 156880 68536
rect 156932 68524 156938 68536
rect 320174 68524 320180 68536
rect 156932 68496 320180 68524
rect 156932 68484 156938 68496
rect 320174 68484 320180 68496
rect 320232 68484 320238 68536
rect 153746 68416 153752 68468
rect 153804 68456 153810 68468
rect 362954 68456 362960 68468
rect 153804 68428 362960 68456
rect 153804 68416 153810 68428
rect 362954 68416 362960 68428
rect 363012 68416 363018 68468
rect 159266 68348 159272 68400
rect 159324 68388 159330 68400
rect 427814 68388 427820 68400
rect 159324 68360 427820 68388
rect 159324 68348 159330 68360
rect 427814 68348 427820 68360
rect 427872 68348 427878 68400
rect 169478 68280 169484 68332
rect 169536 68320 169542 68332
rect 564526 68320 564532 68332
rect 169536 68292 564532 68320
rect 169536 68280 169542 68292
rect 564526 68280 564532 68292
rect 564584 68280 564590 68332
rect 139946 67396 139952 67448
rect 140004 67436 140010 67448
rect 189074 67436 189080 67448
rect 140004 67408 189080 67436
rect 140004 67396 140010 67408
rect 189074 67396 189080 67408
rect 189132 67396 189138 67448
rect 147122 67328 147128 67380
rect 147180 67368 147186 67380
rect 270494 67368 270500 67380
rect 147180 67340 270500 67368
rect 147180 67328 147186 67340
rect 270494 67328 270500 67340
rect 270552 67328 270558 67380
rect 149698 67260 149704 67312
rect 149756 67300 149762 67312
rect 306374 67300 306380 67312
rect 149756 67272 306380 67300
rect 149756 67260 149762 67272
rect 306374 67260 306380 67272
rect 306432 67260 306438 67312
rect 161014 67192 161020 67244
rect 161072 67232 161078 67244
rect 347774 67232 347780 67244
rect 161072 67204 347780 67232
rect 161072 67192 161078 67204
rect 347774 67192 347780 67204
rect 347832 67192 347838 67244
rect 152458 67124 152464 67176
rect 152516 67164 152522 67176
rect 340966 67164 340972 67176
rect 152516 67136 340972 67164
rect 152516 67124 152522 67136
rect 340966 67124 340972 67136
rect 341024 67124 341030 67176
rect 159174 67056 159180 67108
rect 159232 67096 159238 67108
rect 437474 67096 437480 67108
rect 159232 67068 437480 67096
rect 159232 67056 159238 67068
rect 437474 67056 437480 67068
rect 437532 67056 437538 67108
rect 162026 66988 162032 67040
rect 162084 67028 162090 67040
rect 462314 67028 462320 67040
rect 162084 67000 462320 67028
rect 162084 66988 162090 67000
rect 462314 66988 462320 67000
rect 462372 66988 462378 67040
rect 167730 66920 167736 66972
rect 167788 66960 167794 66972
rect 539594 66960 539600 66972
rect 167788 66932 539600 66960
rect 167788 66920 167794 66932
rect 539594 66920 539600 66932
rect 539652 66920 539658 66972
rect 167638 66852 167644 66904
rect 167696 66892 167702 66904
rect 543734 66892 543740 66904
rect 167696 66864 543740 66892
rect 167696 66852 167702 66864
rect 543734 66852 543740 66864
rect 543792 66852 543798 66904
rect 137278 66172 137284 66224
rect 137336 66212 137342 66224
rect 140038 66212 140044 66224
rect 137336 66184 140044 66212
rect 137336 66172 137342 66184
rect 140038 66172 140044 66184
rect 140096 66172 140102 66224
rect 138566 66104 138572 66156
rect 138624 66144 138630 66156
rect 141510 66144 141516 66156
rect 138624 66116 141516 66144
rect 138624 66104 138630 66116
rect 141510 66104 141516 66116
rect 141568 66104 141574 66156
rect 141418 65900 141424 65952
rect 141476 65940 141482 65952
rect 202874 65940 202880 65952
rect 141476 65912 202880 65940
rect 141476 65900 141482 65912
rect 202874 65900 202880 65912
rect 202932 65900 202938 65952
rect 141326 65832 141332 65884
rect 141384 65872 141390 65884
rect 207014 65872 207020 65884
rect 141384 65844 207020 65872
rect 141384 65832 141390 65844
rect 207014 65832 207020 65844
rect 207072 65832 207078 65884
rect 142614 65764 142620 65816
rect 142672 65804 142678 65816
rect 220814 65804 220820 65816
rect 142672 65776 220820 65804
rect 142672 65764 142678 65776
rect 220814 65764 220820 65776
rect 220872 65764 220878 65816
rect 145466 65696 145472 65748
rect 145524 65736 145530 65748
rect 251266 65736 251272 65748
rect 145524 65708 251272 65736
rect 145524 65696 145530 65708
rect 251266 65696 251272 65708
rect 251324 65696 251330 65748
rect 145558 65628 145564 65680
rect 145616 65668 145622 65680
rect 256694 65668 256700 65680
rect 145616 65640 256700 65668
rect 145616 65628 145622 65640
rect 256694 65628 256700 65640
rect 256752 65628 256758 65680
rect 153654 65560 153660 65612
rect 153712 65600 153718 65612
rect 358814 65600 358820 65612
rect 153712 65572 358820 65600
rect 153712 65560 153718 65572
rect 358814 65560 358820 65572
rect 358872 65560 358878 65612
rect 102226 65492 102232 65544
rect 102284 65532 102290 65544
rect 125318 65532 125324 65544
rect 102284 65504 125324 65532
rect 102284 65492 102290 65504
rect 125318 65492 125324 65504
rect 125376 65492 125382 65544
rect 155218 65492 155224 65544
rect 155276 65532 155282 65544
rect 376754 65532 376760 65544
rect 155276 65504 376760 65532
rect 155276 65492 155282 65504
rect 376754 65492 376760 65504
rect 376812 65492 376818 65544
rect 144270 64472 144276 64524
rect 144328 64512 144334 64524
rect 234614 64512 234620 64524
rect 144328 64484 234620 64512
rect 144328 64472 144334 64484
rect 234614 64472 234620 64484
rect 234672 64472 234678 64524
rect 144178 64404 144184 64456
rect 144236 64444 144242 64456
rect 238754 64444 238760 64456
rect 144236 64416 238760 64444
rect 144236 64404 144242 64416
rect 238754 64404 238760 64416
rect 238812 64404 238818 64456
rect 148226 64336 148232 64388
rect 148284 64376 148290 64388
rect 292574 64376 292580 64388
rect 148284 64348 292580 64376
rect 148284 64336 148290 64348
rect 292574 64336 292580 64348
rect 292632 64336 292638 64388
rect 152366 64268 152372 64320
rect 152424 64308 152430 64320
rect 338114 64308 338120 64320
rect 152424 64280 338120 64308
rect 152424 64268 152430 64280
rect 338114 64268 338120 64280
rect 338172 64268 338178 64320
rect 162210 64200 162216 64252
rect 162268 64240 162274 64252
rect 368474 64240 368480 64252
rect 162268 64212 368480 64240
rect 162268 64200 162274 64212
rect 368474 64200 368480 64212
rect 368532 64200 368538 64252
rect 169018 64132 169024 64184
rect 169076 64172 169082 64184
rect 561674 64172 561680 64184
rect 169076 64144 561680 64172
rect 169076 64132 169082 64144
rect 561674 64132 561680 64144
rect 561732 64132 561738 64184
rect 147030 63112 147036 63164
rect 147088 63152 147094 63164
rect 274634 63152 274640 63164
rect 147088 63124 274640 63152
rect 147088 63112 147094 63124
rect 274634 63112 274640 63124
rect 274692 63112 274698 63164
rect 149606 63044 149612 63096
rect 149664 63084 149670 63096
rect 309134 63084 309140 63096
rect 149664 63056 309140 63084
rect 149664 63044 149670 63056
rect 309134 63044 309140 63056
rect 309192 63044 309198 63096
rect 155126 62976 155132 63028
rect 155184 63016 155190 63028
rect 373994 63016 374000 63028
rect 155184 62988 374000 63016
rect 155184 62976 155190 62988
rect 373994 62976 374000 62988
rect 374052 62976 374058 63028
rect 157978 62908 157984 62960
rect 158036 62948 158042 62960
rect 408494 62948 408500 62960
rect 158036 62920 408500 62948
rect 158036 62908 158042 62920
rect 408494 62908 408500 62920
rect 408552 62908 408558 62960
rect 163590 62840 163596 62892
rect 163648 62880 163654 62892
rect 488534 62880 488540 62892
rect 163648 62852 488540 62880
rect 163648 62840 163654 62852
rect 488534 62840 488540 62852
rect 488592 62840 488598 62892
rect 168926 62772 168932 62824
rect 168984 62812 168990 62824
rect 557534 62812 557540 62824
rect 168984 62784 557540 62812
rect 168984 62772 168990 62784
rect 557534 62772 557540 62784
rect 557592 62772 557598 62824
rect 139854 61480 139860 61532
rect 139912 61520 139918 61532
rect 185026 61520 185032 61532
rect 139912 61492 185032 61520
rect 139912 61480 139918 61492
rect 185026 61480 185032 61492
rect 185084 61480 185090 61532
rect 157886 61412 157892 61464
rect 157944 61452 157950 61464
rect 412634 61452 412640 61464
rect 157944 61424 412640 61452
rect 157944 61412 157950 61424
rect 412634 61412 412640 61424
rect 412692 61412 412698 61464
rect 166350 61344 166356 61396
rect 166408 61384 166414 61396
rect 525794 61384 525800 61396
rect 166408 61356 525800 61384
rect 166408 61344 166414 61356
rect 525794 61344 525800 61356
rect 525852 61344 525858 61396
rect 118510 60664 118516 60716
rect 118568 60704 118574 60716
rect 580166 60704 580172 60716
rect 118568 60676 580172 60704
rect 118568 60664 118574 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 137186 59984 137192 60036
rect 137244 60024 137250 60036
rect 138658 60024 138664 60036
rect 137244 59996 138664 60024
rect 137244 59984 137250 59996
rect 138658 59984 138664 59996
rect 138716 59984 138722 60036
rect 159082 59984 159088 60036
rect 159140 60024 159146 60036
rect 433334 60024 433340 60036
rect 159140 59996 433340 60024
rect 159140 59984 159146 59996
rect 433334 59984 433340 59996
rect 433392 59984 433398 60036
rect 156506 58624 156512 58676
rect 156564 58664 156570 58676
rect 401594 58664 401600 58676
rect 156564 58636 401600 58664
rect 156564 58624 156570 58636
rect 401594 58624 401600 58636
rect 401652 58624 401658 58676
rect 163498 57264 163504 57316
rect 163556 57304 163562 57316
rect 481634 57304 481640 57316
rect 163556 57276 481640 57304
rect 163556 57264 163562 57276
rect 481634 57264 481640 57276
rect 481692 57264 481698 57316
rect 164786 57196 164792 57248
rect 164844 57236 164850 57248
rect 507854 57236 507860 57248
rect 164844 57208 507860 57236
rect 164844 57196 164850 57208
rect 507854 57196 507860 57208
rect 507912 57196 507918 57248
rect 95234 53048 95240 53100
rect 95292 53088 95298 53100
rect 125226 53088 125232 53100
rect 95292 53060 125232 53088
rect 95292 53048 95298 53060
rect 125226 53048 125232 53060
rect 125284 53048 125290 53100
rect 182818 46860 182824 46912
rect 182876 46900 182882 46912
rect 580166 46900 580172 46912
rect 182876 46872 580172 46900
rect 182876 46860 182882 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 139762 46180 139768 46232
rect 139820 46220 139826 46232
rect 180794 46220 180800 46232
rect 139820 46192 180800 46220
rect 139820 46180 139826 46192
rect 180794 46180 180800 46192
rect 180852 46180 180858 46232
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 174078 45540 174084 45552
rect 3476 45512 174084 45540
rect 3476 45500 3482 45512
rect 174078 45500 174084 45512
rect 174136 45500 174142 45552
rect 135990 44956 135996 45008
rect 136048 44996 136054 45008
rect 142614 44996 142620 45008
rect 136048 44968 142620 44996
rect 136048 44956 136054 44968
rect 142614 44956 142620 44968
rect 142672 44956 142678 45008
rect 70394 44888 70400 44940
rect 70452 44928 70458 44940
rect 130286 44928 130292 44940
rect 70452 44900 130292 44928
rect 70452 44888 70458 44900
rect 130286 44888 130292 44900
rect 130344 44888 130350 44940
rect 34514 44820 34520 44872
rect 34572 44860 34578 44872
rect 127342 44860 127348 44872
rect 34572 44832 127348 44860
rect 34572 44820 34578 44832
rect 127342 44820 127348 44832
rect 127400 44820 127406 44872
rect 138474 44820 138480 44872
rect 138532 44860 138538 44872
rect 147030 44860 147036 44872
rect 138532 44832 147036 44860
rect 138532 44820 138538 44832
rect 147030 44820 147036 44832
rect 147088 44820 147094 44872
rect 171594 43392 171600 43444
rect 171652 43432 171658 43444
rect 411254 43432 411260 43444
rect 171652 43404 411260 43432
rect 171652 43392 171658 43404
rect 411254 43392 411260 43404
rect 411312 43392 411318 43444
rect 19334 42032 19340 42084
rect 19392 42072 19398 42084
rect 125134 42072 125140 42084
rect 19392 42044 125140 42072
rect 19392 42032 19398 42044
rect 125134 42032 125140 42044
rect 125192 42032 125198 42084
rect 162486 42032 162492 42084
rect 162544 42072 162550 42084
rect 390646 42072 390652 42084
rect 162544 42044 390652 42072
rect 162544 42032 162550 42044
rect 390646 42032 390652 42044
rect 390704 42032 390710 42084
rect 172422 40672 172428 40724
rect 172480 40712 172486 40724
rect 418154 40712 418160 40724
rect 172480 40684 418160 40712
rect 172480 40672 172486 40684
rect 418154 40672 418160 40684
rect 418212 40672 418218 40724
rect 120074 40264 120080 40316
rect 120132 40304 120138 40316
rect 123478 40304 123484 40316
rect 120132 40276 123484 40304
rect 120132 40264 120138 40276
rect 123478 40264 123484 40276
rect 123536 40264 123542 40316
rect 172330 39312 172336 39364
rect 172388 39352 172394 39364
rect 404354 39352 404360 39364
rect 172388 39324 404360 39352
rect 172388 39312 172394 39324
rect 404354 39312 404360 39324
rect 404412 39312 404418 39364
rect 172146 37884 172152 37936
rect 172204 37924 172210 37936
rect 397454 37924 397460 37936
rect 172204 37896 397460 37924
rect 172204 37884 172210 37896
rect 397454 37884 397460 37896
rect 397512 37884 397518 37936
rect 88334 36524 88340 36576
rect 88392 36564 88398 36576
rect 125042 36564 125048 36576
rect 88392 36536 125048 36564
rect 88392 36524 88398 36536
rect 125042 36524 125048 36536
rect 125100 36524 125106 36576
rect 145374 35572 145380 35624
rect 145432 35612 145438 35624
rect 259454 35612 259460 35624
rect 145432 35584 259460 35612
rect 145432 35572 145438 35584
rect 259454 35572 259460 35584
rect 259512 35572 259518 35624
rect 146938 35504 146944 35556
rect 146996 35544 147002 35556
rect 276014 35544 276020 35556
rect 146996 35516 276020 35544
rect 146996 35504 147002 35516
rect 276014 35504 276020 35516
rect 276072 35504 276078 35556
rect 148134 35436 148140 35488
rect 148192 35476 148198 35488
rect 287054 35476 287060 35488
rect 148192 35448 287060 35476
rect 148192 35436 148198 35448
rect 287054 35436 287060 35448
rect 287112 35436 287118 35488
rect 148042 35368 148048 35420
rect 148100 35408 148106 35420
rect 293954 35408 293960 35420
rect 148100 35380 293960 35408
rect 148100 35368 148106 35380
rect 293954 35368 293960 35380
rect 294012 35368 294018 35420
rect 149422 35300 149428 35352
rect 149480 35340 149486 35352
rect 304994 35340 305000 35352
rect 149480 35312 305000 35340
rect 149480 35300 149486 35312
rect 304994 35300 305000 35312
rect 305052 35300 305058 35352
rect 149514 35232 149520 35284
rect 149572 35272 149578 35284
rect 307754 35272 307760 35284
rect 149572 35244 307760 35272
rect 149572 35232 149578 35244
rect 307754 35232 307760 35244
rect 307812 35232 307818 35284
rect 159726 35164 159732 35216
rect 159784 35204 159790 35216
rect 382366 35204 382372 35216
rect 159784 35176 382372 35204
rect 159784 35164 159790 35176
rect 382366 35164 382372 35176
rect 382424 35164 382430 35216
rect 139670 34076 139676 34128
rect 139728 34116 139734 34128
rect 187694 34116 187700 34128
rect 139728 34088 187700 34116
rect 139728 34076 139734 34088
rect 187694 34076 187700 34088
rect 187752 34076 187758 34128
rect 141050 34008 141056 34060
rect 141108 34048 141114 34060
rect 198734 34048 198740 34060
rect 141108 34020 198740 34048
rect 141108 34008 141114 34020
rect 198734 34008 198740 34020
rect 198792 34008 198798 34060
rect 141234 33940 141240 33992
rect 141292 33980 141298 33992
rect 201494 33980 201500 33992
rect 141292 33952 201500 33980
rect 141292 33940 141298 33952
rect 201494 33940 201500 33952
rect 201552 33940 201558 33992
rect 141142 33872 141148 33924
rect 141200 33912 141206 33924
rect 205634 33912 205640 33924
rect 141200 33884 205640 33912
rect 141200 33872 141206 33884
rect 205634 33872 205640 33884
rect 205692 33872 205698 33924
rect 144086 33804 144092 33856
rect 144144 33844 144150 33856
rect 234706 33844 234712 33856
rect 144144 33816 234712 33844
rect 144144 33804 144150 33816
rect 234706 33804 234712 33816
rect 234764 33804 234770 33856
rect 146846 33736 146852 33788
rect 146904 33776 146910 33788
rect 269114 33776 269120 33788
rect 146904 33748 269120 33776
rect 146904 33736 146910 33748
rect 269114 33736 269120 33748
rect 269172 33736 269178 33788
rect 171686 33056 171692 33108
rect 171744 33096 171750 33108
rect 580166 33096 580172 33108
rect 171744 33068 580172 33096
rect 171744 33056 171750 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 3418 32988 3424 33040
rect 3476 33028 3482 33040
rect 181254 33028 181260 33040
rect 3476 33000 181260 33028
rect 3476 32988 3482 33000
rect 181254 32988 181260 33000
rect 181312 32988 181318 33040
rect 156414 32716 156420 32768
rect 156472 32756 156478 32768
rect 391934 32756 391940 32768
rect 156472 32728 391940 32756
rect 156472 32716 156478 32728
rect 391934 32716 391940 32728
rect 391992 32716 391998 32768
rect 160002 32648 160008 32700
rect 160060 32688 160066 32700
rect 434714 32688 434720 32700
rect 160060 32660 434720 32688
rect 160060 32648 160066 32660
rect 434714 32648 434720 32660
rect 434772 32648 434778 32700
rect 161934 32580 161940 32632
rect 161992 32620 161998 32632
rect 463694 32620 463700 32632
rect 161992 32592 463700 32620
rect 161992 32580 161998 32592
rect 463694 32580 463700 32592
rect 463752 32580 463758 32632
rect 163406 32512 163412 32564
rect 163464 32552 163470 32564
rect 481726 32552 481732 32564
rect 163464 32524 481732 32552
rect 163464 32512 163470 32524
rect 481726 32512 481732 32524
rect 481784 32512 481790 32564
rect 167546 32444 167552 32496
rect 167604 32484 167610 32496
rect 539686 32484 539692 32496
rect 167604 32456 539692 32484
rect 167604 32444 167610 32456
rect 539686 32444 539692 32456
rect 539744 32444 539750 32496
rect 170122 32376 170128 32428
rect 170180 32416 170186 32428
rect 574094 32416 574100 32428
rect 170180 32388 574100 32416
rect 170180 32376 170186 32388
rect 574094 32376 574100 32388
rect 574152 32376 574158 32428
rect 143994 31424 144000 31476
rect 144052 31464 144058 31476
rect 242894 31464 242900 31476
rect 144052 31436 242900 31464
rect 144052 31424 144058 31436
rect 242894 31424 242900 31436
rect 242952 31424 242958 31476
rect 146754 31356 146760 31408
rect 146812 31396 146818 31408
rect 267826 31396 267832 31408
rect 146812 31368 267832 31396
rect 146812 31356 146818 31368
rect 267826 31356 267832 31368
rect 267884 31356 267890 31408
rect 147950 31288 147956 31340
rect 148008 31328 148014 31340
rect 289814 31328 289820 31340
rect 148008 31300 289820 31328
rect 148008 31288 148014 31300
rect 289814 31288 289820 31300
rect 289872 31288 289878 31340
rect 154114 31220 154120 31272
rect 154172 31260 154178 31272
rect 332594 31260 332600 31272
rect 154172 31232 332600 31260
rect 154172 31220 154178 31232
rect 332594 31220 332600 31232
rect 332652 31220 332658 31272
rect 153562 31152 153568 31204
rect 153620 31192 153626 31204
rect 357526 31192 357532 31204
rect 153620 31164 357532 31192
rect 153620 31152 153626 31164
rect 357526 31152 357532 31164
rect 357584 31152 357590 31204
rect 156966 31084 156972 31136
rect 157024 31124 157030 31136
rect 389174 31124 389180 31136
rect 157024 31096 389180 31124
rect 157024 31084 157030 31096
rect 389174 31084 389180 31096
rect 389232 31084 389238 31136
rect 166258 31016 166264 31068
rect 166316 31056 166322 31068
rect 524414 31056 524420 31068
rect 166316 31028 524420 31056
rect 166316 31016 166322 31028
rect 524414 31016 524420 31028
rect 524472 31016 524478 31068
rect 140958 30064 140964 30116
rect 141016 30104 141022 30116
rect 204254 30104 204260 30116
rect 141016 30076 204260 30104
rect 141016 30064 141022 30076
rect 204254 30064 204260 30076
rect 204312 30064 204318 30116
rect 140866 29996 140872 30048
rect 140924 30036 140930 30048
rect 208394 30036 208400 30048
rect 140924 30008 208400 30036
rect 140924 29996 140930 30008
rect 208394 29996 208400 30008
rect 208452 29996 208458 30048
rect 143902 29928 143908 29980
rect 143960 29968 143966 29980
rect 233234 29968 233240 29980
rect 143960 29940 233240 29968
rect 143960 29928 143966 29940
rect 233234 29928 233240 29940
rect 233292 29928 233298 29980
rect 143810 29860 143816 29912
rect 143868 29900 143874 29912
rect 235994 29900 236000 29912
rect 143868 29872 236000 29900
rect 143868 29860 143874 29872
rect 235994 29860 236000 29872
rect 236052 29860 236058 29912
rect 145190 29792 145196 29844
rect 145248 29832 145254 29844
rect 253934 29832 253940 29844
rect 145248 29804 253940 29832
rect 145248 29792 145254 29804
rect 253934 29792 253940 29804
rect 253992 29792 253998 29844
rect 145282 29724 145288 29776
rect 145340 29764 145346 29776
rect 258074 29764 258080 29776
rect 145340 29736 258080 29764
rect 145340 29724 145346 29736
rect 258074 29724 258080 29736
rect 258132 29724 258138 29776
rect 166166 29656 166172 29708
rect 166224 29696 166230 29708
rect 521654 29696 521660 29708
rect 166224 29668 521660 29696
rect 166224 29656 166230 29668
rect 521654 29656 521660 29668
rect 521712 29656 521718 29708
rect 167454 29588 167460 29640
rect 167512 29628 167518 29640
rect 542354 29628 542360 29640
rect 167512 29600 542360 29628
rect 167512 29588 167518 29600
rect 542354 29588 542360 29600
rect 542412 29588 542418 29640
rect 148686 28500 148692 28552
rect 148744 28540 148750 28552
rect 190454 28540 190460 28552
rect 148744 28512 190460 28540
rect 148744 28500 148750 28512
rect 190454 28500 190460 28512
rect 190512 28500 190518 28552
rect 139578 28432 139584 28484
rect 139636 28472 139642 28484
rect 186314 28472 186320 28484
rect 139636 28444 186320 28472
rect 139636 28432 139642 28444
rect 186314 28432 186320 28444
rect 186372 28432 186378 28484
rect 140774 28364 140780 28416
rect 140832 28404 140838 28416
rect 201586 28404 201592 28416
rect 140832 28376 201592 28404
rect 140832 28364 140838 28376
rect 201586 28364 201592 28376
rect 201644 28364 201650 28416
rect 146662 28296 146668 28348
rect 146720 28336 146726 28348
rect 271874 28336 271880 28348
rect 146720 28308 271880 28336
rect 146720 28296 146726 28308
rect 271874 28296 271880 28308
rect 271932 28296 271938 28348
rect 147858 28228 147864 28280
rect 147916 28268 147922 28280
rect 285674 28268 285680 28280
rect 147916 28240 285680 28268
rect 147916 28228 147922 28240
rect 285674 28228 285680 28240
rect 285732 28228 285738 28280
rect 322198 28228 322204 28280
rect 322256 28268 322262 28280
rect 580994 28268 581000 28280
rect 322256 28240 581000 28268
rect 322256 28228 322262 28240
rect 580994 28228 581000 28240
rect 581052 28228 581058 28280
rect 140498 27276 140504 27328
rect 140556 27316 140562 27328
rect 176746 27316 176752 27328
rect 140556 27288 176752 27316
rect 140556 27276 140562 27288
rect 176746 27276 176752 27288
rect 176804 27276 176810 27328
rect 139486 27208 139492 27260
rect 139544 27248 139550 27260
rect 179414 27248 179420 27260
rect 139544 27220 179420 27248
rect 139544 27208 139550 27220
rect 179414 27208 179420 27220
rect 179472 27208 179478 27260
rect 139394 27140 139400 27192
rect 139452 27180 139458 27192
rect 183554 27180 183560 27192
rect 139452 27152 183560 27180
rect 139452 27140 139458 27152
rect 183554 27140 183560 27152
rect 183612 27140 183618 27192
rect 146570 27072 146576 27124
rect 146628 27112 146634 27124
rect 276106 27112 276112 27124
rect 146628 27084 276112 27112
rect 146628 27072 146634 27084
rect 276106 27072 276112 27084
rect 276164 27072 276170 27124
rect 149330 27004 149336 27056
rect 149388 27044 149394 27056
rect 310514 27044 310520 27056
rect 149388 27016 310520 27044
rect 149388 27004 149394 27016
rect 310514 27004 310520 27016
rect 310572 27004 310578 27056
rect 152274 26936 152280 26988
rect 152332 26976 152338 26988
rect 339494 26976 339500 26988
rect 152332 26948 339500 26976
rect 152332 26936 152338 26948
rect 339494 26936 339500 26948
rect 339552 26936 339558 26988
rect 164694 26868 164700 26920
rect 164752 26908 164758 26920
rect 506474 26908 506480 26920
rect 164752 26880 506480 26908
rect 164752 26868 164758 26880
rect 506474 26868 506480 26880
rect 506532 26868 506538 26920
rect 142522 25984 142528 26036
rect 142580 26024 142586 26036
rect 222194 26024 222200 26036
rect 142580 25996 222200 26024
rect 142580 25984 142586 25996
rect 222194 25984 222200 25996
rect 222252 25984 222258 26036
rect 146478 25916 146484 25968
rect 146536 25956 146542 25968
rect 278774 25956 278780 25968
rect 146536 25928 278780 25956
rect 146536 25916 146542 25928
rect 278774 25916 278780 25928
rect 278832 25916 278838 25968
rect 149238 25848 149244 25900
rect 149296 25888 149302 25900
rect 307846 25888 307852 25900
rect 149296 25860 307852 25888
rect 149296 25848 149302 25860
rect 307846 25848 307852 25860
rect 307904 25848 307910 25900
rect 152182 25780 152188 25832
rect 152240 25820 152246 25832
rect 346394 25820 346400 25832
rect 152240 25792 346400 25820
rect 152240 25780 152246 25792
rect 346394 25780 346400 25792
rect 346452 25780 346458 25832
rect 166074 25712 166080 25764
rect 166132 25752 166138 25764
rect 517514 25752 517520 25764
rect 166132 25724 517520 25752
rect 166132 25712 166138 25724
rect 517514 25712 517520 25724
rect 517572 25712 517578 25764
rect 170674 25644 170680 25696
rect 170732 25684 170738 25696
rect 558914 25684 558920 25696
rect 170732 25656 558920 25684
rect 170732 25644 170738 25656
rect 558914 25644 558920 25656
rect 558972 25644 558978 25696
rect 168834 25576 168840 25628
rect 168892 25616 168898 25628
rect 563054 25616 563060 25628
rect 168892 25588 563060 25616
rect 168892 25576 168898 25588
rect 563054 25576 563060 25588
rect 563112 25576 563118 25628
rect 170030 25508 170036 25560
rect 170088 25548 170094 25560
rect 572714 25548 572720 25560
rect 170088 25520 572720 25548
rect 170088 25508 170094 25520
rect 572714 25508 572720 25520
rect 572772 25508 572778 25560
rect 142338 24556 142344 24608
rect 142396 24596 142402 24608
rect 215294 24596 215300 24608
rect 142396 24568 215300 24596
rect 142396 24556 142402 24568
rect 215294 24556 215300 24568
rect 215352 24556 215358 24608
rect 142430 24488 142436 24540
rect 142488 24528 142494 24540
rect 218146 24528 218152 24540
rect 142488 24500 218152 24528
rect 142488 24488 142494 24500
rect 218146 24488 218152 24500
rect 218204 24488 218210 24540
rect 147766 24420 147772 24472
rect 147824 24460 147830 24472
rect 292666 24460 292672 24472
rect 147824 24432 292672 24460
rect 147824 24420 147830 24432
rect 292666 24420 292672 24432
rect 292724 24420 292730 24472
rect 155034 24352 155040 24404
rect 155092 24392 155098 24404
rect 374086 24392 374092 24404
rect 155092 24364 374092 24392
rect 155092 24352 155098 24364
rect 374086 24352 374092 24364
rect 374144 24352 374150 24404
rect 167178 24284 167184 24336
rect 167236 24324 167242 24336
rect 467098 24324 467104 24336
rect 167236 24296 467104 24324
rect 167236 24284 167242 24296
rect 467098 24284 467104 24296
rect 467156 24284 467162 24336
rect 167270 24216 167276 24268
rect 167328 24256 167334 24268
rect 535454 24256 535460 24268
rect 167328 24228 535460 24256
rect 167328 24216 167334 24228
rect 535454 24216 535460 24228
rect 535512 24216 535518 24268
rect 167362 24148 167368 24200
rect 167420 24188 167426 24200
rect 538214 24188 538220 24200
rect 167420 24160 538220 24188
rect 167420 24148 167426 24160
rect 538214 24148 538220 24160
rect 538272 24148 538278 24200
rect 168742 24080 168748 24132
rect 168800 24120 168806 24132
rect 552014 24120 552020 24132
rect 168800 24092 552020 24120
rect 168800 24080 168806 24092
rect 552014 24080 552020 24092
rect 552072 24080 552078 24132
rect 149146 23332 149152 23384
rect 149204 23372 149210 23384
rect 303614 23372 303620 23384
rect 149204 23344 303620 23372
rect 149204 23332 149210 23344
rect 303614 23332 303620 23344
rect 303672 23332 303678 23384
rect 3418 23264 3424 23316
rect 3476 23304 3482 23316
rect 173986 23304 173992 23316
rect 3476 23276 173992 23304
rect 3476 23264 3482 23276
rect 173986 23264 173992 23276
rect 174044 23264 174050 23316
rect 153470 23196 153476 23248
rect 153528 23236 153534 23248
rect 360194 23236 360200 23248
rect 153528 23208 360200 23236
rect 153528 23196 153534 23208
rect 360194 23196 360200 23208
rect 360252 23196 360258 23248
rect 154942 23128 154948 23180
rect 155000 23168 155006 23180
rect 379514 23168 379520 23180
rect 155000 23140 379520 23168
rect 155000 23128 155006 23140
rect 379514 23128 379520 23140
rect 379572 23128 379578 23180
rect 164602 23060 164608 23112
rect 164660 23100 164666 23112
rect 498286 23100 498292 23112
rect 164660 23072 498292 23100
rect 164660 23060 164666 23072
rect 498286 23060 498292 23072
rect 498344 23060 498350 23112
rect 164510 22992 164516 23044
rect 164568 23032 164574 23044
rect 509234 23032 509240 23044
rect 164568 23004 509240 23032
rect 164568 22992 164574 23004
rect 509234 22992 509240 23004
rect 509292 22992 509298 23044
rect 165890 22924 165896 22976
rect 165948 22964 165954 22976
rect 516134 22964 516140 22976
rect 165948 22936 516140 22964
rect 165948 22924 165954 22936
rect 516134 22924 516140 22936
rect 516192 22924 516198 22976
rect 165982 22856 165988 22908
rect 166040 22896 166046 22908
rect 520274 22896 520280 22908
rect 166040 22868 520280 22896
rect 166040 22856 166046 22868
rect 520274 22856 520280 22868
rect 520332 22856 520338 22908
rect 74534 22788 74540 22840
rect 74592 22828 74598 22840
rect 129182 22828 129188 22840
rect 74592 22800 129188 22828
rect 74592 22788 74598 22800
rect 129182 22788 129188 22800
rect 129240 22788 129246 22840
rect 168650 22788 168656 22840
rect 168708 22828 168714 22840
rect 556154 22828 556160 22840
rect 168708 22800 556160 22828
rect 168708 22788 168714 22800
rect 556154 22788 556160 22800
rect 556212 22788 556218 22840
rect 118418 22720 118424 22772
rect 118476 22760 118482 22772
rect 580166 22760 580172 22772
rect 118476 22732 580172 22760
rect 118476 22720 118482 22732
rect 580166 22720 580172 22732
rect 580224 22720 580230 22772
rect 152090 21632 152096 21684
rect 152148 21672 152154 21684
rect 343634 21672 343640 21684
rect 152148 21644 343640 21672
rect 152148 21632 152154 21644
rect 343634 21632 343640 21644
rect 343692 21632 343698 21684
rect 160646 21564 160652 21616
rect 160704 21604 160710 21616
rect 447134 21604 447140 21616
rect 160704 21576 447140 21604
rect 160704 21564 160710 21576
rect 447134 21564 447140 21576
rect 447192 21564 447198 21616
rect 161842 21496 161848 21548
rect 161900 21536 161906 21548
rect 473354 21536 473360 21548
rect 161900 21508 473360 21536
rect 161900 21496 161906 21508
rect 473354 21496 473360 21508
rect 473412 21496 473418 21548
rect 163314 21428 163320 21480
rect 163372 21468 163378 21480
rect 484394 21468 484400 21480
rect 163372 21440 484400 21468
rect 163372 21428 163378 21440
rect 484394 21428 484400 21440
rect 484452 21428 484458 21480
rect 124306 21360 124312 21412
rect 124364 21400 124370 21412
rect 134334 21400 134340 21412
rect 124364 21372 134340 21400
rect 124364 21360 124370 21372
rect 134334 21360 134340 21372
rect 134392 21360 134398 21412
rect 164418 21360 164424 21412
rect 164476 21400 164482 21412
rect 506566 21400 506572 21412
rect 164476 21372 506572 21400
rect 164476 21360 164482 21372
rect 506566 21360 506572 21372
rect 506624 21360 506630 21412
rect 145098 20340 145104 20392
rect 145156 20380 145162 20392
rect 255314 20380 255320 20392
rect 145156 20352 255320 20380
rect 145156 20340 145162 20352
rect 255314 20340 255320 20352
rect 255372 20340 255378 20392
rect 145006 20272 145012 20324
rect 145064 20312 145070 20324
rect 262214 20312 262220 20324
rect 145064 20284 262220 20312
rect 145064 20272 145070 20284
rect 262214 20272 262220 20284
rect 262272 20272 262278 20324
rect 146386 20204 146392 20256
rect 146444 20244 146450 20256
rect 273254 20244 273260 20256
rect 146444 20216 273260 20244
rect 146444 20204 146450 20216
rect 273254 20204 273260 20216
rect 273312 20204 273318 20256
rect 247678 20136 247684 20188
rect 247736 20176 247742 20188
rect 456794 20176 456800 20188
rect 247736 20148 456800 20176
rect 247736 20136 247742 20148
rect 456794 20136 456800 20148
rect 456852 20136 456858 20188
rect 138382 20068 138388 20120
rect 138440 20108 138446 20120
rect 162854 20108 162860 20120
rect 138440 20080 162860 20108
rect 138440 20068 138446 20080
rect 162854 20068 162860 20080
rect 162912 20068 162918 20120
rect 253198 20068 253204 20120
rect 253256 20108 253262 20120
rect 465074 20108 465080 20120
rect 253256 20080 465080 20108
rect 253256 20068 253262 20080
rect 465074 20068 465080 20080
rect 465132 20068 465138 20120
rect 85574 20000 85580 20052
rect 85632 20040 85638 20052
rect 131666 20040 131672 20052
rect 85632 20012 131672 20040
rect 85632 20000 85638 20012
rect 131666 20000 131672 20012
rect 131724 20000 131730 20052
rect 160554 20000 160560 20052
rect 160612 20040 160618 20052
rect 455414 20040 455420 20052
rect 160612 20012 455420 20040
rect 160612 20000 160618 20012
rect 455414 20000 455420 20012
rect 455472 20000 455478 20052
rect 45554 19932 45560 19984
rect 45612 19972 45618 19984
rect 120810 19972 120816 19984
rect 45612 19944 120816 19972
rect 45612 19932 45618 19944
rect 120810 19932 120816 19944
rect 120868 19932 120874 19984
rect 161750 19932 161756 19984
rect 161808 19972 161814 19984
rect 465166 19972 465172 19984
rect 161808 19944 465172 19972
rect 161808 19932 161814 19944
rect 465166 19932 465172 19944
rect 465224 19932 465230 19984
rect 160462 18844 160468 18896
rect 160520 18884 160526 18896
rect 448514 18884 448520 18896
rect 160520 18856 448520 18884
rect 160520 18844 160526 18856
rect 448514 18844 448520 18856
rect 448572 18844 448578 18896
rect 160370 18776 160376 18828
rect 160428 18816 160434 18828
rect 451274 18816 451280 18828
rect 160428 18788 451280 18816
rect 160428 18776 160434 18788
rect 451274 18776 451280 18788
rect 451332 18776 451338 18828
rect 117314 18708 117320 18760
rect 117372 18748 117378 18760
rect 134242 18748 134248 18760
rect 117372 18720 134248 18748
rect 117372 18708 117378 18720
rect 134242 18708 134248 18720
rect 134300 18708 134306 18760
rect 168466 18708 168472 18760
rect 168524 18748 168530 18760
rect 553394 18748 553400 18760
rect 168524 18720 553400 18748
rect 168524 18708 168530 18720
rect 553394 18708 553400 18720
rect 553452 18708 553458 18760
rect 31754 18640 31760 18692
rect 31812 18680 31818 18692
rect 122282 18680 122288 18692
rect 31812 18652 122288 18680
rect 31812 18640 31818 18652
rect 122282 18640 122288 18652
rect 122340 18640 122346 18692
rect 168374 18640 168380 18692
rect 168432 18680 168438 18692
rect 556246 18680 556252 18692
rect 168432 18652 556252 18680
rect 168432 18640 168438 18652
rect 556246 18640 556252 18652
rect 556304 18640 556310 18692
rect 4154 18572 4160 18624
rect 4212 18612 4218 18624
rect 126238 18612 126244 18624
rect 4212 18584 126244 18612
rect 4212 18572 4218 18584
rect 126238 18572 126244 18584
rect 126296 18572 126302 18624
rect 168558 18572 168564 18624
rect 168616 18612 168622 18624
rect 560294 18612 560300 18624
rect 168616 18584 560300 18612
rect 168616 18572 168622 18584
rect 560294 18572 560300 18584
rect 560352 18572 560358 18624
rect 157794 17552 157800 17604
rect 157852 17592 157858 17604
rect 415394 17592 415400 17604
rect 157852 17564 415400 17592
rect 157852 17552 157858 17564
rect 415394 17552 415400 17564
rect 415452 17552 415458 17604
rect 157702 17484 157708 17536
rect 157760 17524 157766 17536
rect 419534 17524 419540 17536
rect 157760 17496 419540 17524
rect 157760 17484 157766 17496
rect 419534 17484 419540 17496
rect 419592 17484 419598 17536
rect 171962 17416 171968 17468
rect 172020 17456 172026 17468
rect 440234 17456 440240 17468
rect 172020 17428 440240 17456
rect 172020 17416 172026 17428
rect 440234 17416 440240 17428
rect 440292 17416 440298 17468
rect 160278 17348 160284 17400
rect 160336 17388 160342 17400
rect 448606 17388 448612 17400
rect 160336 17360 448612 17388
rect 160336 17348 160342 17360
rect 448606 17348 448612 17360
rect 448664 17348 448670 17400
rect 163222 17280 163228 17332
rect 163280 17320 163286 17332
rect 492674 17320 492680 17332
rect 163280 17292 492680 17320
rect 163280 17280 163286 17292
rect 492674 17280 492680 17292
rect 492732 17280 492738 17332
rect 167086 17212 167092 17264
rect 167144 17252 167150 17264
rect 545114 17252 545120 17264
rect 167144 17224 545120 17252
rect 167144 17212 167150 17224
rect 545114 17212 545120 17224
rect 545172 17212 545178 17264
rect 154850 16124 154856 16176
rect 154908 16164 154914 16176
rect 378410 16164 378416 16176
rect 154908 16136 378416 16164
rect 154908 16124 154914 16136
rect 378410 16124 378416 16136
rect 378468 16124 378474 16176
rect 156230 16056 156236 16108
rect 156288 16096 156294 16108
rect 395338 16096 395344 16108
rect 156288 16068 395344 16096
rect 156288 16056 156294 16068
rect 395338 16056 395344 16068
rect 395396 16056 395402 16108
rect 156322 15988 156328 16040
rect 156380 16028 156386 16040
rect 398834 16028 398840 16040
rect 156380 16000 398840 16028
rect 156380 15988 156386 16000
rect 398834 15988 398840 16000
rect 398892 15988 398898 16040
rect 174538 15920 174544 15972
rect 174596 15960 174602 15972
rect 425698 15960 425704 15972
rect 174596 15932 425704 15960
rect 174596 15920 174602 15932
rect 425698 15920 425704 15932
rect 425756 15920 425762 15972
rect 14274 15852 14280 15904
rect 14332 15892 14338 15904
rect 124950 15892 124956 15904
rect 14332 15864 124956 15892
rect 14332 15852 14338 15864
rect 124950 15852 124956 15864
rect 125008 15852 125014 15904
rect 166994 15852 167000 15904
rect 167052 15892 167058 15904
rect 541986 15892 541992 15904
rect 167052 15864 541992 15892
rect 167052 15852 167058 15864
rect 541986 15852 541992 15864
rect 542044 15852 542050 15904
rect 143718 14764 143724 14816
rect 143776 14804 143782 14816
rect 241698 14804 241704 14816
rect 143776 14776 241704 14804
rect 143776 14764 143782 14776
rect 241698 14764 241704 14776
rect 241756 14764 241762 14816
rect 154666 14696 154672 14748
rect 154724 14736 154730 14748
rect 381170 14736 381176 14748
rect 154724 14708 381176 14736
rect 154724 14696 154730 14708
rect 381170 14696 381176 14708
rect 381228 14696 381234 14748
rect 154758 14628 154764 14680
rect 154816 14668 154822 14680
rect 384298 14668 384304 14680
rect 154816 14640 384304 14668
rect 154816 14628 154822 14640
rect 384298 14628 384304 14640
rect 384356 14628 384362 14680
rect 154574 14560 154580 14612
rect 154632 14600 154638 14612
rect 385954 14600 385960 14612
rect 154632 14572 385960 14600
rect 154632 14560 154638 14572
rect 385954 14560 385960 14572
rect 386012 14560 386018 14612
rect 114002 14492 114008 14544
rect 114060 14532 114066 14544
rect 134150 14532 134156 14544
rect 114060 14504 134156 14532
rect 114060 14492 114066 14504
rect 134150 14492 134156 14504
rect 134208 14492 134214 14544
rect 158898 14492 158904 14544
rect 158956 14532 158962 14544
rect 436738 14532 436744 14544
rect 158956 14504 436744 14532
rect 158956 14492 158962 14504
rect 436738 14492 436744 14504
rect 436796 14492 436802 14544
rect 39114 14424 39120 14476
rect 39172 14464 39178 14476
rect 120718 14464 120724 14476
rect 39172 14436 120724 14464
rect 39172 14424 39178 14436
rect 120718 14424 120724 14436
rect 120776 14424 120782 14476
rect 164326 14424 164332 14476
rect 164384 14464 164390 14476
rect 502978 14464 502984 14476
rect 164384 14436 502984 14464
rect 164384 14424 164390 14436
rect 502978 14424 502984 14436
rect 503036 14424 503042 14476
rect 151906 13404 151912 13456
rect 151964 13444 151970 13456
rect 345290 13444 345296 13456
rect 151964 13416 345296 13444
rect 151964 13404 151970 13416
rect 345290 13404 345296 13416
rect 345348 13404 345354 13456
rect 151998 13336 152004 13388
rect 152056 13376 152062 13388
rect 349154 13376 349160 13388
rect 152056 13348 349160 13376
rect 152056 13336 152062 13348
rect 349154 13336 349160 13348
rect 349212 13336 349218 13388
rect 153378 13268 153384 13320
rect 153436 13308 153442 13320
rect 365714 13308 365720 13320
rect 153436 13280 365720 13308
rect 153436 13268 153442 13280
rect 365714 13268 365720 13280
rect 365772 13268 365778 13320
rect 157610 13200 157616 13252
rect 157668 13240 157674 13252
rect 417418 13240 417424 13252
rect 157668 13212 417424 13240
rect 157668 13200 157674 13212
rect 417418 13200 417424 13212
rect 417476 13200 417482 13252
rect 158806 13132 158812 13184
rect 158864 13172 158870 13184
rect 429194 13172 429200 13184
rect 158864 13144 429200 13172
rect 158864 13132 158870 13144
rect 429194 13132 429200 13144
rect 429252 13132 429258 13184
rect 160186 13064 160192 13116
rect 160244 13104 160250 13116
rect 453298 13104 453304 13116
rect 160244 13076 453304 13104
rect 160244 13064 160250 13076
rect 453298 13064 453304 13076
rect 453356 13064 453362 13116
rect 143626 11976 143632 12028
rect 143684 12016 143690 12028
rect 237650 12016 237656 12028
rect 143684 11988 237656 12016
rect 143684 11976 143690 11988
rect 237650 11976 237656 11988
rect 237708 11976 237714 12028
rect 150342 11908 150348 11960
rect 150400 11948 150406 11960
rect 313826 11948 313832 11960
rect 150400 11920 313832 11948
rect 150400 11908 150406 11920
rect 313826 11908 313832 11920
rect 313884 11908 313890 11960
rect 157518 11840 157524 11892
rect 157576 11880 157582 11892
rect 414290 11880 414296 11892
rect 157576 11852 414296 11880
rect 157576 11840 157582 11852
rect 414290 11840 414296 11852
rect 414348 11840 414354 11892
rect 157426 11772 157432 11824
rect 157484 11812 157490 11824
rect 415486 11812 415492 11824
rect 157484 11784 415492 11812
rect 157484 11772 157490 11784
rect 415486 11772 415492 11784
rect 415544 11772 415550 11824
rect 165798 11704 165804 11756
rect 165856 11744 165862 11756
rect 523770 11744 523776 11756
rect 165856 11716 523776 11744
rect 165856 11704 165862 11716
rect 523770 11704 523776 11716
rect 523828 11704 523834 11756
rect 176654 11636 176660 11688
rect 176712 11676 176718 11688
rect 177850 11676 177856 11688
rect 176712 11648 177856 11676
rect 176712 11636 176718 11648
rect 177850 11636 177856 11648
rect 177908 11636 177914 11688
rect 184934 11636 184940 11688
rect 184992 11676 184998 11688
rect 186130 11676 186136 11688
rect 184992 11648 186136 11676
rect 184992 11636 184998 11648
rect 186130 11636 186136 11648
rect 186188 11636 186194 11688
rect 201494 11636 201500 11688
rect 201552 11676 201558 11688
rect 202690 11676 202696 11688
rect 201552 11648 202696 11676
rect 201552 11636 201558 11648
rect 202690 11636 202696 11648
rect 202748 11636 202754 11688
rect 234614 11636 234620 11688
rect 234672 11676 234678 11688
rect 235810 11676 235816 11688
rect 234672 11648 235816 11676
rect 234672 11636 234678 11648
rect 235810 11636 235816 11648
rect 235868 11636 235874 11688
rect 106458 10616 106464 10668
rect 106516 10656 106522 10668
rect 133046 10656 133052 10668
rect 106516 10628 133052 10656
rect 106516 10616 106522 10628
rect 133046 10616 133052 10628
rect 133104 10616 133110 10668
rect 99834 10548 99840 10600
rect 99892 10588 99898 10600
rect 132954 10588 132960 10600
rect 99892 10560 132960 10588
rect 99892 10548 99898 10560
rect 132954 10548 132960 10560
rect 133012 10548 133018 10600
rect 147674 10548 147680 10600
rect 147732 10588 147738 10600
rect 295610 10588 295616 10600
rect 147732 10560 295616 10588
rect 147732 10548 147738 10560
rect 295610 10548 295616 10560
rect 295668 10548 295674 10600
rect 81618 10480 81624 10532
rect 81676 10520 81682 10532
rect 131574 10520 131580 10532
rect 81676 10492 131580 10520
rect 81676 10480 81682 10492
rect 131574 10480 131580 10492
rect 131632 10480 131638 10532
rect 153286 10480 153292 10532
rect 153344 10520 153350 10532
rect 364610 10520 364616 10532
rect 153344 10492 364616 10520
rect 153344 10480 153350 10492
rect 364610 10480 364616 10492
rect 364668 10480 364674 10532
rect 35986 10412 35992 10464
rect 36044 10452 36050 10464
rect 127250 10452 127256 10464
rect 36044 10424 127256 10452
rect 36044 10412 36050 10424
rect 127250 10412 127256 10424
rect 127308 10412 127314 10464
rect 156046 10412 156052 10464
rect 156104 10452 156110 10464
rect 394234 10452 394240 10464
rect 156104 10424 394240 10452
rect 156104 10412 156110 10424
rect 394234 10412 394240 10424
rect 394292 10412 394298 10464
rect 28442 10344 28448 10396
rect 28500 10384 28506 10396
rect 127158 10384 127164 10396
rect 28500 10356 127164 10384
rect 28500 10344 28506 10356
rect 127158 10344 127164 10356
rect 127216 10344 127222 10396
rect 156138 10344 156144 10396
rect 156196 10384 156202 10396
rect 398926 10384 398932 10396
rect 156196 10356 398932 10384
rect 156196 10344 156202 10356
rect 398926 10344 398932 10356
rect 398984 10344 398990 10396
rect 11146 10276 11152 10328
rect 11204 10316 11210 10328
rect 126146 10316 126152 10328
rect 11204 10288 126152 10316
rect 11204 10276 11210 10288
rect 126146 10276 126152 10288
rect 126204 10276 126210 10328
rect 163130 10276 163136 10328
rect 163188 10316 163194 10328
rect 486418 10316 486424 10328
rect 163188 10288 486424 10316
rect 163188 10276 163194 10288
rect 486418 10276 486424 10288
rect 486476 10276 486482 10328
rect 67910 9324 67916 9376
rect 67968 9364 67974 9376
rect 130194 9364 130200 9376
rect 67968 9336 130200 9364
rect 67968 9324 67974 9336
rect 130194 9324 130200 9336
rect 130252 9324 130258 9376
rect 64322 9256 64328 9308
rect 64380 9296 64386 9308
rect 126330 9296 126336 9308
rect 64380 9268 126336 9296
rect 64380 9256 64386 9268
rect 126330 9256 126336 9268
rect 126388 9256 126394 9308
rect 144914 9256 144920 9308
rect 144972 9296 144978 9308
rect 260650 9296 260656 9308
rect 144972 9268 260656 9296
rect 144972 9256 144978 9268
rect 260650 9256 260656 9268
rect 260708 9256 260714 9308
rect 63218 9188 63224 9240
rect 63276 9228 63282 9240
rect 130102 9228 130108 9240
rect 63276 9200 130108 9228
rect 63276 9188 63282 9200
rect 130102 9188 130108 9200
rect 130160 9188 130166 9240
rect 146294 9188 146300 9240
rect 146352 9228 146358 9240
rect 278314 9228 278320 9240
rect 146352 9200 278320 9228
rect 146352 9188 146358 9200
rect 278314 9188 278320 9200
rect 278372 9188 278378 9240
rect 60826 9120 60832 9172
rect 60884 9160 60890 9172
rect 129090 9160 129096 9172
rect 60884 9132 129096 9160
rect 60884 9120 60890 9132
rect 129090 9120 129096 9132
rect 129148 9120 129154 9172
rect 151814 9120 151820 9172
rect 151872 9160 151878 9172
rect 343358 9160 343364 9172
rect 151872 9132 343364 9160
rect 151872 9120 151878 9132
rect 343358 9120 343364 9132
rect 343416 9120 343422 9172
rect 53742 9052 53748 9104
rect 53800 9092 53806 9104
rect 128722 9092 128728 9104
rect 53800 9064 128728 9092
rect 53800 9052 53806 9064
rect 128722 9052 128728 9064
rect 128780 9052 128786 9104
rect 161658 9052 161664 9104
rect 161716 9092 161722 9104
rect 471054 9092 471060 9104
rect 161716 9064 471060 9092
rect 161716 9052 161722 9064
rect 471054 9052 471060 9064
rect 471112 9052 471118 9104
rect 50154 8984 50160 9036
rect 50212 9024 50218 9036
rect 127710 9024 127716 9036
rect 50212 8996 127716 9024
rect 50212 8984 50218 8996
rect 127710 8984 127716 8996
rect 127768 8984 127774 9036
rect 163038 8984 163044 9036
rect 163096 9024 163102 9036
rect 492306 9024 492312 9036
rect 163096 8996 492312 9024
rect 163096 8984 163102 8996
rect 492306 8984 492312 8996
rect 492364 8984 492370 9036
rect 566 8916 572 8968
rect 624 8956 630 8968
rect 124214 8956 124220 8968
rect 624 8928 124220 8956
rect 624 8916 630 8928
rect 124214 8916 124220 8928
rect 124272 8916 124278 8968
rect 169938 8916 169944 8968
rect 169996 8956 170002 8968
rect 571518 8956 571524 8968
rect 169996 8928 571524 8956
rect 169996 8916 170002 8928
rect 571518 8916 571524 8928
rect 571576 8916 571582 8968
rect 116394 7896 116400 7948
rect 116452 7936 116458 7948
rect 134058 7936 134064 7948
rect 116452 7908 134064 7936
rect 116452 7896 116458 7908
rect 134058 7896 134064 7908
rect 134116 7896 134122 7948
rect 142246 7896 142252 7948
rect 142304 7936 142310 7948
rect 225138 7936 225144 7948
rect 142304 7908 225144 7936
rect 142304 7896 142310 7908
rect 225138 7896 225144 7908
rect 225196 7896 225202 7948
rect 105722 7828 105728 7880
rect 105780 7868 105786 7880
rect 132770 7868 132776 7880
rect 105780 7840 132776 7868
rect 105780 7828 105786 7840
rect 132770 7828 132776 7840
rect 132828 7828 132834 7880
rect 143534 7828 143540 7880
rect 143592 7868 143598 7880
rect 242986 7868 242992 7880
rect 143592 7840 242992 7868
rect 143592 7828 143598 7840
rect 242986 7828 242992 7840
rect 243044 7828 243050 7880
rect 98638 7760 98644 7812
rect 98696 7800 98702 7812
rect 132862 7800 132868 7812
rect 98696 7772 132868 7800
rect 98696 7760 98702 7772
rect 132862 7760 132868 7772
rect 132920 7760 132926 7812
rect 155954 7760 155960 7812
rect 156012 7800 156018 7812
rect 401318 7800 401324 7812
rect 156012 7772 401324 7800
rect 156012 7760 156018 7772
rect 401318 7760 401324 7772
rect 401376 7760 401382 7812
rect 48958 7692 48964 7744
rect 49016 7732 49022 7744
rect 128538 7732 128544 7744
rect 49016 7704 128544 7732
rect 49016 7692 49022 7704
rect 128538 7692 128544 7704
rect 128596 7692 128602 7744
rect 160094 7692 160100 7744
rect 160152 7732 160158 7744
rect 446214 7732 446220 7744
rect 160152 7704 446220 7732
rect 160152 7692 160158 7704
rect 446214 7692 446220 7704
rect 446272 7692 446278 7744
rect 44266 7624 44272 7676
rect 44324 7664 44330 7676
rect 128630 7664 128636 7676
rect 44324 7636 128636 7664
rect 44324 7624 44330 7636
rect 128630 7624 128636 7636
rect 128688 7624 128694 7676
rect 161566 7624 161572 7676
rect 161624 7664 161630 7676
rect 469858 7664 469864 7676
rect 161624 7636 469864 7664
rect 161624 7624 161630 7636
rect 469858 7624 469864 7636
rect 469916 7624 469922 7676
rect 9950 7556 9956 7608
rect 10008 7596 10014 7608
rect 126054 7596 126060 7608
rect 10008 7568 126060 7596
rect 10008 7556 10014 7568
rect 126054 7556 126060 7568
rect 126112 7556 126118 7608
rect 164234 7556 164240 7608
rect 164292 7596 164298 7608
rect 504174 7596 504180 7608
rect 164292 7568 504180 7596
rect 164292 7556 164298 7568
rect 504174 7556 504180 7568
rect 504232 7556 504238 7608
rect 555418 6808 555424 6860
rect 555476 6848 555482 6860
rect 580166 6848 580172 6860
rect 555476 6820 580172 6848
rect 555476 6808 555482 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 150802 6740 150808 6792
rect 150860 6780 150866 6792
rect 323302 6780 323308 6792
rect 150860 6752 323308 6780
rect 150860 6740 150866 6752
rect 323302 6740 323308 6752
rect 323360 6740 323366 6792
rect 150986 6672 150992 6724
rect 151044 6712 151050 6724
rect 326798 6712 326804 6724
rect 151044 6684 326804 6712
rect 151044 6672 151050 6684
rect 326798 6672 326804 6684
rect 326856 6672 326862 6724
rect 115198 6604 115204 6656
rect 115256 6644 115262 6656
rect 134702 6644 134708 6656
rect 115256 6616 134708 6644
rect 115256 6604 115262 6616
rect 134702 6604 134708 6616
rect 134760 6604 134766 6656
rect 150894 6604 150900 6656
rect 150952 6644 150958 6656
rect 329190 6644 329196 6656
rect 150952 6616 329196 6644
rect 150952 6604 150958 6616
rect 329190 6604 329196 6616
rect 329248 6604 329254 6656
rect 104526 6536 104532 6588
rect 104584 6576 104590 6588
rect 132678 6576 132684 6588
rect 104584 6548 132684 6576
rect 104584 6536 104590 6548
rect 132678 6536 132684 6548
rect 132736 6536 132742 6588
rect 151078 6536 151084 6588
rect 151136 6576 151142 6588
rect 330386 6576 330392 6588
rect 151136 6548 330392 6576
rect 151136 6536 151142 6548
rect 330386 6536 330392 6548
rect 330444 6536 330450 6588
rect 84470 6468 84476 6520
rect 84528 6508 84534 6520
rect 131298 6508 131304 6520
rect 84528 6480 131304 6508
rect 84528 6468 84534 6480
rect 131298 6468 131304 6480
rect 131356 6468 131362 6520
rect 158530 6468 158536 6520
rect 158588 6508 158594 6520
rect 410794 6508 410800 6520
rect 158588 6480 410800 6508
rect 158588 6468 158594 6480
rect 410794 6468 410800 6480
rect 410852 6468 410858 6520
rect 80882 6400 80888 6452
rect 80940 6440 80946 6452
rect 131390 6440 131396 6452
rect 80940 6412 131396 6440
rect 80940 6400 80946 6412
rect 131390 6400 131396 6412
rect 131448 6400 131454 6452
rect 175918 6400 175924 6452
rect 175976 6440 175982 6452
rect 433242 6440 433248 6452
rect 175976 6412 433248 6440
rect 175976 6400 175982 6412
rect 433242 6400 433248 6412
rect 433300 6400 433306 6452
rect 77386 6332 77392 6384
rect 77444 6372 77450 6384
rect 131482 6372 131488 6384
rect 77444 6344 131488 6372
rect 77444 6332 77450 6344
rect 131482 6332 131488 6344
rect 131540 6332 131546 6384
rect 158714 6332 158720 6384
rect 158772 6372 158778 6384
rect 441522 6372 441528 6384
rect 158772 6344 441528 6372
rect 158772 6332 158778 6344
rect 441522 6332 441528 6344
rect 441580 6332 441586 6384
rect 25314 6264 25320 6316
rect 25372 6304 25378 6316
rect 57238 6304 57244 6316
rect 25372 6276 57244 6304
rect 25372 6264 25378 6276
rect 57238 6264 57244 6276
rect 57296 6264 57302 6316
rect 66714 6264 66720 6316
rect 66772 6304 66778 6316
rect 130010 6304 130016 6316
rect 66772 6276 130016 6304
rect 66772 6264 66778 6276
rect 130010 6264 130016 6276
rect 130068 6264 130074 6316
rect 161474 6264 161480 6316
rect 161532 6304 161538 6316
rect 467466 6304 467472 6316
rect 161532 6276 467472 6304
rect 161532 6264 161538 6276
rect 467466 6264 467472 6276
rect 467524 6264 467530 6316
rect 33594 6196 33600 6248
rect 33652 6236 33658 6248
rect 127526 6236 127532 6248
rect 33652 6208 127532 6236
rect 33652 6196 33658 6208
rect 127526 6196 127532 6208
rect 127584 6196 127590 6248
rect 140406 6196 140412 6248
rect 140464 6236 140470 6248
rect 156598 6236 156604 6248
rect 140464 6208 156604 6236
rect 140464 6196 140470 6208
rect 156598 6196 156604 6208
rect 156656 6196 156662 6248
rect 169754 6196 169760 6248
rect 169812 6236 169818 6248
rect 572714 6236 572720 6248
rect 169812 6208 572720 6236
rect 169812 6196 169818 6208
rect 572714 6196 572720 6208
rect 572772 6196 572778 6248
rect 18230 6128 18236 6180
rect 18288 6168 18294 6180
rect 125962 6168 125968 6180
rect 18288 6140 125968 6168
rect 18288 6128 18294 6140
rect 125962 6128 125968 6140
rect 126020 6128 126026 6180
rect 138290 6128 138296 6180
rect 138348 6168 138354 6180
rect 162486 6168 162492 6180
rect 138348 6140 162492 6168
rect 138348 6128 138354 6140
rect 162486 6128 162492 6140
rect 162544 6128 162550 6180
rect 169846 6128 169852 6180
rect 169904 6168 169910 6180
rect 576302 6168 576308 6180
rect 169904 6140 576308 6168
rect 169904 6128 169910 6140
rect 576302 6128 576308 6140
rect 576360 6128 576366 6180
rect 101030 5312 101036 5364
rect 101088 5352 101094 5364
rect 133138 5352 133144 5364
rect 101088 5324 133144 5352
rect 101088 5312 101094 5324
rect 133138 5312 133144 5324
rect 133196 5312 133202 5364
rect 97442 5244 97448 5296
rect 97500 5284 97506 5296
rect 132586 5284 132592 5296
rect 97500 5256 132592 5284
rect 97500 5244 97506 5256
rect 132586 5244 132592 5256
rect 132644 5244 132650 5296
rect 86862 5176 86868 5228
rect 86920 5216 86926 5228
rect 132402 5216 132408 5228
rect 86920 5188 132408 5216
rect 86920 5176 86926 5188
rect 132402 5176 132408 5188
rect 132460 5176 132466 5228
rect 138014 5176 138020 5228
rect 138072 5216 138078 5228
rect 169570 5216 169576 5228
rect 138072 5188 169576 5216
rect 138072 5176 138078 5188
rect 169570 5176 169576 5188
rect 169628 5176 169634 5228
rect 28966 5120 38654 5148
rect 15930 5040 15936 5092
rect 15988 5080 15994 5092
rect 28966 5080 28994 5120
rect 15988 5052 28994 5080
rect 38626 5080 38654 5120
rect 59630 5108 59636 5160
rect 59688 5148 59694 5160
rect 129918 5148 129924 5160
rect 59688 5120 129924 5148
rect 59688 5108 59694 5120
rect 129918 5108 129924 5120
rect 129976 5108 129982 5160
rect 142154 5108 142160 5160
rect 142212 5148 142218 5160
rect 220446 5148 220452 5160
rect 142212 5120 220452 5148
rect 142212 5108 142218 5120
rect 220446 5108 220452 5120
rect 220504 5108 220510 5160
rect 46198 5080 46204 5092
rect 38626 5052 46204 5080
rect 15988 5040 15994 5052
rect 46198 5040 46204 5052
rect 46256 5040 46262 5092
rect 52546 5040 52552 5092
rect 52604 5080 52610 5092
rect 128446 5080 128452 5092
rect 52604 5052 128452 5080
rect 52604 5040 52610 5052
rect 128446 5040 128452 5052
rect 128504 5040 128510 5092
rect 136910 5040 136916 5092
rect 136968 5080 136974 5092
rect 148318 5080 148324 5092
rect 136968 5052 148324 5080
rect 136968 5040 136974 5052
rect 148318 5040 148324 5052
rect 148376 5040 148382 5092
rect 154482 5040 154488 5092
rect 154540 5080 154546 5092
rect 365806 5080 365812 5092
rect 154540 5052 365812 5080
rect 154540 5040 154546 5052
rect 365806 5040 365812 5052
rect 365864 5040 365870 5092
rect 33226 4972 33232 5024
rect 33284 5012 33290 5024
rect 127434 5012 127440 5024
rect 33284 4984 127440 5012
rect 33284 4972 33290 4984
rect 127434 4972 127440 4984
rect 127492 4972 127498 5024
rect 138198 4972 138204 5024
rect 138256 5012 138262 5024
rect 171962 5012 171968 5024
rect 138256 4984 171968 5012
rect 138256 4972 138262 4984
rect 171962 4972 171968 4984
rect 172020 4972 172026 5024
rect 180058 4972 180064 5024
rect 180116 5012 180122 5024
rect 450906 5012 450912 5024
rect 180116 4984 450912 5012
rect 180116 4972 180122 4984
rect 450906 4972 450912 4984
rect 450964 4972 450970 5024
rect 6454 4904 6460 4956
rect 6512 4944 6518 4956
rect 22738 4944 22744 4956
rect 6512 4916 22744 4944
rect 6512 4904 6518 4916
rect 22738 4904 22744 4916
rect 22796 4904 22802 4956
rect 24210 4904 24216 4956
rect 24268 4944 24274 4956
rect 122098 4944 122104 4956
rect 24268 4916 122104 4944
rect 24268 4904 24274 4916
rect 122098 4904 122104 4916
rect 122156 4904 122162 4956
rect 137002 4904 137008 4956
rect 137060 4944 137066 4956
rect 150618 4944 150624 4956
rect 137060 4916 150624 4944
rect 137060 4904 137066 4916
rect 150618 4904 150624 4916
rect 150676 4904 150682 4956
rect 162946 4904 162952 4956
rect 163004 4944 163010 4956
rect 487614 4944 487620 4956
rect 163004 4916 487620 4944
rect 163004 4904 163010 4916
rect 487614 4904 487620 4916
rect 487672 4904 487678 4956
rect 13538 4836 13544 4888
rect 13596 4876 13602 4888
rect 125870 4876 125876 4888
rect 13596 4848 125876 4876
rect 13596 4836 13602 4848
rect 125870 4836 125876 4848
rect 125928 4836 125934 4888
rect 137094 4836 137100 4888
rect 137152 4876 137158 4888
rect 157794 4876 157800 4888
rect 137152 4848 157800 4876
rect 137152 4836 137158 4848
rect 157794 4836 157800 4848
rect 157852 4836 157858 4888
rect 165614 4836 165620 4888
rect 165672 4876 165678 4888
rect 523034 4876 523040 4888
rect 165672 4848 523040 4876
rect 165672 4836 165678 4848
rect 523034 4836 523040 4848
rect 523092 4836 523098 4888
rect 8754 4768 8760 4820
rect 8812 4808 8818 4820
rect 125778 4808 125784 4820
rect 8812 4780 125784 4808
rect 8812 4768 8818 4780
rect 125778 4768 125784 4780
rect 125836 4768 125842 4820
rect 138106 4768 138112 4820
rect 138164 4808 138170 4820
rect 164878 4808 164884 4820
rect 138164 4780 164884 4808
rect 138164 4768 138170 4780
rect 164878 4768 164884 4780
rect 164936 4768 164942 4820
rect 165706 4768 165712 4820
rect 165764 4808 165770 4820
rect 527818 4808 527824 4820
rect 165764 4780 527824 4808
rect 165764 4768 165770 4780
rect 527818 4768 527824 4780
rect 527876 4768 527882 4820
rect 138934 4360 138940 4412
rect 138992 4400 138998 4412
rect 143534 4400 143540 4412
rect 138992 4372 143540 4400
rect 138992 4360 138998 4372
rect 143534 4360 143540 4372
rect 143592 4360 143598 4412
rect 242894 4156 242900 4208
rect 242952 4196 242958 4208
rect 244090 4196 244096 4208
rect 242952 4168 244096 4196
rect 242952 4156 242958 4168
rect 244090 4156 244096 4168
rect 244148 4156 244154 4208
rect 251174 4156 251180 4208
rect 251232 4196 251238 4208
rect 252370 4196 252376 4208
rect 251232 4168 252376 4196
rect 251232 4156 251238 4168
rect 252370 4156 252376 4168
rect 252428 4156 252434 4208
rect 276014 4156 276020 4208
rect 276072 4196 276078 4208
rect 276750 4196 276756 4208
rect 276072 4168 276756 4196
rect 276072 4156 276078 4168
rect 276750 4156 276756 4168
rect 276808 4156 276814 4208
rect 119890 4088 119896 4140
rect 119948 4128 119954 4140
rect 124858 4128 124864 4140
rect 119948 4100 124864 4128
rect 119948 4088 119954 4100
rect 124858 4088 124864 4100
rect 124916 4088 124922 4140
rect 125870 4088 125876 4140
rect 125928 4128 125934 4140
rect 134518 4128 134524 4140
rect 125928 4100 134524 4128
rect 125928 4088 125934 4100
rect 134518 4088 134524 4100
rect 134576 4088 134582 4140
rect 151538 4088 151544 4140
rect 151596 4128 151602 4140
rect 325602 4128 325608 4140
rect 151596 4100 325608 4128
rect 151596 4088 151602 4100
rect 325602 4088 325608 4100
rect 325660 4088 325666 4140
rect 138658 4020 138664 4072
rect 138716 4060 138722 4072
rect 145926 4060 145932 4072
rect 138716 4032 145932 4060
rect 138716 4020 138722 4032
rect 145926 4020 145932 4032
rect 145984 4020 145990 4072
rect 150894 4020 150900 4072
rect 150952 4060 150958 4072
rect 327994 4060 328000 4072
rect 150952 4032 328000 4060
rect 150952 4020 150958 4032
rect 327994 4020 328000 4032
rect 328052 4020 328058 4072
rect 12342 3952 12348 4004
rect 12400 3992 12406 4004
rect 126422 3992 126428 4004
rect 12400 3964 126428 3992
rect 12400 3952 12406 3964
rect 126422 3952 126428 3964
rect 126480 3952 126486 4004
rect 150526 3952 150532 4004
rect 150584 3992 150590 4004
rect 331582 3992 331588 4004
rect 150584 3964 331588 3992
rect 150584 3952 150590 3964
rect 331582 3952 331588 3964
rect 331640 3952 331646 4004
rect 136818 3884 136824 3936
rect 136876 3924 136882 3936
rect 144730 3924 144736 3936
rect 136876 3896 144736 3924
rect 136876 3884 136882 3896
rect 144730 3884 144736 3896
rect 144788 3884 144794 3936
rect 172054 3884 172060 3936
rect 172112 3924 172118 3936
rect 356330 3924 356336 3936
rect 172112 3896 356336 3924
rect 172112 3884 172118 3896
rect 356330 3884 356336 3896
rect 356388 3884 356394 3936
rect 467098 3884 467104 3936
rect 467156 3924 467162 3936
rect 534902 3924 534908 3936
rect 467156 3896 534908 3924
rect 467156 3884 467162 3896
rect 534902 3884 534908 3896
rect 534960 3884 534966 3936
rect 83274 3816 83280 3868
rect 83332 3856 83338 3868
rect 131850 3856 131856 3868
rect 83332 3828 131856 3856
rect 83332 3816 83338 3828
rect 131850 3816 131856 3828
rect 131908 3816 131914 3868
rect 142982 3816 142988 3868
rect 143040 3856 143046 3868
rect 151814 3856 151820 3868
rect 143040 3828 151820 3856
rect 143040 3816 143046 3828
rect 151814 3816 151820 3828
rect 151872 3816 151878 3868
rect 172238 3816 172244 3868
rect 172296 3856 172302 3868
rect 303154 3856 303160 3868
rect 172296 3828 303160 3856
rect 172296 3816 172302 3828
rect 303154 3816 303160 3828
rect 303212 3816 303218 3868
rect 319438 3816 319444 3868
rect 319496 3856 319502 3868
rect 583386 3856 583392 3868
rect 319496 3828 583392 3856
rect 319496 3816 319502 3828
rect 583386 3816 583392 3828
rect 583444 3816 583450 3868
rect 76190 3748 76196 3800
rect 76248 3788 76254 3800
rect 128998 3788 129004 3800
rect 76248 3760 129004 3788
rect 76248 3748 76254 3760
rect 128998 3748 129004 3760
rect 129056 3748 129062 3800
rect 140038 3748 140044 3800
rect 140096 3788 140102 3800
rect 149514 3788 149520 3800
rect 140096 3760 149520 3788
rect 140096 3748 140102 3760
rect 149514 3748 149520 3760
rect 149572 3748 149578 3800
rect 152550 3748 152556 3800
rect 152608 3788 152614 3800
rect 168374 3788 168380 3800
rect 152608 3760 168380 3788
rect 152608 3748 152614 3760
rect 168374 3748 168380 3760
rect 168432 3748 168438 3800
rect 178678 3748 178684 3800
rect 178736 3788 178742 3800
rect 475746 3788 475752 3800
rect 178736 3760 475752 3788
rect 178736 3748 178742 3760
rect 475746 3748 475752 3760
rect 475804 3748 475810 3800
rect 69106 3680 69112 3732
rect 69164 3720 69170 3732
rect 130654 3720 130660 3732
rect 69164 3692 130660 3720
rect 69164 3680 69170 3692
rect 130654 3680 130660 3692
rect 130712 3680 130718 3732
rect 137738 3680 137744 3732
rect 137796 3720 137802 3732
rect 154206 3720 154212 3732
rect 137796 3692 154212 3720
rect 137796 3680 137802 3692
rect 154206 3680 154212 3692
rect 154264 3680 154270 3732
rect 163958 3680 163964 3732
rect 164016 3720 164022 3732
rect 491110 3720 491116 3732
rect 164016 3692 491116 3720
rect 164016 3680 164022 3692
rect 491110 3680 491116 3692
rect 491168 3680 491174 3732
rect 62022 3612 62028 3664
rect 62080 3652 62086 3664
rect 122190 3652 122196 3664
rect 62080 3624 122196 3652
rect 62080 3612 62086 3624
rect 122190 3612 122196 3624
rect 122248 3612 122254 3664
rect 127618 3652 127624 3664
rect 122806 3624 127624 3652
rect 47854 3544 47860 3596
rect 47912 3584 47918 3596
rect 122806 3584 122834 3624
rect 127618 3612 127624 3624
rect 127676 3612 127682 3664
rect 136726 3612 136732 3664
rect 136784 3652 136790 3664
rect 155402 3652 155408 3664
rect 136784 3624 155408 3652
rect 136784 3612 136790 3624
rect 155402 3612 155408 3624
rect 155460 3612 155466 3664
rect 171870 3612 171876 3664
rect 171928 3652 171934 3664
rect 501782 3652 501788 3664
rect 171928 3624 501788 3652
rect 171928 3612 171934 3624
rect 501782 3612 501788 3624
rect 501840 3612 501846 3664
rect 47912 3556 122834 3584
rect 47912 3544 47918 3556
rect 126974 3544 126980 3596
rect 127032 3584 127038 3596
rect 130378 3584 130384 3596
rect 127032 3556 130384 3584
rect 127032 3544 127038 3556
rect 130378 3544 130384 3556
rect 130436 3544 130442 3596
rect 133782 3544 133788 3596
rect 133840 3584 133846 3596
rect 147122 3584 147128 3596
rect 133840 3556 147128 3584
rect 133840 3544 133846 3556
rect 147122 3544 147128 3556
rect 147180 3544 147186 3596
rect 147214 3544 147220 3596
rect 147272 3584 147278 3596
rect 167178 3584 167184 3596
rect 147272 3556 167184 3584
rect 147272 3544 147278 3556
rect 167178 3544 167184 3556
rect 167236 3544 167242 3596
rect 171778 3544 171784 3596
rect 171836 3584 171842 3596
rect 515950 3584 515956 3596
rect 171836 3556 515956 3584
rect 171836 3544 171842 3556
rect 515950 3544 515956 3556
rect 516008 3544 516014 3596
rect 17034 3476 17040 3528
rect 17092 3516 17098 3528
rect 125686 3516 125692 3528
rect 17092 3488 125692 3516
rect 17092 3476 17098 3488
rect 125686 3476 125692 3488
rect 125744 3476 125750 3528
rect 131758 3476 131764 3528
rect 131816 3516 131822 3528
rect 135622 3516 135628 3528
rect 131816 3488 135628 3516
rect 131816 3476 131822 3488
rect 135622 3476 135628 3488
rect 135680 3476 135686 3528
rect 141510 3476 141516 3528
rect 141568 3516 141574 3528
rect 166074 3516 166080 3528
rect 141568 3488 166080 3516
rect 141568 3476 141574 3488
rect 166074 3476 166080 3488
rect 166132 3476 166138 3528
rect 173158 3476 173164 3528
rect 173216 3516 173222 3528
rect 173216 3488 531176 3516
rect 173216 3476 173222 3488
rect 93854 3408 93860 3460
rect 93912 3448 93918 3460
rect 94774 3448 94780 3460
rect 93912 3420 94780 3448
rect 93912 3408 93918 3420
rect 94774 3408 94780 3420
rect 94832 3408 94838 3460
rect 142798 3408 142804 3460
rect 142856 3448 142862 3460
rect 170766 3448 170772 3460
rect 142856 3420 170772 3448
rect 142856 3408 142862 3420
rect 170766 3408 170772 3420
rect 170824 3408 170830 3460
rect 173342 3408 173348 3460
rect 173400 3448 173406 3460
rect 531148 3448 531176 3488
rect 531314 3476 531320 3528
rect 531372 3516 531378 3528
rect 532142 3516 532148 3528
rect 531372 3488 532148 3516
rect 531372 3476 531378 3488
rect 532142 3476 532148 3488
rect 532200 3476 532206 3528
rect 539594 3476 539600 3528
rect 539652 3516 539658 3528
rect 540422 3516 540428 3528
rect 539652 3488 540428 3516
rect 539652 3476 539658 3488
rect 540422 3476 540428 3488
rect 540480 3476 540486 3528
rect 533706 3448 533712 3460
rect 173400 3420 528554 3448
rect 531148 3420 533712 3448
rect 173400 3408 173406 3420
rect 150802 3340 150808 3392
rect 150860 3380 150866 3392
rect 322106 3380 322112 3392
rect 150860 3352 322112 3380
rect 150860 3340 150866 3352
rect 322106 3340 322112 3352
rect 322164 3340 322170 3392
rect 340966 3340 340972 3392
rect 341024 3380 341030 3392
rect 342162 3380 342168 3392
rect 341024 3352 342168 3380
rect 341024 3340 341030 3352
rect 342162 3340 342168 3352
rect 342220 3340 342226 3392
rect 349246 3340 349252 3392
rect 349304 3380 349310 3392
rect 350442 3380 350448 3392
rect 349304 3352 350448 3380
rect 349304 3340 349310 3352
rect 350442 3340 350448 3352
rect 350500 3340 350506 3392
rect 357434 3340 357440 3392
rect 357492 3380 357498 3392
rect 358722 3380 358728 3392
rect 357492 3352 358728 3380
rect 357492 3340 357498 3352
rect 358722 3340 358728 3352
rect 358780 3340 358786 3392
rect 365714 3340 365720 3392
rect 365772 3380 365778 3392
rect 367002 3380 367008 3392
rect 365772 3352 367008 3380
rect 365772 3340 365778 3352
rect 367002 3340 367008 3352
rect 367060 3340 367066 3392
rect 374086 3340 374092 3392
rect 374144 3380 374150 3392
rect 375282 3380 375288 3392
rect 374144 3352 375288 3380
rect 374144 3340 374150 3352
rect 375282 3340 375288 3352
rect 375340 3340 375346 3392
rect 382366 3340 382372 3392
rect 382424 3380 382430 3392
rect 383562 3380 383568 3392
rect 382424 3352 383568 3380
rect 382424 3340 382430 3352
rect 383562 3340 383568 3352
rect 383620 3340 383626 3392
rect 398926 3340 398932 3392
rect 398984 3380 398990 3392
rect 400122 3380 400128 3392
rect 398984 3352 400128 3380
rect 398984 3340 398990 3352
rect 400122 3340 400128 3352
rect 400180 3340 400186 3392
rect 415394 3340 415400 3392
rect 415452 3380 415458 3392
rect 416682 3380 416688 3392
rect 415452 3352 416688 3380
rect 415452 3340 415458 3352
rect 416682 3340 416688 3352
rect 416740 3340 416746 3392
rect 423766 3340 423772 3392
rect 423824 3380 423830 3392
rect 424962 3380 424968 3392
rect 423824 3352 424968 3380
rect 423824 3340 423830 3352
rect 424962 3340 424968 3352
rect 425020 3340 425026 3392
rect 448606 3340 448612 3392
rect 448664 3380 448670 3392
rect 449802 3380 449808 3392
rect 448664 3352 449808 3380
rect 448664 3340 448670 3352
rect 449802 3340 449808 3352
rect 449860 3340 449866 3392
rect 456794 3340 456800 3392
rect 456852 3380 456858 3392
rect 458082 3380 458088 3392
rect 456852 3352 458088 3380
rect 456852 3340 456858 3352
rect 458082 3340 458088 3352
rect 458140 3340 458146 3392
rect 506474 3340 506480 3392
rect 506532 3380 506538 3392
rect 507302 3380 507308 3392
rect 506532 3352 507308 3380
rect 506532 3340 506538 3352
rect 507302 3340 507308 3352
rect 507360 3340 507366 3392
rect 528526 3380 528554 3420
rect 533706 3408 533712 3420
rect 533764 3408 533770 3460
rect 537202 3380 537208 3392
rect 528526 3352 537208 3380
rect 537202 3340 537208 3352
rect 537260 3340 537266 3392
rect 135714 3272 135720 3324
rect 135772 3312 135778 3324
rect 138842 3312 138848 3324
rect 135772 3284 138848 3312
rect 135772 3272 135778 3284
rect 138842 3272 138848 3284
rect 138900 3272 138906 3324
rect 144454 3272 144460 3324
rect 144512 3312 144518 3324
rect 153010 3312 153016 3324
rect 144512 3284 153016 3312
rect 144512 3272 144518 3284
rect 153010 3272 153016 3284
rect 153068 3272 153074 3324
rect 173250 3272 173256 3324
rect 173308 3312 173314 3324
rect 212166 3312 212172 3324
rect 173308 3284 212172 3312
rect 173308 3272 173314 3284
rect 212166 3272 212172 3284
rect 212224 3272 212230 3324
rect 362310 3312 362316 3324
rect 219406 3284 362316 3312
rect 211798 3204 211804 3256
rect 211856 3244 211862 3256
rect 219406 3244 219434 3284
rect 362310 3272 362316 3284
rect 362368 3272 362374 3324
rect 211856 3216 219434 3244
rect 211856 3204 211862 3216
rect 307754 3204 307760 3256
rect 307812 3244 307818 3256
rect 309042 3244 309048 3256
rect 307812 3216 309048 3244
rect 307812 3204 307818 3216
rect 309042 3204 309048 3216
rect 309100 3204 309106 3256
rect 316034 3204 316040 3256
rect 316092 3244 316098 3256
rect 317322 3244 317328 3256
rect 316092 3216 317328 3244
rect 316092 3204 316098 3216
rect 317322 3204 317328 3216
rect 317380 3204 317386 3256
rect 135530 3136 135536 3188
rect 135588 3176 135594 3188
rect 140038 3176 140044 3188
rect 135588 3148 140044 3176
rect 135588 3136 135594 3148
rect 140038 3136 140044 3148
rect 140096 3136 140102 3188
rect 132954 3068 132960 3120
rect 133012 3108 133018 3120
rect 135438 3108 135444 3120
rect 133012 3080 135444 3108
rect 133012 3068 133018 3080
rect 135438 3068 135444 3080
rect 135496 3068 135502 3120
rect 135806 3068 135812 3120
rect 135864 3108 135870 3120
rect 137646 3108 137652 3120
rect 135864 3080 137652 3108
rect 135864 3068 135870 3080
rect 137646 3068 137652 3080
rect 137704 3068 137710 3120
rect 135898 3000 135904 3052
rect 135956 3040 135962 3052
rect 141234 3040 141240 3052
rect 135956 3012 141240 3040
rect 135956 3000 135962 3012
rect 141234 3000 141240 3012
rect 141292 3000 141298 3052
rect 390554 1232 390560 1284
rect 390612 1272 390618 1284
rect 391842 1272 391848 1284
rect 390612 1244 391848 1272
rect 390612 1232 390618 1244
rect 391842 1232 391848 1244
rect 391900 1232 391906 1284
rect 30098 1096 30104 1148
rect 30156 1136 30162 1148
rect 33226 1136 33232 1148
rect 30156 1108 33232 1136
rect 30156 1096 30162 1108
rect 33226 1096 33232 1108
rect 33284 1096 33290 1148
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 331220 702992 331272 703044
rect 332508 702992 332560 703044
rect 410524 700408 410576 700460
rect 429844 700408 429896 700460
rect 300124 700340 300176 700392
rect 303252 700340 303304 700392
rect 409144 700340 409196 700392
rect 494796 700340 494848 700392
rect 254584 700272 254636 700324
rect 267648 700272 267700 700324
rect 407764 700272 407816 700324
rect 559656 700272 559708 700324
rect 348792 699796 348844 699848
rect 351184 699796 351236 699848
rect 152464 699660 152516 699712
rect 154120 699660 154172 699712
rect 196624 699660 196676 699712
rect 202788 699660 202840 699712
rect 217324 699660 217376 699712
rect 218980 699660 219032 699712
rect 282184 697552 282236 697604
rect 283840 697552 283892 697604
rect 303252 693404 303304 693456
rect 316040 693404 316092 693456
rect 351184 692044 351236 692096
rect 358084 692044 358136 692096
rect 364340 690412 364392 690464
rect 369860 690412 369912 690464
rect 150440 689256 150492 689308
rect 152464 689256 152516 689308
rect 239036 689256 239088 689308
rect 254584 689256 254636 689308
rect 331220 688848 331272 688900
rect 334624 688848 334676 688900
rect 213184 688576 213236 688628
rect 217324 688644 217376 688696
rect 316040 688168 316092 688220
rect 323584 688168 323636 688220
rect 369860 688168 369912 688220
rect 372620 688168 372672 688220
rect 224224 685108 224276 685160
rect 239036 685108 239088 685160
rect 2780 683680 2832 683732
rect 4804 683680 4856 683732
rect 149060 683680 149112 683732
rect 150440 683680 150492 683732
rect 372620 683612 372672 683664
rect 375380 683612 375432 683664
rect 358084 681028 358136 681080
rect 360476 681028 360528 681080
rect 261484 680960 261536 681012
rect 282184 680960 282236 681012
rect 375380 680960 375432 681012
rect 389180 680960 389232 681012
rect 360476 678240 360528 678292
rect 369124 678240 369176 678292
rect 146208 676336 146260 676388
rect 148968 676336 149020 676388
rect 369124 675452 369176 675504
rect 378784 675452 378836 675504
rect 389180 675180 389232 675232
rect 393320 675180 393372 675232
rect 143540 674432 143592 674484
rect 146208 674432 146260 674484
rect 220820 673752 220872 673804
rect 224224 673752 224276 673804
rect 393320 673208 393372 673260
rect 396448 673208 396500 673260
rect 211528 672052 211580 672104
rect 213184 672052 213236 672104
rect 3516 670692 3568 670744
rect 15844 670692 15896 670744
rect 208400 670692 208452 670744
rect 211528 670692 211580 670744
rect 406384 670692 406436 670744
rect 580172 670692 580224 670744
rect 140044 667836 140096 667888
rect 143540 667904 143592 667956
rect 218704 667632 218756 667684
rect 220820 667632 220872 667684
rect 258724 666476 258776 666528
rect 261484 666544 261536 666596
rect 206284 665864 206336 665916
rect 208308 665864 208360 665916
rect 378784 664436 378836 664488
rect 387064 664436 387116 664488
rect 215300 662396 215352 662448
rect 218704 662396 218756 662448
rect 323584 662328 323636 662380
rect 326620 662328 326672 662380
rect 326620 659200 326672 659252
rect 330024 659200 330076 659252
rect 211804 657568 211856 657620
rect 215300 657568 215352 657620
rect 330024 656140 330076 656192
rect 336740 656140 336792 656192
rect 257436 654100 257488 654152
rect 258724 654100 258776 654152
rect 387064 652264 387116 652316
rect 395344 652264 395396 652316
rect 138664 651380 138716 651432
rect 140044 651380 140096 651432
rect 255320 651380 255372 651432
rect 257436 651380 257488 651432
rect 336740 649272 336792 649324
rect 345664 649272 345716 649324
rect 201408 647844 201460 647896
rect 211804 647844 211856 647896
rect 204904 647164 204956 647216
rect 206284 647164 206336 647216
rect 334624 646484 334676 646536
rect 342904 646484 342956 646536
rect 189724 645124 189776 645176
rect 201408 645124 201460 645176
rect 245568 645124 245620 645176
rect 255320 645124 255372 645176
rect 345664 644308 345716 644360
rect 353944 644308 353996 644360
rect 135904 641724 135956 641776
rect 138664 641724 138716 641776
rect 243544 640296 243596 640348
rect 245568 640296 245620 640348
rect 179420 636828 179472 636880
rect 189724 636828 189776 636880
rect 2780 632068 2832 632120
rect 4896 632068 4948 632120
rect 174452 630640 174504 630692
rect 179420 630640 179472 630692
rect 171784 629008 171836 629060
rect 174452 629008 174504 629060
rect 193864 623772 193916 623824
rect 196624 623772 196676 623824
rect 239956 623704 240008 623756
rect 243544 623772 243596 623824
rect 353944 622344 353996 622396
rect 356704 622344 356756 622396
rect 237380 620984 237432 621036
rect 239956 620984 240008 621036
rect 3516 618264 3568 618316
rect 19984 618264 20036 618316
rect 233884 616768 233936 616820
rect 237380 616836 237432 616888
rect 405004 616836 405056 616888
rect 579712 616836 579764 616888
rect 342904 616088 342956 616140
rect 360844 616088 360896 616140
rect 191104 610648 191156 610700
rect 193864 610648 193916 610700
rect 232596 610240 232648 610292
rect 234620 610240 234672 610292
rect 356704 607860 356756 607912
rect 369124 607860 369176 607912
rect 153844 605072 153896 605124
rect 171784 605072 171836 605124
rect 134524 603100 134576 603152
rect 135904 603100 135956 603152
rect 232504 603100 232556 603152
rect 233884 603100 233936 603152
rect 203616 601672 203668 601724
rect 204904 601672 204956 601724
rect 224408 600924 224460 600976
rect 232596 600924 232648 600976
rect 184204 599836 184256 599888
rect 191104 599836 191156 599888
rect 202144 599632 202196 599684
rect 203616 599632 203668 599684
rect 220820 598136 220872 598188
rect 224408 598136 224460 598188
rect 214564 594804 214616 594856
rect 220820 594804 220872 594856
rect 360844 594396 360896 594448
rect 366364 594396 366416 594448
rect 181444 592016 181496 592068
rect 184204 592016 184256 592068
rect 369124 590588 369176 590640
rect 371884 590588 371936 590640
rect 371884 585760 371936 585812
rect 380164 585760 380216 585812
rect 130384 583652 130436 583704
rect 134524 583720 134576 583772
rect 3516 579640 3568 579692
rect 10324 579640 10376 579692
rect 211804 578144 211856 578196
rect 214564 578144 214616 578196
rect 149060 575220 149112 575272
rect 153844 575220 153896 575272
rect 366364 574064 366416 574116
rect 369124 574064 369176 574116
rect 231124 572704 231176 572756
rect 232504 572704 232556 572756
rect 137284 571956 137336 572008
rect 149060 571956 149112 572008
rect 380164 570596 380216 570648
rect 392584 570596 392636 570648
rect 127624 567808 127676 567860
rect 137284 567808 137336 567860
rect 3056 565836 3108 565888
rect 37924 565836 37976 565888
rect 209044 564952 209096 565004
rect 211804 564952 211856 565004
rect 229928 564680 229980 564732
rect 231124 564680 231176 564732
rect 392584 564340 392636 564392
rect 395436 564340 395488 564392
rect 403624 563048 403676 563100
rect 580172 563048 580224 563100
rect 228364 562640 228416 562692
rect 229928 562640 229980 562692
rect 189080 560940 189132 560992
rect 202144 560940 202196 560992
rect 184940 558968 184992 559020
rect 189080 558968 189132 559020
rect 124864 558832 124916 558884
rect 127624 558832 127676 558884
rect 201224 556180 201276 556232
rect 209044 556180 209096 556232
rect 163504 554004 163556 554056
rect 181444 554004 181496 554056
rect 193864 552848 193916 552900
rect 201224 552848 201276 552900
rect 183192 552644 183244 552696
rect 184848 552644 184900 552696
rect 226984 552644 227036 552696
rect 228364 552644 228416 552696
rect 181444 550400 181496 550452
rect 183192 550400 183244 550452
rect 129004 550196 129056 550248
rect 130384 550196 130436 550248
rect 146116 547136 146168 547188
rect 163504 547136 163556 547188
rect 224960 546456 225012 546508
rect 226984 546456 227036 546508
rect 170404 545708 170456 545760
rect 193864 545708 193916 545760
rect 122104 545572 122156 545624
rect 124864 545572 124916 545624
rect 133144 544348 133196 544400
rect 146116 544348 146168 544400
rect 223028 540064 223080 540116
rect 224868 540064 224920 540116
rect 156604 537480 156656 537532
rect 170404 537480 170456 537532
rect 123484 536052 123536 536104
rect 133144 536052 133196 536104
rect 220360 535440 220412 535492
rect 223028 535440 223080 535492
rect 180064 534012 180116 534064
rect 181444 534012 181496 534064
rect 218704 532312 218756 532364
rect 220360 532312 220412 532364
rect 117136 527144 117188 527196
rect 122104 527144 122156 527196
rect 106924 525036 106976 525088
rect 129004 525036 129056 525088
rect 101404 519528 101456 519580
rect 117136 519528 117188 519580
rect 127624 516740 127676 516792
rect 156604 516740 156656 516792
rect 3332 514768 3384 514820
rect 43444 514768 43496 514820
rect 105544 514020 105596 514072
rect 106924 514020 106976 514072
rect 98644 511912 98696 511964
rect 101404 511912 101456 511964
rect 400864 510620 400916 510672
rect 580172 510620 580224 510672
rect 113824 508512 113876 508564
rect 123484 508512 123536 508564
rect 178684 505112 178736 505164
rect 180064 505112 180116 505164
rect 102784 499536 102836 499588
rect 105544 499536 105596 499588
rect 175280 498176 175332 498228
rect 178684 498176 178736 498228
rect 173164 493280 173216 493332
rect 175188 493280 175240 493332
rect 217324 493280 217376 493332
rect 218704 493280 218756 493332
rect 369124 490356 369176 490408
rect 376024 490356 376076 490408
rect 171140 482808 171192 482860
rect 173164 482808 173216 482860
rect 215944 482672 215996 482724
rect 217324 482672 217376 482724
rect 119344 482264 119396 482316
rect 127624 482264 127676 482316
rect 171140 478864 171192 478916
rect 167644 478796 167696 478848
rect 101404 477504 101456 477556
rect 102784 477504 102836 477556
rect 116584 469208 116636 469260
rect 119344 469208 119396 469260
rect 213184 469208 213236 469260
rect 215944 469208 215996 469260
rect 95884 466420 95936 466472
rect 98644 466420 98696 466472
rect 2780 462544 2832 462596
rect 4988 462544 5040 462596
rect 399484 456764 399536 456816
rect 580172 456764 580224 456816
rect 376024 456016 376076 456068
rect 385684 456016 385736 456068
rect 210516 453976 210568 454028
rect 213184 454044 213236 454096
rect 97264 452548 97316 452600
rect 101404 452616 101456 452668
rect 108304 447720 108356 447772
rect 113824 447720 113876 447772
rect 209044 446360 209096 446412
rect 210516 446360 210568 446412
rect 207664 438880 207716 438932
rect 209044 438880 209096 438932
rect 204904 430584 204956 430636
rect 207664 430584 207716 430636
rect 396724 430584 396776 430636
rect 579988 430584 580040 430636
rect 93124 429700 93176 429752
rect 95884 429700 95936 429752
rect 100024 424328 100076 424380
rect 108304 424328 108356 424380
rect 166264 423580 166316 423632
rect 167644 423580 167696 423632
rect 3148 422900 3200 422952
rect 6184 422900 6236 422952
rect 398104 418140 398156 418192
rect 580172 418140 580224 418192
rect 164792 415080 164844 415132
rect 166264 415080 166316 415132
rect 95884 415012 95936 415064
rect 97264 415012 97316 415064
rect 108304 411884 108356 411936
rect 116584 411884 116636 411936
rect 3332 409912 3384 409964
rect 8944 409912 8996 409964
rect 161848 407124 161900 407176
rect 164792 407124 164844 407176
rect 93216 406376 93268 406428
rect 100024 406376 100076 406428
rect 160100 406376 160152 406428
rect 161848 406376 161900 406428
rect 157340 404268 157392 404320
rect 160100 404336 160152 404388
rect 421564 404336 421616 404388
rect 580172 404336 580224 404388
rect 153844 400120 153896 400172
rect 157340 400188 157392 400240
rect 69664 396720 69716 396772
rect 136640 396720 136692 396772
rect 105544 394612 105596 394664
rect 108304 394612 108356 394664
rect 93308 393320 93360 393372
rect 95884 393320 95936 393372
rect 146944 391892 146996 391944
rect 153844 391960 153896 392012
rect 385684 388492 385736 388544
rect 389272 388492 389324 388544
rect 199384 388424 199436 388476
rect 204904 388424 204956 388476
rect 97540 385024 97592 385076
rect 105544 385024 105596 385076
rect 68284 384956 68336 385008
rect 69664 384956 69716 385008
rect 389272 384956 389324 385008
rect 392768 384956 392820 385008
rect 88984 384412 89036 384464
rect 93216 384412 93268 384464
rect 86868 382916 86920 382968
rect 97540 382916 97592 382968
rect 392768 382168 392820 382220
rect 395528 382168 395580 382220
rect 91928 379516 91980 379568
rect 93308 379516 93360 379568
rect 79324 379040 79376 379092
rect 86868 379040 86920 379092
rect 396908 378156 396960 378208
rect 579804 378156 579856 378208
rect 90364 377816 90416 377868
rect 91928 377816 91980 377868
rect 197360 372580 197412 372632
rect 199384 372580 199436 372632
rect 3332 371220 3384 371272
rect 10416 371220 10468 371272
rect 192484 369792 192536 369844
rect 197360 369860 197412 369912
rect 87512 364488 87564 364540
rect 90364 364488 90416 364540
rect 73804 359456 73856 359508
rect 88984 359456 89036 359508
rect 65708 359048 65760 359100
rect 68284 359048 68336 359100
rect 86224 358912 86276 358964
rect 87512 358912 87564 358964
rect 142804 358708 142856 358760
rect 146944 358776 146996 358828
rect 64144 358164 64196 358216
rect 65708 358164 65760 358216
rect 54484 358028 54536 358080
rect 79324 358028 79376 358080
rect 3332 357416 3384 357468
rect 24124 357416 24176 357468
rect 85028 353268 85080 353320
rect 86224 353268 86276 353320
rect 140780 353268 140832 353320
rect 142804 353268 142856 353320
rect 418804 351908 418856 351960
rect 580080 351908 580132 351960
rect 82820 351296 82872 351348
rect 85028 351296 85080 351348
rect 137284 350548 137336 350600
rect 140780 350548 140832 350600
rect 51724 349460 51776 349512
rect 54484 349460 54536 349512
rect 78680 346332 78732 346384
rect 82820 346400 82872 346452
rect 2780 345176 2832 345228
rect 5080 345176 5132 345228
rect 189724 345040 189776 345092
rect 192484 345040 192536 345092
rect 395528 343612 395580 343664
rect 397552 343612 397604 343664
rect 75920 340892 75972 340944
rect 78588 340892 78640 340944
rect 62120 340144 62172 340196
rect 73804 340144 73856 340196
rect 53840 337356 53892 337408
rect 62120 337356 62172 337408
rect 73160 336744 73212 336796
rect 75828 336744 75880 336796
rect 186228 336676 186280 336728
rect 189724 336744 189776 336796
rect 46388 333956 46440 334008
rect 53840 333956 53892 334008
rect 70308 332528 70360 332580
rect 73068 332596 73120 332648
rect 62856 331848 62908 331900
rect 88340 331848 88392 331900
rect 44916 331508 44968 331560
rect 46388 331508 46440 331560
rect 45008 330488 45060 330540
rect 51724 330488 51776 330540
rect 183560 330012 183612 330064
rect 186228 330012 186280 330064
rect 134524 329536 134576 329588
rect 137284 329536 137336 329588
rect 68192 328040 68244 328092
rect 70308 328040 70360 328092
rect 182824 326408 182876 326460
rect 183560 326408 183612 326460
rect 397092 324300 397144 324352
rect 580080 324300 580132 324352
rect 66904 320084 66956 320136
rect 68192 320084 68244 320136
rect 126244 320084 126296 320136
rect 134524 320152 134576 320204
rect 62764 319404 62816 319456
rect 64144 319404 64196 319456
rect 3148 318792 3200 318844
rect 33784 318792 33836 318844
rect 61476 318384 61528 318436
rect 62856 318384 62908 318436
rect 84844 315256 84896 315308
rect 104900 315256 104952 315308
rect 62120 312128 62172 312180
rect 66904 312128 66956 312180
rect 90364 311856 90416 311908
rect 93124 311856 93176 311908
rect 398196 311856 398248 311908
rect 580080 311856 580132 311908
rect 60004 311176 60056 311228
rect 61476 311176 61528 311228
rect 60096 307232 60148 307284
rect 62120 307232 62172 307284
rect 179604 306348 179656 306400
rect 182824 306348 182876 306400
rect 178684 301384 178736 301436
rect 179604 301384 179656 301436
rect 61568 299072 61620 299124
rect 62764 299072 62816 299124
rect 417424 298120 417476 298172
rect 580080 298120 580132 298172
rect 73160 294584 73212 294636
rect 90364 294584 90416 294636
rect 60188 293972 60240 294024
rect 61568 293972 61620 294024
rect 175280 293972 175332 294024
rect 178684 293972 178736 294024
rect 124864 292544 124916 292596
rect 126244 292544 126296 292596
rect 66996 291184 67048 291236
rect 73160 291184 73212 291236
rect 58624 291116 58676 291168
rect 60004 291116 60056 291168
rect 55220 289756 55272 289808
rect 60096 289824 60148 289876
rect 55864 289076 55916 289128
rect 66996 289076 67048 289128
rect 57244 287648 57296 287700
rect 71780 287648 71832 287700
rect 56508 284248 56560 284300
rect 58624 284316 58676 284368
rect 82084 284248 82136 284300
rect 84844 284316 84896 284368
rect 57980 282888 58032 282940
rect 60188 282888 60240 282940
rect 173164 281800 173216 281852
rect 174912 281800 174964 281852
rect 54208 281392 54260 281444
rect 56508 281392 56560 281444
rect 53288 280780 53340 280832
rect 169760 280780 169812 280832
rect 53380 280168 53432 280220
rect 55128 280168 55180 280220
rect 53104 279420 53156 279472
rect 54208 279420 54260 279472
rect 54484 278740 54536 278792
rect 57888 278740 57940 278792
rect 53840 277312 53892 277364
rect 57244 277380 57296 277432
rect 55956 276632 56008 276684
rect 82084 276632 82136 276684
rect 50344 274864 50396 274916
rect 55864 274864 55916 274916
rect 50436 274728 50488 274780
rect 53380 274728 53432 274780
rect 53196 274660 53248 274712
rect 53840 274660 53892 274712
rect 118700 273164 118752 273216
rect 124864 273232 124916 273284
rect 51724 272008 51776 272060
rect 53104 272008 53156 272060
rect 396816 271872 396868 271924
rect 579804 271872 579856 271924
rect 167644 271804 167696 271856
rect 173164 271804 173216 271856
rect 116768 270512 116820 270564
rect 118700 270512 118752 270564
rect 51080 270444 51132 270496
rect 53288 270444 53340 270496
rect 45284 268336 45336 268388
rect 50344 268336 50396 268388
rect 112168 268336 112220 268388
rect 116768 268336 116820 268388
rect 3148 266704 3200 266756
rect 9036 266704 9088 266756
rect 165620 266568 165672 266620
rect 167644 266568 167696 266620
rect 53196 266432 53248 266484
rect 54484 266432 54536 266484
rect 46204 266296 46256 266348
rect 50436 266364 50488 266416
rect 48320 266296 48372 266348
rect 51080 266364 51132 266416
rect 54208 266364 54260 266416
rect 55956 266364 56008 266416
rect 109040 266364 109092 266416
rect 112168 266364 112220 266416
rect 158720 265616 158772 265668
rect 165620 265616 165672 265668
rect 49700 263576 49752 263628
rect 51724 263576 51776 263628
rect 53288 263576 53340 263628
rect 54208 263576 54260 263628
rect 107016 260448 107068 260500
rect 108948 260448 109000 260500
rect 151820 259224 151872 259276
rect 158720 259224 158772 259276
rect 45744 259088 45796 259140
rect 48228 259088 48280 259140
rect 46940 258544 46992 258596
rect 49700 258544 49752 258596
rect 418896 258068 418948 258120
rect 579988 258068 580040 258120
rect 45192 256708 45244 256760
rect 46204 256708 46256 256760
rect 50436 256640 50488 256692
rect 53288 256708 53340 256760
rect 104900 256708 104952 256760
rect 107016 256708 107068 256760
rect 45652 255280 45704 255332
rect 46940 255280 46992 255332
rect 101404 255212 101456 255264
rect 104900 255280 104952 255332
rect 3148 253920 3200 253972
rect 22744 253920 22796 253972
rect 46204 253852 46256 253904
rect 53196 253988 53248 254040
rect 47584 253920 47636 253972
rect 50436 253920 50488 253972
rect 146944 253852 146996 253904
rect 151728 253920 151780 253972
rect 51080 252832 51132 252884
rect 53104 252832 53156 252884
rect 50344 250384 50396 250436
rect 51080 250384 51132 250436
rect 143264 247052 143316 247104
rect 146944 247052 146996 247104
rect 45836 245624 45888 245676
rect 47584 245624 47636 245676
rect 44824 244944 44876 244996
rect 46204 244944 46256 244996
rect 414664 244264 414716 244316
rect 579988 244264 580040 244316
rect 45100 240796 45152 240848
rect 101404 240796 101456 240848
rect 45468 240728 45520 240780
rect 143264 240728 143316 240780
rect 45652 240524 45704 240576
rect 50344 240524 50396 240576
rect 2780 240184 2832 240236
rect 5172 240184 5224 240236
rect 395436 240048 395488 240100
rect 396540 240048 396592 240100
rect 395344 239776 395396 239828
rect 45376 238756 45428 238808
rect 45836 238756 45888 238808
rect 396540 238756 396592 238808
rect 396632 238688 396684 238740
rect 396540 238620 396592 238672
rect 45744 233316 45796 233368
rect 45560 233248 45612 233300
rect 45376 233180 45428 233232
rect 45100 233112 45152 233164
rect 45836 233112 45888 233164
rect 45560 232840 45612 232892
rect 45468 232772 45520 232824
rect 45744 232772 45796 232824
rect 62764 232364 62816 232416
rect 82084 232364 82136 232416
rect 395436 232364 395488 232416
rect 396632 232364 396684 232416
rect 395344 232296 395396 232348
rect 396448 232296 396500 232348
rect 391204 232228 391256 232280
rect 396540 232228 396592 232280
rect 393964 231820 394016 231872
rect 580080 231820 580132 231872
rect 45836 231140 45888 231192
rect 134156 231140 134208 231192
rect 4068 231072 4120 231124
rect 180800 231072 180852 231124
rect 44824 231004 44876 231056
rect 84844 231004 84896 231056
rect 44916 230528 44968 230580
rect 47676 230528 47728 230580
rect 45744 230392 45796 230444
rect 47584 230392 47636 230444
rect 45560 230324 45612 230376
rect 55128 230324 55180 230376
rect 134156 230052 134208 230104
rect 136364 230052 136416 230104
rect 3884 229712 3936 229764
rect 179420 229712 179472 229764
rect 45008 228352 45060 228404
rect 49976 228352 50028 228404
rect 157984 228352 158036 228404
rect 266544 228352 266596 228404
rect 267004 228352 267056 228404
rect 356520 228352 356572 228404
rect 3148 227740 3200 227792
rect 138664 227740 138716 227792
rect 388444 227740 388496 227792
rect 391204 227740 391256 227792
rect 391296 227740 391348 227792
rect 395436 227740 395488 227792
rect 82084 227672 82136 227724
rect 85488 227672 85540 227724
rect 62764 227128 62816 227180
rect 65800 227128 65852 227180
rect 45192 226244 45244 226296
rect 48228 226244 48280 226296
rect 136364 225156 136416 225208
rect 138756 225156 138808 225208
rect 49976 224952 50028 225004
rect 53840 224952 53892 225004
rect 389088 224952 389140 225004
rect 391296 224952 391348 225004
rect 85488 224204 85540 224256
rect 100024 224204 100076 224256
rect 55220 224136 55272 224188
rect 59360 224136 59412 224188
rect 394056 223524 394108 223576
rect 395344 223524 395396 223576
rect 118700 222844 118752 222896
rect 580172 222844 580224 222896
rect 48228 222164 48280 222216
rect 47584 222096 47636 222148
rect 48320 222096 48372 222148
rect 53196 222096 53248 222148
rect 65800 222096 65852 222148
rect 69664 222096 69716 222148
rect 53840 221416 53892 221468
rect 59268 221416 59320 221468
rect 59360 220736 59412 220788
rect 62764 220736 62816 220788
rect 84844 220736 84896 220788
rect 85764 220736 85816 220788
rect 385040 220736 385092 220788
rect 389088 220736 389140 220788
rect 48320 219444 48372 219496
rect 55128 219376 55180 219428
rect 138756 218696 138808 218748
rect 158720 218696 158772 218748
rect 394424 218084 394476 218136
rect 397552 218084 397604 218136
rect 85764 218016 85816 218068
rect 87604 218016 87656 218068
rect 118608 218016 118660 218068
rect 579988 218016 580040 218068
rect 380900 217880 380952 217932
rect 385040 217880 385092 217932
rect 45284 217608 45336 217660
rect 47584 217608 47636 217660
rect 47676 216724 47728 216776
rect 50344 216724 50396 216776
rect 158720 215976 158772 216028
rect 162768 215976 162820 216028
rect 100024 215908 100076 215960
rect 111064 215908 111116 215960
rect 59268 215704 59320 215756
rect 61384 215704 61436 215756
rect 375472 215432 375524 215484
rect 380900 215432 380952 215484
rect 53196 215228 53248 215280
rect 53840 215228 53892 215280
rect 3148 213936 3200 213988
rect 179512 213936 179564 213988
rect 371884 213868 371936 213920
rect 375472 213936 375524 213988
rect 55220 213188 55272 213240
rect 68284 213188 68336 213240
rect 391204 213120 391256 213172
rect 394424 213120 394476 213172
rect 162768 212848 162820 212900
rect 164884 212848 164936 212900
rect 53840 211692 53892 211744
rect 55220 211692 55272 211744
rect 69664 209516 69716 209568
rect 77024 209516 77076 209568
rect 55220 208836 55272 208888
rect 56876 208836 56928 208888
rect 164884 208360 164936 208412
rect 166264 208360 166316 208412
rect 45560 207612 45612 207664
rect 50436 207612 50488 207664
rect 77024 205776 77076 205828
rect 78680 205776 78732 205828
rect 50344 205708 50396 205760
rect 54484 205708 54536 205760
rect 370504 205708 370556 205760
rect 371884 205708 371936 205760
rect 56876 205640 56928 205692
rect 188344 205640 188396 205692
rect 580172 205640 580224 205692
rect 60004 205572 60056 205624
rect 384396 205436 384448 205488
rect 388444 205436 388496 205488
rect 61384 204892 61436 204944
rect 75184 204892 75236 204944
rect 68284 204212 68336 204264
rect 69664 204212 69716 204264
rect 385684 204212 385736 204264
rect 391204 204212 391256 204264
rect 382924 203328 382976 203380
rect 384396 203328 384448 203380
rect 87604 202784 87656 202836
rect 93124 202784 93176 202836
rect 78680 202104 78732 202156
rect 88064 202104 88116 202156
rect 111064 202104 111116 202156
rect 126888 202104 126940 202156
rect 147772 202104 147824 202156
rect 176660 202104 176712 202156
rect 50436 201900 50488 201952
rect 57244 201900 57296 201952
rect 3148 201832 3200 201884
rect 7564 201832 7616 201884
rect 155960 199384 156012 199436
rect 296720 199384 296772 199436
rect 88064 198704 88116 198756
rect 90364 198704 90416 198756
rect 148968 197956 149020 198008
rect 207020 197956 207072 198008
rect 154488 197412 154540 197464
rect 155960 197412 156012 197464
rect 166264 197344 166316 197396
rect 167644 197344 167696 197396
rect 60004 197276 60056 197328
rect 65524 197276 65576 197328
rect 152740 197276 152792 197328
rect 157984 197276 158036 197328
rect 380900 196868 380952 196920
rect 382924 196868 382976 196920
rect 138664 196732 138716 196784
rect 164240 196732 164292 196784
rect 151176 196664 151228 196716
rect 236000 196664 236052 196716
rect 155960 196596 156012 196648
rect 327080 196596 327132 196648
rect 126888 196324 126940 196376
rect 129004 196324 129056 196376
rect 56600 195916 56652 195968
rect 138112 195916 138164 195968
rect 160100 195916 160152 195968
rect 386420 195916 386472 195968
rect 86960 195848 87012 195900
rect 139400 195848 139452 195900
rect 157616 195848 157668 195900
rect 267004 195848 267056 195900
rect 115940 194556 115992 194608
rect 140780 194556 140832 194608
rect 47584 194488 47636 194540
rect 54576 194488 54628 194540
rect 380164 193944 380216 193996
rect 385684 193944 385736 193996
rect 166172 193808 166224 193860
rect 380900 193808 380952 193860
rect 54484 192448 54536 192500
rect 58624 192448 58676 192500
rect 180064 191836 180116 191888
rect 580172 191836 580224 191888
rect 144736 190476 144788 190528
rect 145012 190272 145064 190324
rect 54576 189728 54628 189780
rect 60740 189728 60792 189780
rect 93124 189252 93176 189304
rect 94504 189252 94556 189304
rect 387064 189048 387116 189100
rect 394056 189048 394108 189100
rect 144736 188912 144788 188964
rect 145012 188912 145064 188964
rect 75184 187756 75236 187808
rect 80060 187756 80112 187808
rect 2780 187688 2832 187740
rect 5264 187688 5316 187740
rect 69664 186328 69716 186380
rect 71136 186328 71188 186380
rect 62764 186056 62816 186108
rect 64144 186056 64196 186108
rect 129004 185580 129056 185632
rect 132408 185580 132460 185632
rect 60740 184832 60792 184884
rect 65616 184832 65668 184884
rect 94504 184832 94556 184884
rect 97264 184832 97316 184884
rect 57244 184152 57296 184204
rect 65800 184152 65852 184204
rect 71136 183472 71188 183524
rect 72516 183472 72568 183524
rect 167644 183472 167696 183524
rect 169116 183472 169168 183524
rect 132408 183268 132460 183320
rect 135904 183268 135956 183320
rect 80060 182792 80112 182844
rect 88984 182792 89036 182844
rect 58624 182452 58676 182504
rect 64880 182452 64932 182504
rect 90364 181432 90416 181484
rect 100024 181432 100076 181484
rect 144920 180956 144972 181008
rect 153936 180752 153988 180804
rect 154396 180616 154448 180668
rect 65800 180548 65852 180600
rect 68376 180548 68428 180600
rect 121460 180072 121512 180124
rect 136364 180072 136416 180124
rect 157800 180072 157852 180124
rect 158628 180072 158680 180124
rect 165620 180072 165672 180124
rect 65524 179868 65576 179920
rect 66996 179868 67048 179920
rect 135996 178848 136048 178900
rect 136548 178848 136600 178900
rect 122840 178644 122892 178696
rect 136456 178644 136508 178696
rect 72516 178032 72568 178084
rect 73804 178032 73856 178084
rect 166540 178032 166592 178084
rect 580172 178032 580224 178084
rect 159456 177828 159508 177880
rect 167644 177828 167696 177880
rect 124220 177284 124272 177336
rect 135996 177284 136048 177336
rect 64880 177148 64932 177200
rect 68468 177148 68520 177200
rect 149336 176468 149388 176520
rect 153936 176400 153988 176452
rect 154396 176400 154448 176452
rect 126980 176060 127032 176112
rect 136272 176060 136324 176112
rect 125600 175924 125652 175976
rect 136180 175924 136232 175976
rect 144092 175924 144144 175976
rect 149336 175924 149388 175976
rect 169116 176332 169168 176384
rect 169760 176332 169812 176384
rect 162492 175924 162544 175976
rect 144460 175516 144512 175568
rect 149980 175516 150032 175568
rect 128360 175176 128412 175228
rect 136364 175176 136416 175228
rect 141608 174700 141660 174752
rect 143080 174700 143132 174752
rect 152464 174632 152516 174684
rect 156512 174632 156564 174684
rect 161480 174496 161532 174548
rect 366364 174496 366416 174548
rect 380164 174496 380216 174548
rect 385684 174496 385736 174548
rect 387064 174496 387116 174548
rect 167000 174292 167052 174344
rect 133880 173884 133932 173936
rect 137376 173884 137428 173936
rect 135904 173136 135956 173188
rect 148324 172932 148376 172984
rect 149060 172932 149112 172984
rect 149336 172932 149388 172984
rect 151452 172932 151504 172984
rect 162492 172932 162544 172984
rect 165436 172932 165488 172984
rect 148968 172864 149020 172916
rect 131120 172524 131172 172576
rect 136548 172524 136600 172576
rect 66996 172456 67048 172508
rect 68284 172456 68336 172508
rect 65616 172388 65668 172440
rect 71044 172388 71096 172440
rect 138020 172116 138072 172168
rect 140780 172116 140832 172168
rect 135260 171640 135312 171692
rect 138664 171640 138716 171692
rect 169760 171368 169812 171420
rect 171784 171368 171836 171420
rect 132500 171096 132552 171148
rect 136732 171096 136784 171148
rect 148968 170348 149020 170400
rect 162676 170348 162728 170400
rect 118424 168988 118476 169040
rect 158444 168988 158496 169040
rect 68468 168036 68520 168088
rect 71504 168036 71556 168088
rect 162676 167696 162728 167748
rect 172244 167696 172296 167748
rect 118792 167628 118844 167680
rect 580264 167628 580316 167680
rect 384304 167084 384356 167136
rect 385684 167084 385736 167136
rect 68376 166948 68428 167000
rect 71780 166948 71832 167000
rect 142436 166268 142488 166320
rect 142620 166268 142672 166320
rect 226984 165588 227036 165640
rect 580172 165588 580224 165640
rect 97264 165520 97316 165572
rect 98644 165520 98696 165572
rect 380900 165248 380952 165300
rect 384304 165248 384356 165300
rect 172244 164160 172296 164212
rect 175188 164160 175240 164212
rect 71504 163548 71556 163600
rect 82820 163548 82872 163600
rect 71780 163480 71832 163532
rect 86224 163480 86276 163532
rect 380256 163072 380308 163124
rect 380900 163072 380952 163124
rect 3148 162868 3200 162920
rect 180892 162868 180944 162920
rect 9036 162120 9088 162172
rect 182180 162120 182232 162172
rect 118884 160692 118936 160744
rect 580448 160692 580500 160744
rect 73804 160080 73856 160132
rect 76564 160012 76616 160064
rect 64144 159332 64196 159384
rect 66168 159332 66220 159384
rect 82820 159060 82872 159112
rect 86592 159060 86644 159112
rect 175188 158856 175240 158908
rect 177304 158856 177356 158908
rect 88984 158652 89036 158704
rect 96528 158652 96580 158704
rect 154488 157972 154540 158024
rect 165620 157972 165672 158024
rect 378876 157360 378928 157412
rect 380256 157360 380308 157412
rect 71044 154504 71096 154556
rect 74172 154504 74224 154556
rect 165620 154504 165672 154556
rect 168380 154504 168432 154556
rect 377404 154096 377456 154148
rect 378876 154096 378928 154148
rect 96528 153824 96580 153876
rect 109684 153824 109736 153876
rect 118976 153824 119028 153876
rect 580632 153824 580684 153876
rect 86592 153144 86644 153196
rect 89628 153144 89680 153196
rect 180156 151784 180208 151836
rect 580172 151784 580224 151836
rect 66260 151444 66312 151496
rect 68376 151444 68428 151496
rect 3240 149676 3292 149728
rect 22836 149676 22888 149728
rect 118516 148316 118568 148368
rect 166448 148316 166500 148368
rect 86224 147908 86276 147960
rect 88984 147908 89036 147960
rect 76564 147568 76616 147620
rect 79968 147568 80020 147620
rect 171784 146956 171836 147008
rect 172520 146956 172572 147008
rect 89628 146888 89680 146940
rect 106004 146888 106056 146940
rect 141700 146208 141752 146260
rect 142436 146208 142488 146260
rect 139492 146072 139544 146124
rect 142252 146072 142304 146124
rect 74172 145528 74224 145580
rect 78680 145528 78732 145580
rect 177304 144848 177356 144900
rect 180248 144848 180300 144900
rect 106004 144576 106056 144628
rect 109776 144576 109828 144628
rect 33784 144440 33836 144492
rect 182272 144440 182324 144492
rect 10416 144372 10468 144424
rect 182548 144372 182600 144424
rect 6184 144304 6236 144356
rect 182456 144304 182508 144356
rect 118056 144236 118108 144288
rect 398104 144236 398156 144288
rect 119252 144168 119304 144220
rect 477500 144168 477552 144220
rect 79968 143556 80020 143608
rect 78680 143488 78732 143540
rect 82084 143488 82136 143540
rect 84200 143488 84252 143540
rect 146484 143488 146536 143540
rect 148048 143488 148100 143540
rect 153476 143488 153528 143540
rect 158996 143488 159048 143540
rect 167644 143488 167696 143540
rect 169944 143488 169996 143540
rect 172520 143488 172572 143540
rect 176476 143488 176528 143540
rect 137744 143420 137796 143472
rect 139584 143420 139636 143472
rect 152464 143420 152516 143472
rect 157432 143420 157484 143472
rect 163596 143148 163648 143200
rect 174636 143148 174688 143200
rect 150532 143080 150584 143132
rect 154580 143080 154632 143132
rect 164516 143080 164568 143132
rect 176200 143080 176252 143132
rect 144460 143012 144512 143064
rect 160560 143012 160612 143064
rect 163504 143012 163556 143064
rect 178040 143012 178092 143064
rect 142528 142944 142580 142996
rect 173072 142944 173124 142996
rect 118148 142876 118200 142928
rect 398196 142876 398248 142928
rect 118240 142808 118292 142860
rect 418896 142808 418948 142860
rect 149520 142196 149572 142248
rect 152740 142128 152792 142180
rect 157340 142128 157392 142180
rect 163688 142128 163740 142180
rect 40040 141720 40092 141772
rect 181168 141720 181220 141772
rect 4896 141652 4948 141704
rect 182824 141652 182876 141704
rect 119344 141584 119396 141636
rect 412640 141584 412692 141636
rect 120724 141516 120776 141568
rect 542360 141516 542412 141568
rect 119160 141448 119212 141500
rect 580816 141448 580868 141500
rect 119068 141380 119120 141432
rect 580908 141380 580960 141432
rect 176476 141312 176528 141364
rect 181076 141312 181128 141364
rect 367376 140768 367428 140820
rect 370504 140768 370556 140820
rect 109684 140156 109736 140208
rect 180340 140156 180392 140208
rect 10324 140088 10376 140140
rect 182732 140088 182784 140140
rect 4804 140020 4856 140072
rect 182640 140020 182692 140072
rect 375012 139816 375064 139868
rect 377404 139816 377456 139868
rect 98644 139612 98696 139664
rect 100852 139612 100904 139664
rect 62764 139476 62816 139528
rect 182364 139476 182416 139528
rect 118332 139408 118384 139460
rect 580172 139408 580224 139460
rect 3884 138660 3936 138712
rect 25504 138660 25556 138712
rect 88984 138660 89036 138712
rect 97264 138660 97316 138712
rect 373264 137368 373316 137420
rect 375012 137368 375064 137420
rect 84200 137300 84252 137352
rect 87604 137300 87656 137352
rect 3240 136688 3292 136740
rect 116584 136688 116636 136740
rect 3884 136620 3936 136672
rect 117320 136620 117372 136672
rect 365536 136212 365588 136264
rect 367376 136212 367428 136264
rect 4068 135260 4120 135312
rect 117320 135260 117372 135312
rect 100852 135192 100904 135244
rect 102876 135192 102928 135244
rect 182364 134444 182416 134496
rect 182640 134444 182692 134496
rect 3240 133900 3292 133952
rect 117320 133900 117372 133952
rect 362224 133900 362276 133952
rect 365536 133900 365588 133952
rect 25504 132404 25556 132456
rect 117320 132404 117372 132456
rect 68284 132132 68336 132184
rect 69020 132132 69072 132184
rect 109776 131724 109828 131776
rect 117964 131724 118016 131776
rect 7564 131044 7616 131096
rect 117320 131044 117372 131096
rect 69020 130976 69072 131028
rect 74908 130976 74960 131028
rect 87604 129752 87656 129804
rect 90364 129752 90416 129804
rect 22744 129684 22796 129736
rect 117320 129684 117372 129736
rect 369860 129684 369912 129736
rect 373264 129752 373316 129804
rect 102876 129616 102928 129668
rect 104164 129616 104216 129668
rect 68376 129004 68428 129056
rect 69664 129004 69716 129056
rect 74908 129004 74960 129056
rect 84844 129004 84896 129056
rect 22836 128256 22888 128308
rect 117320 128256 117372 128308
rect 180340 128256 180392 128308
rect 182180 128256 182232 128308
rect 24124 126896 24176 126948
rect 117320 126896 117372 126948
rect 184204 125604 184256 125656
rect 580080 125604 580132 125656
rect 8944 125536 8996 125588
rect 117320 125536 117372 125588
rect 367744 125128 367796 125180
rect 369768 125128 369820 125180
rect 4988 124108 5040 124160
rect 117320 124108 117372 124160
rect 97264 124040 97316 124092
rect 100116 124040 100168 124092
rect 82084 123428 82136 123480
rect 90456 123428 90508 123480
rect 43444 122748 43496 122800
rect 117320 122748 117372 122800
rect 100024 122068 100076 122120
rect 110420 122068 110472 122120
rect 37924 121388 37976 121440
rect 117320 121388 117372 121440
rect 69664 120844 69716 120896
rect 71688 120844 71740 120896
rect 19984 120028 20036 120080
rect 117320 120028 117372 120080
rect 180248 120028 180300 120080
rect 182272 120028 182324 120080
rect 110420 119960 110472 120012
rect 114468 119960 114520 120012
rect 71688 119892 71740 119944
rect 73160 119892 73212 119944
rect 355968 119348 356020 119400
rect 366364 119348 366416 119400
rect 15844 118600 15896 118652
rect 117320 118600 117372 118652
rect 104164 118532 104216 118584
rect 108304 118532 108356 118584
rect 23480 117240 23532 117292
rect 117320 117240 117372 117292
rect 352564 116832 352616 116884
rect 355968 116832 356020 116884
rect 73160 114860 73212 114912
rect 74908 114860 74960 114912
rect 114468 114452 114520 114504
rect 117320 114452 117372 114504
rect 100116 113772 100168 113824
rect 111800 113772 111852 113824
rect 84844 113092 84896 113144
rect 117320 113092 117372 113144
rect 90364 112140 90416 112192
rect 91836 112140 91888 112192
rect 74908 111800 74960 111852
rect 3148 111732 3200 111784
rect 62764 111732 62816 111784
rect 180248 111800 180300 111852
rect 580172 111800 580224 111852
rect 117320 111732 117372 111784
rect 183284 111732 183336 111784
rect 362224 111732 362276 111784
rect 91836 111052 91888 111104
rect 97908 111052 97960 111104
rect 90456 110508 90508 110560
rect 93124 110508 93176 110560
rect 349528 110440 349580 110492
rect 352564 110440 352616 110492
rect 97908 110372 97960 110424
rect 117320 110372 117372 110424
rect 183468 110372 183520 110424
rect 367744 110372 367796 110424
rect 182272 108944 182324 108996
rect 410524 108944 410576 108996
rect 108304 108264 108356 108316
rect 109776 108264 109828 108316
rect 111800 106904 111852 106956
rect 119436 106904 119488 106956
rect 183468 106224 183520 106276
rect 409144 106224 409196 106276
rect 346400 105544 346452 105596
rect 349528 105544 349580 105596
rect 109776 104796 109828 104848
rect 111156 104796 111208 104848
rect 183468 104796 183520 104848
rect 407764 104796 407816 104848
rect 183468 103436 183520 103488
rect 406384 103436 406436 103488
rect 343640 102144 343692 102196
rect 346400 102144 346452 102196
rect 182916 102076 182968 102128
rect 405004 102076 405056 102128
rect 93124 101396 93176 101448
rect 102140 101396 102192 101448
rect 182916 100648 182968 100700
rect 403624 100648 403676 100700
rect 117964 99356 118016 99408
rect 120908 99356 120960 99408
rect 180340 99356 180392 99408
rect 580172 99356 580224 99408
rect 102140 99288 102192 99340
rect 105544 99288 105596 99340
rect 183100 99288 183152 99340
rect 400864 99288 400916 99340
rect 111156 97928 111208 97980
rect 112444 97928 112496 97980
rect 183468 97928 183520 97980
rect 399484 97928 399536 97980
rect 183192 96568 183244 96620
rect 421564 96568 421616 96620
rect 183284 95140 183336 95192
rect 418804 95140 418856 95192
rect 339224 94936 339276 94988
rect 343640 94936 343692 94988
rect 183284 93780 183336 93832
rect 417424 93780 417476 93832
rect 183468 92420 183520 92472
rect 414664 92420 414716 92472
rect 112444 92216 112496 92268
rect 113916 92216 113968 92268
rect 329104 91740 329156 91792
rect 339224 91740 339276 91792
rect 182180 89632 182232 89684
rect 188344 89632 188396 89684
rect 180984 88272 181036 88324
rect 226984 88272 227036 88324
rect 113916 86912 113968 86964
rect 116676 86912 116728 86964
rect 182180 86708 182232 86760
rect 184204 86708 184256 86760
rect 105544 86232 105596 86284
rect 120724 86232 120776 86284
rect 182640 85552 182692 85604
rect 580172 85552 580224 85604
rect 3148 84804 3200 84856
rect 3332 84804 3384 84856
rect 3424 84804 3476 84856
rect 3608 84804 3660 84856
rect 3976 84736 4028 84788
rect 3608 84668 3660 84720
rect 3792 84668 3844 84720
rect 3792 84532 3844 84584
rect 3976 84192 4028 84244
rect 120448 84192 120500 84244
rect 116676 82356 116728 82408
rect 119988 82356 120040 82408
rect 182456 81404 182508 81456
rect 555424 81404 555476 81456
rect 119436 80724 119488 80776
rect 5264 80656 5316 80708
rect 119988 80044 120040 80096
rect 124128 79976 124180 80028
rect 125830 79908 125882 79960
rect 125922 79908 125974 79960
rect 126014 79908 126066 79960
rect 126382 79908 126434 79960
rect 126566 79908 126618 79960
rect 125876 79772 125928 79824
rect 125692 79704 125744 79756
rect 5172 79568 5224 79620
rect 125968 79568 126020 79620
rect 126152 79568 126204 79620
rect 126474 79840 126526 79892
rect 126934 79840 126986 79892
rect 127118 79840 127170 79892
rect 126612 79704 126664 79756
rect 127302 79840 127354 79892
rect 127164 79704 127216 79756
rect 127256 79704 127308 79756
rect 127762 79908 127814 79960
rect 128038 79908 128090 79960
rect 127854 79840 127906 79892
rect 127946 79840 127998 79892
rect 128222 79908 128274 79960
rect 128866 79908 128918 79960
rect 128958 79908 129010 79960
rect 128084 79772 128136 79824
rect 127900 79704 127952 79756
rect 127992 79704 128044 79756
rect 128406 79840 128458 79892
rect 128590 79840 128642 79892
rect 128268 79636 128320 79688
rect 128682 79772 128734 79824
rect 128820 79704 128872 79756
rect 128728 79636 128780 79688
rect 128360 79568 128412 79620
rect 128452 79568 128504 79620
rect 128636 79568 128688 79620
rect 129602 79840 129654 79892
rect 130062 79908 130114 79960
rect 130338 79908 130390 79960
rect 129878 79772 129930 79824
rect 130246 79840 130298 79892
rect 130430 79840 130482 79892
rect 130154 79772 130206 79824
rect 130016 79704 130068 79756
rect 130292 79704 130344 79756
rect 130384 79704 130436 79756
rect 130614 79908 130666 79960
rect 130706 79908 130758 79960
rect 130798 79908 130850 79960
rect 130982 79908 131034 79960
rect 129832 79636 129884 79688
rect 130108 79636 130160 79688
rect 130476 79636 130528 79688
rect 130660 79636 130712 79688
rect 129556 79568 129608 79620
rect 129740 79568 129792 79620
rect 130752 79568 130804 79620
rect 126428 79500 126480 79552
rect 126888 79500 126940 79552
rect 127348 79500 127400 79552
rect 116584 79432 116636 79484
rect 127900 79432 127952 79484
rect 130936 79500 130988 79552
rect 3332 79296 3384 79348
rect 127440 79364 127492 79416
rect 127624 79296 127676 79348
rect 127900 79296 127952 79348
rect 129464 79432 129516 79484
rect 131350 79908 131402 79960
rect 131534 79908 131586 79960
rect 132638 79908 132690 79960
rect 133006 79908 133058 79960
rect 131166 79840 131218 79892
rect 131258 79840 131310 79892
rect 131350 79772 131402 79824
rect 131304 79568 131356 79620
rect 131994 79840 132046 79892
rect 131810 79772 131862 79824
rect 132178 79772 132230 79824
rect 132454 79772 132506 79824
rect 131948 79704 132000 79756
rect 131856 79636 131908 79688
rect 132132 79568 132184 79620
rect 132684 79704 132736 79756
rect 132960 79704 133012 79756
rect 132592 79636 132644 79688
rect 133466 79908 133518 79960
rect 133834 79908 133886 79960
rect 134110 79908 134162 79960
rect 134202 79908 134254 79960
rect 133282 79840 133334 79892
rect 133190 79772 133242 79824
rect 131212 79500 131264 79552
rect 131488 79500 131540 79552
rect 132408 79500 132460 79552
rect 133236 79568 133288 79620
rect 133052 79500 133104 79552
rect 133558 79772 133610 79824
rect 133650 79772 133702 79824
rect 133926 79840 133978 79892
rect 133788 79704 133840 79756
rect 133880 79704 133932 79756
rect 133972 79704 134024 79756
rect 134386 79840 134438 79892
rect 134248 79772 134300 79824
rect 133604 79636 133656 79688
rect 134340 79568 134392 79620
rect 133420 79500 133472 79552
rect 134064 79500 134116 79552
rect 134570 79908 134622 79960
rect 134846 79908 134898 79960
rect 135030 79908 135082 79960
rect 135122 79908 135174 79960
rect 135582 79908 135634 79960
rect 135674 79908 135726 79960
rect 136042 79908 136094 79960
rect 136134 79908 136186 79960
rect 136226 79908 136278 79960
rect 136318 79908 136370 79960
rect 136502 79908 136554 79960
rect 134662 79840 134714 79892
rect 134754 79840 134806 79892
rect 134616 79704 134668 79756
rect 134708 79704 134760 79756
rect 134800 79704 134852 79756
rect 134984 79636 135036 79688
rect 135076 79636 135128 79688
rect 135536 79636 135588 79688
rect 133236 79432 133288 79484
rect 135950 79840 136002 79892
rect 135766 79772 135818 79824
rect 135720 79636 135772 79688
rect 135996 79704 136048 79756
rect 136088 79704 136140 79756
rect 135904 79568 135956 79620
rect 135812 79500 135864 79552
rect 136456 79772 136508 79824
rect 136778 79908 136830 79960
rect 137146 79908 137198 79960
rect 137238 79908 137290 79960
rect 136870 79840 136922 79892
rect 136962 79772 137014 79824
rect 137100 79772 137152 79824
rect 136916 79636 136968 79688
rect 137008 79636 137060 79688
rect 137330 79840 137382 79892
rect 138066 79908 138118 79960
rect 138158 79908 138210 79960
rect 138434 79908 138486 79960
rect 138710 79908 138762 79960
rect 138802 79908 138854 79960
rect 138894 79908 138946 79960
rect 137606 79840 137658 79892
rect 136364 79568 136416 79620
rect 136640 79568 136692 79620
rect 137376 79568 137428 79620
rect 137468 79568 137520 79620
rect 137974 79840 138026 79892
rect 137882 79772 137934 79824
rect 138342 79840 138394 79892
rect 138388 79704 138440 79756
rect 138296 79568 138348 79620
rect 137928 79500 137980 79552
rect 138020 79500 138072 79552
rect 136732 79432 136784 79484
rect 137284 79432 137336 79484
rect 137652 79432 137704 79484
rect 137836 79432 137888 79484
rect 138112 79432 138164 79484
rect 138572 79636 138624 79688
rect 138848 79568 138900 79620
rect 138664 79500 138716 79552
rect 139170 79908 139222 79960
rect 139262 79908 139314 79960
rect 139446 79840 139498 79892
rect 139216 79772 139268 79824
rect 139032 79636 139084 79688
rect 139124 79636 139176 79688
rect 139400 79568 139452 79620
rect 139814 79908 139866 79960
rect 140182 79908 140234 79960
rect 140274 79908 140326 79960
rect 140366 79908 140418 79960
rect 140826 79908 140878 79960
rect 140918 79908 140970 79960
rect 141378 79908 141430 79960
rect 141470 79908 141522 79960
rect 141562 79908 141614 79960
rect 141930 79908 141982 79960
rect 139906 79840 139958 79892
rect 139998 79772 140050 79824
rect 139860 79704 139912 79756
rect 139952 79636 140004 79688
rect 140642 79840 140694 79892
rect 140412 79636 140464 79688
rect 139584 79500 139636 79552
rect 140320 79568 140372 79620
rect 140688 79636 140740 79688
rect 141194 79840 141246 79892
rect 141102 79772 141154 79824
rect 140872 79636 140924 79688
rect 141056 79636 141108 79688
rect 140780 79568 140832 79620
rect 141332 79636 141384 79688
rect 141746 79840 141798 79892
rect 141792 79704 141844 79756
rect 141608 79636 141660 79688
rect 142022 79840 142074 79892
rect 141516 79568 141568 79620
rect 141884 79568 141936 79620
rect 140320 79432 140372 79484
rect 131120 79364 131172 79416
rect 132868 79364 132920 79416
rect 133144 79364 133196 79416
rect 134892 79364 134944 79416
rect 140504 79364 140556 79416
rect 131120 79228 131172 79280
rect 141332 79296 141384 79348
rect 141700 79296 141752 79348
rect 142206 79908 142258 79960
rect 142298 79908 142350 79960
rect 142482 79908 142534 79960
rect 143218 79908 143270 79960
rect 143310 79908 143362 79960
rect 143494 79908 143546 79960
rect 143586 79908 143638 79960
rect 144230 79908 144282 79960
rect 144506 79908 144558 79960
rect 144598 79908 144650 79960
rect 142252 79704 142304 79756
rect 142666 79840 142718 79892
rect 142850 79840 142902 79892
rect 142436 79636 142488 79688
rect 142942 79772 142994 79824
rect 142896 79636 142948 79688
rect 142804 79568 142856 79620
rect 143356 79772 143408 79824
rect 143264 79636 143316 79688
rect 143448 79636 143500 79688
rect 143678 79840 143730 79892
rect 143540 79568 143592 79620
rect 142988 79500 143040 79552
rect 143954 79772 144006 79824
rect 143632 79432 143684 79484
rect 142160 79296 142212 79348
rect 143908 79636 143960 79688
rect 144414 79840 144466 79892
rect 144460 79636 144512 79688
rect 144552 79636 144604 79688
rect 144276 79568 144328 79620
rect 144092 79500 144144 79552
rect 143816 79432 143868 79484
rect 145334 79908 145386 79960
rect 145610 79908 145662 79960
rect 144966 79840 145018 79892
rect 145150 79840 145202 79892
rect 144920 79704 144972 79756
rect 145104 79636 145156 79688
rect 144736 79500 144788 79552
rect 145288 79500 145340 79552
rect 146254 79908 146306 79960
rect 146438 79908 146490 79960
rect 146622 79908 146674 79960
rect 146530 79840 146582 79892
rect 146392 79704 146444 79756
rect 146484 79704 146536 79756
rect 146300 79636 146352 79688
rect 146208 79568 146260 79620
rect 146806 79840 146858 79892
rect 146668 79500 146720 79552
rect 146208 79432 146260 79484
rect 146392 79432 146444 79484
rect 147266 79908 147318 79960
rect 147450 79908 147502 79960
rect 147542 79908 147594 79960
rect 147634 79908 147686 79960
rect 147726 79908 147778 79960
rect 147910 79908 147962 79960
rect 148002 79908 148054 79960
rect 148094 79908 148146 79960
rect 148370 79908 148422 79960
rect 148462 79908 148514 79960
rect 148738 79908 148790 79960
rect 149106 79908 149158 79960
rect 146990 79840 147042 79892
rect 147036 79568 147088 79620
rect 147358 79840 147410 79892
rect 147312 79704 147364 79756
rect 147404 79704 147456 79756
rect 147496 79636 147548 79688
rect 146944 79500 146996 79552
rect 147128 79432 147180 79484
rect 147588 79568 147640 79620
rect 147864 79704 147916 79756
rect 147956 79704 148008 79756
rect 148048 79704 148100 79756
rect 148324 79568 148376 79620
rect 149474 79908 149526 79960
rect 149658 79908 149710 79960
rect 149750 79908 149802 79960
rect 149290 79840 149342 79892
rect 149336 79636 149388 79688
rect 149704 79772 149756 79824
rect 149612 79636 149664 79688
rect 148600 79568 148652 79620
rect 148784 79568 148836 79620
rect 149428 79568 149480 79620
rect 150026 79908 150078 79960
rect 150854 79908 150906 79960
rect 151038 79908 151090 79960
rect 149934 79840 149986 79892
rect 150394 79840 150446 79892
rect 150348 79636 150400 79688
rect 150716 79636 150768 79688
rect 151222 79840 151274 79892
rect 151176 79636 151228 79688
rect 151590 79908 151642 79960
rect 151498 79840 151550 79892
rect 149980 79568 150032 79620
rect 150532 79568 150584 79620
rect 151360 79568 151412 79620
rect 150072 79500 150124 79552
rect 147680 79432 147732 79484
rect 151682 79840 151734 79892
rect 152234 79908 152286 79960
rect 152050 79840 152102 79892
rect 151728 79568 151780 79620
rect 151820 79568 151872 79620
rect 152694 79908 152746 79960
rect 152878 79908 152930 79960
rect 152970 79908 153022 79960
rect 153062 79908 153114 79960
rect 153246 79908 153298 79960
rect 152648 79772 152700 79824
rect 152740 79704 152792 79756
rect 153016 79772 153068 79824
rect 152832 79636 152884 79688
rect 152924 79568 152976 79620
rect 151636 79500 151688 79552
rect 153614 79840 153666 79892
rect 153568 79568 153620 79620
rect 154120 79500 154172 79552
rect 153384 79432 153436 79484
rect 154810 79908 154862 79960
rect 155362 79840 155414 79892
rect 155224 79432 155276 79484
rect 155822 79840 155874 79892
rect 155776 79704 155828 79756
rect 156190 79908 156242 79960
rect 156374 79908 156426 79960
rect 156466 79908 156518 79960
rect 156834 79908 156886 79960
rect 156006 79840 156058 79892
rect 156282 79840 156334 79892
rect 156374 79772 156426 79824
rect 156742 79840 156794 79892
rect 156650 79772 156702 79824
rect 156052 79636 156104 79688
rect 156144 79636 156196 79688
rect 156236 79636 156288 79688
rect 156604 79636 156656 79688
rect 156328 79500 156380 79552
rect 156512 79568 156564 79620
rect 156926 79772 156978 79824
rect 156972 79500 157024 79552
rect 155868 79432 155920 79484
rect 157386 79840 157438 79892
rect 157846 79840 157898 79892
rect 157294 79772 157346 79824
rect 157478 79772 157530 79824
rect 157156 79636 157208 79688
rect 157248 79636 157300 79688
rect 157340 79636 157392 79688
rect 157432 79568 157484 79620
rect 157616 79500 157668 79552
rect 158122 79840 158174 79892
rect 157984 79568 158036 79620
rect 158352 79568 158404 79620
rect 157892 79432 157944 79484
rect 143908 79296 143960 79348
rect 144368 79296 144420 79348
rect 148416 79296 148468 79348
rect 155040 79296 155092 79348
rect 120448 79160 120500 79212
rect 139032 79160 139084 79212
rect 141976 79228 142028 79280
rect 145472 79228 145524 79280
rect 156696 79364 156748 79416
rect 396816 80724 396868 80776
rect 158674 79908 158726 79960
rect 158766 79908 158818 79960
rect 158628 79568 158680 79620
rect 158904 79568 158956 79620
rect 174820 80656 174872 80708
rect 174912 80656 174964 80708
rect 175924 80588 175976 80640
rect 580356 80656 580408 80708
rect 174728 80452 174780 80504
rect 393964 80588 394016 80640
rect 175096 80384 175148 80436
rect 180248 80384 180300 80436
rect 159226 79840 159278 79892
rect 159180 79636 159232 79688
rect 159594 79908 159646 79960
rect 159778 79908 159830 79960
rect 159410 79840 159462 79892
rect 159732 79568 159784 79620
rect 159916 79568 159968 79620
rect 160008 79568 160060 79620
rect 160606 79908 160658 79960
rect 161342 79908 161394 79960
rect 161894 79908 161946 79960
rect 161986 79908 162038 79960
rect 160330 79840 160382 79892
rect 160652 79772 160704 79824
rect 160790 79772 160842 79824
rect 161066 79772 161118 79824
rect 160836 79636 160888 79688
rect 160376 79568 160428 79620
rect 159916 79432 159968 79484
rect 160284 79500 160336 79552
rect 161296 79636 161348 79688
rect 161112 79568 161164 79620
rect 161480 79568 161532 79620
rect 161848 79568 161900 79620
rect 161020 79500 161072 79552
rect 162262 79840 162314 79892
rect 162722 79908 162774 79960
rect 162998 79908 163050 79960
rect 162538 79840 162590 79892
rect 162492 79704 162544 79756
rect 162676 79636 162728 79688
rect 163366 79840 163418 79892
rect 162860 79568 162912 79620
rect 163136 79568 163188 79620
rect 163642 79908 163694 79960
rect 163826 79840 163878 79892
rect 163504 79568 163556 79620
rect 163688 79568 163740 79620
rect 164746 79908 164798 79960
rect 166034 79908 166086 79960
rect 166126 79908 166178 79960
rect 166218 79908 166270 79960
rect 164378 79840 164430 79892
rect 165758 79840 165810 79892
rect 165206 79772 165258 79824
rect 164608 79636 164660 79688
rect 164240 79568 164292 79620
rect 165988 79772 166040 79824
rect 166080 79704 166132 79756
rect 165896 79636 165948 79688
rect 165344 79568 165396 79620
rect 165620 79568 165672 79620
rect 166310 79840 166362 79892
rect 162952 79500 163004 79552
rect 163412 79500 163464 79552
rect 165804 79500 165856 79552
rect 166678 79908 166730 79960
rect 167598 79908 167650 79960
rect 167690 79908 167742 79960
rect 167782 79908 167834 79960
rect 167874 79908 167926 79960
rect 168150 79908 168202 79960
rect 168334 79908 168386 79960
rect 168794 79908 168846 79960
rect 168978 79908 169030 79960
rect 167552 79636 167604 79688
rect 166908 79568 166960 79620
rect 167000 79568 167052 79620
rect 167460 79568 167512 79620
rect 167736 79636 167788 79688
rect 168196 79636 168248 79688
rect 168518 79840 168570 79892
rect 168610 79840 168662 79892
rect 168380 79704 168432 79756
rect 168472 79636 168524 79688
rect 168886 79840 168938 79892
rect 168748 79636 168800 79688
rect 169070 79840 169122 79892
rect 169162 79840 169214 79892
rect 168932 79704 168984 79756
rect 169024 79704 169076 79756
rect 169116 79636 169168 79688
rect 168840 79568 168892 79620
rect 167828 79500 167880 79552
rect 168288 79500 168340 79552
rect 169530 79840 169582 79892
rect 169484 79636 169536 79688
rect 169806 79908 169858 79960
rect 169668 79568 169720 79620
rect 170174 79908 170226 79960
rect 170358 79908 170410 79960
rect 170450 79908 170502 79960
rect 170634 79908 170686 79960
rect 170726 79908 170778 79960
rect 170036 79636 170088 79688
rect 170542 79840 170594 79892
rect 170404 79704 170456 79756
rect 170910 79840 170962 79892
rect 171002 79840 171054 79892
rect 171186 79840 171238 79892
rect 170772 79772 170824 79824
rect 170864 79704 170916 79756
rect 170312 79636 170364 79688
rect 171830 79840 171882 79892
rect 174452 80248 174504 80300
rect 182180 80248 182232 80300
rect 172014 79908 172066 79960
rect 172290 79908 172342 79960
rect 175740 80112 175792 80164
rect 200120 80180 200172 80232
rect 177028 80112 177080 80164
rect 231860 80112 231912 80164
rect 172934 79908 172986 79960
rect 171968 79772 172020 79824
rect 171876 79704 171928 79756
rect 175924 80044 175976 80096
rect 252560 80044 252612 80096
rect 174820 79976 174872 80028
rect 173486 79908 173538 79960
rect 173854 79908 173906 79960
rect 173946 79908 173998 79960
rect 174038 79908 174090 79960
rect 174130 79908 174182 79960
rect 173394 79840 173446 79892
rect 171140 79636 171192 79688
rect 171370 79636 171422 79688
rect 171600 79636 171652 79688
rect 173256 79636 173308 79688
rect 173762 79840 173814 79892
rect 173900 79772 173952 79824
rect 173992 79772 174044 79824
rect 174176 79772 174228 79824
rect 173808 79704 173860 79756
rect 173624 79636 173676 79688
rect 170496 79568 170548 79620
rect 170956 79568 171008 79620
rect 174728 79568 174780 79620
rect 170404 79500 170456 79552
rect 163228 79432 163280 79484
rect 166448 79432 166500 79484
rect 169392 79432 169444 79484
rect 159456 79364 159508 79416
rect 160008 79364 160060 79416
rect 164332 79364 164384 79416
rect 167644 79364 167696 79416
rect 163228 79296 163280 79348
rect 163412 79296 163464 79348
rect 174176 79500 174228 79552
rect 170680 79432 170732 79484
rect 171876 79432 171928 79484
rect 173072 79432 173124 79484
rect 171232 79364 171284 79416
rect 171508 79296 171560 79348
rect 174912 79296 174964 79348
rect 180064 79296 180116 79348
rect 580540 79296 580592 79348
rect 148416 79092 148468 79144
rect 127532 79024 127584 79076
rect 127716 79024 127768 79076
rect 141148 79024 141200 79076
rect 141700 79024 141752 79076
rect 155224 79160 155276 79212
rect 156696 79160 156748 79212
rect 157984 79160 158036 79212
rect 158996 79160 159048 79212
rect 164148 79228 164200 79280
rect 178132 79228 178184 79280
rect 173900 79160 173952 79212
rect 164332 79092 164384 79144
rect 195980 79092 196032 79144
rect 164792 79024 164844 79076
rect 165160 79024 165212 79076
rect 249800 79024 249852 79076
rect 5080 78820 5132 78872
rect 140504 78888 140556 78940
rect 144368 78888 144420 78940
rect 164056 78956 164108 79008
rect 213920 78956 213972 79008
rect 147772 78888 147824 78940
rect 267740 78888 267792 78940
rect 127716 78684 127768 78736
rect 129004 78684 129056 78736
rect 155224 78820 155276 78872
rect 161020 78820 161072 78872
rect 173716 78820 173768 78872
rect 176660 78820 176712 78872
rect 329104 78820 329156 78872
rect 166356 78752 166408 78804
rect 444380 78752 444432 78804
rect 168656 78684 168708 78736
rect 554780 78684 554832 78736
rect 126060 78616 126112 78668
rect 126336 78616 126388 78668
rect 128728 78616 128780 78668
rect 129372 78616 129424 78668
rect 137192 78616 137244 78668
rect 137468 78616 137520 78668
rect 145196 78616 145248 78668
rect 158904 78616 158956 78668
rect 163228 78616 163280 78668
rect 171692 78616 171744 78668
rect 171784 78616 171836 78668
rect 178592 78616 178644 78668
rect 139216 78548 139268 78600
rect 140504 78548 140556 78600
rect 144920 78548 144972 78600
rect 165160 78548 165212 78600
rect 166448 78548 166500 78600
rect 171508 78548 171560 78600
rect 172336 78548 172388 78600
rect 176568 78548 176620 78600
rect 126336 78480 126388 78532
rect 130568 78480 130620 78532
rect 140688 78480 140740 78532
rect 164332 78480 164384 78532
rect 170128 78480 170180 78532
rect 170588 78480 170640 78532
rect 141056 78412 141108 78464
rect 155224 78412 155276 78464
rect 161204 78412 161256 78464
rect 146760 78344 146812 78396
rect 164056 78344 164108 78396
rect 125048 78208 125100 78260
rect 132408 78276 132460 78328
rect 154304 78276 154356 78328
rect 162400 78276 162452 78328
rect 164792 78412 164844 78464
rect 173808 78412 173860 78464
rect 165712 78344 165764 78396
rect 171876 78344 171928 78396
rect 173992 78344 174044 78396
rect 174544 78344 174596 78396
rect 247684 78276 247736 78328
rect 133512 78208 133564 78260
rect 136916 78208 136968 78260
rect 146392 78208 146444 78260
rect 147036 78208 147088 78260
rect 161664 78208 161716 78260
rect 253204 78208 253256 78260
rect 89720 78140 89772 78192
rect 132500 78140 132552 78192
rect 148140 78140 148192 78192
rect 148324 78140 148376 78192
rect 153108 78140 153160 78192
rect 161020 78140 161072 78192
rect 171600 78140 171652 78192
rect 322204 78140 322256 78192
rect 46204 78072 46256 78124
rect 126704 78072 126756 78124
rect 136824 78072 136876 78124
rect 137468 78072 137520 78124
rect 140872 78072 140924 78124
rect 150164 78072 150216 78124
rect 158904 78072 158956 78124
rect 159548 78072 159600 78124
rect 162492 78072 162544 78124
rect 471980 78072 472032 78124
rect 57244 78004 57296 78056
rect 127624 78004 127676 78056
rect 149244 78004 149296 78056
rect 149796 78004 149848 78056
rect 163964 78004 164016 78056
rect 480260 78004 480312 78056
rect 22744 77936 22796 77988
rect 125692 77936 125744 77988
rect 134524 77936 134576 77988
rect 135260 77936 135312 77988
rect 147864 77936 147916 77988
rect 148140 77936 148192 77988
rect 150072 77936 150124 77988
rect 157064 77936 157116 77988
rect 167644 77936 167696 77988
rect 498200 77936 498252 77988
rect 125324 77868 125376 77920
rect 133420 77868 133472 77920
rect 152464 77868 152516 77920
rect 159640 77868 159692 77920
rect 161296 77868 161348 77920
rect 180064 77868 180116 77920
rect 125232 77800 125284 77852
rect 129464 77800 129516 77852
rect 159180 77800 159232 77852
rect 170220 77800 170272 77852
rect 123576 77732 123628 77784
rect 132776 77732 132828 77784
rect 158628 77732 158680 77784
rect 174544 77732 174596 77784
rect 120816 77664 120868 77716
rect 129004 77664 129056 77716
rect 129096 77664 129148 77716
rect 130292 77664 130344 77716
rect 141700 77664 141752 77716
rect 120632 77596 120684 77648
rect 128452 77596 128504 77648
rect 122288 77528 122340 77580
rect 128084 77528 128136 77580
rect 129004 77528 129056 77580
rect 131396 77528 131448 77580
rect 143448 77528 143500 77580
rect 158352 77664 158404 77716
rect 172428 77664 172480 77716
rect 157524 77596 157576 77648
rect 171416 77596 171468 77648
rect 174452 77596 174504 77648
rect 122104 77460 122156 77512
rect 125876 77460 125928 77512
rect 127624 77392 127676 77444
rect 129188 77392 129240 77444
rect 172060 77528 172112 77580
rect 580724 77528 580776 77580
rect 155224 77460 155276 77512
rect 164148 77460 164200 77512
rect 164516 77460 164568 77512
rect 166448 77460 166500 77512
rect 170220 77460 170272 77512
rect 175924 77460 175976 77512
rect 177028 77392 177080 77444
rect 124956 77324 125008 77376
rect 126520 77324 126572 77376
rect 129832 77324 129884 77376
rect 134892 77324 134944 77376
rect 139400 77324 139452 77376
rect 155224 77324 155276 77376
rect 120724 77256 120776 77308
rect 125140 77256 125192 77308
rect 126980 77256 127032 77308
rect 132500 77256 132552 77308
rect 133880 77256 133932 77308
rect 153568 77256 153620 77308
rect 164792 77324 164844 77376
rect 168288 77324 168340 77376
rect 169392 77324 169444 77376
rect 156328 77256 156380 77308
rect 165160 77256 165212 77308
rect 167092 77256 167144 77308
rect 173164 77256 173216 77308
rect 153200 77188 153252 77240
rect 153476 77188 153528 77240
rect 156144 77188 156196 77240
rect 156972 77188 157024 77240
rect 162216 77188 162268 77240
rect 167920 77188 167972 77240
rect 168288 77188 168340 77240
rect 168840 77188 168892 77240
rect 175740 77188 175792 77240
rect 527180 77188 527232 77240
rect 172612 77120 172664 77172
rect 145104 77052 145156 77104
rect 147404 77052 147456 77104
rect 150164 77052 150216 77104
rect 197360 77052 197412 77104
rect 124864 76984 124916 77036
rect 134800 76984 134852 77036
rect 152188 76984 152240 77036
rect 152464 76984 152516 77036
rect 153476 76984 153528 77036
rect 154120 76984 154172 77036
rect 157432 76984 157484 77036
rect 158628 76984 158680 77036
rect 162768 76984 162820 77036
rect 211804 76984 211856 77036
rect 133420 76916 133472 76968
rect 135536 76916 135588 76968
rect 143172 76916 143224 76968
rect 226340 76916 226392 76968
rect 122840 76848 122892 76900
rect 135076 76848 135128 76900
rect 144276 76848 144328 76900
rect 240140 76848 240192 76900
rect 102140 76780 102192 76832
rect 86960 76712 87012 76764
rect 123484 76712 123536 76764
rect 131396 76780 131448 76832
rect 131764 76780 131816 76832
rect 134248 76780 134300 76832
rect 134616 76780 134668 76832
rect 145932 76780 145984 76832
rect 260840 76780 260892 76832
rect 133236 76712 133288 76764
rect 133880 76712 133932 76764
rect 135904 76712 135956 76764
rect 140228 76712 140280 76764
rect 140412 76712 140464 76764
rect 147956 76712 148008 76764
rect 288440 76712 288492 76764
rect 69020 76644 69072 76696
rect 130936 76644 130988 76696
rect 133052 76644 133104 76696
rect 133788 76644 133840 76696
rect 148876 76644 148928 76696
rect 296720 76644 296772 76696
rect 44180 76576 44232 76628
rect 128820 76576 128872 76628
rect 134432 76576 134484 76628
rect 135168 76576 135220 76628
rect 135904 76576 135956 76628
rect 136456 76576 136508 76628
rect 136640 76576 136692 76628
rect 136824 76576 136876 76628
rect 137100 76576 137152 76628
rect 137744 76576 137796 76628
rect 150900 76576 150952 76628
rect 151084 76576 151136 76628
rect 152188 76576 152240 76628
rect 152556 76576 152608 76628
rect 153292 76576 153344 76628
rect 153568 76576 153620 76628
rect 154764 76576 154816 76628
rect 155224 76576 155276 76628
rect 156144 76576 156196 76628
rect 156604 76576 156656 76628
rect 156696 76576 156748 76628
rect 157156 76576 157208 76628
rect 157708 76576 157760 76628
rect 157892 76576 157944 76628
rect 159640 76576 159692 76628
rect 324412 76576 324464 76628
rect 30380 76508 30432 76560
rect 127992 76508 128044 76560
rect 124220 76440 124272 76492
rect 123484 76372 123536 76424
rect 132224 76440 132276 76492
rect 151912 76508 151964 76560
rect 152372 76508 152424 76560
rect 158720 76508 158772 76560
rect 159272 76508 159324 76560
rect 160284 76508 160336 76560
rect 160560 76508 160612 76560
rect 161572 76508 161624 76560
rect 162216 76508 162268 76560
rect 163044 76508 163096 76560
rect 163412 76508 163464 76560
rect 164332 76508 164384 76560
rect 164700 76508 164752 76560
rect 165712 76508 165764 76560
rect 166724 76508 166776 76560
rect 167552 76508 167604 76560
rect 167736 76508 167788 76560
rect 167920 76508 167972 76560
rect 454040 76508 454092 76560
rect 172888 76440 172940 76492
rect 120908 76304 120960 76356
rect 172796 76372 172848 76424
rect 131672 76304 131724 76356
rect 132132 76304 132184 76356
rect 151912 76304 151964 76356
rect 152280 76304 152332 76356
rect 154764 76304 154816 76356
rect 155132 76304 155184 76356
rect 163228 76304 163280 76356
rect 163872 76304 163924 76356
rect 164516 76304 164568 76356
rect 165344 76304 165396 76356
rect 168380 76304 168432 76356
rect 168748 76304 168800 76356
rect 169668 76304 169720 76356
rect 172244 76304 172296 76356
rect 144736 76236 144788 76288
rect 145196 76236 145248 76288
rect 154580 76236 154632 76288
rect 162768 76236 162820 76288
rect 163044 76236 163096 76288
rect 163688 76236 163740 76288
rect 164792 76236 164844 76288
rect 172060 76236 172112 76288
rect 135352 76168 135404 76220
rect 135996 76168 136048 76220
rect 143632 76168 143684 76220
rect 148692 76168 148744 76220
rect 152004 76168 152056 76220
rect 152280 76168 152332 76220
rect 154672 76168 154724 76220
rect 155132 76168 155184 76220
rect 160560 76168 160612 76220
rect 160928 76168 160980 76220
rect 142344 76100 142396 76152
rect 145840 76100 145892 76152
rect 150532 76100 150584 76152
rect 158444 76100 158496 76152
rect 160376 76100 160428 76152
rect 160744 76100 160796 76152
rect 142436 76032 142488 76084
rect 142620 76032 142672 76084
rect 143724 76032 143776 76084
rect 144276 76032 144328 76084
rect 145104 76032 145156 76084
rect 145380 76032 145432 76084
rect 137652 75964 137704 76016
rect 144644 75964 144696 76016
rect 144920 75964 144972 76016
rect 145748 75964 145800 76016
rect 139400 75896 139452 75948
rect 139584 75896 139636 75948
rect 139952 75896 140004 75948
rect 140228 75896 140280 75948
rect 141148 75896 141200 75948
rect 141608 75896 141660 75948
rect 143632 75896 143684 75948
rect 144000 75896 144052 75948
rect 145380 75896 145432 75948
rect 145656 75896 145708 75948
rect 157616 75896 157668 75948
rect 158076 75896 158128 75948
rect 161572 75896 161624 75948
rect 162032 75896 162084 75948
rect 169024 75896 169076 75948
rect 170680 75896 170732 75948
rect 125692 75828 125744 75880
rect 126244 75828 126296 75880
rect 140964 75828 141016 75880
rect 141516 75828 141568 75880
rect 142160 75828 142212 75880
rect 142804 75828 142856 75880
rect 143724 75828 143776 75880
rect 144460 75828 144512 75880
rect 147772 75828 147824 75880
rect 148416 75828 148468 75880
rect 155776 75828 155828 75880
rect 156972 75828 157024 75880
rect 169852 75828 169904 75880
rect 170496 75828 170548 75880
rect 139676 75760 139728 75812
rect 140320 75760 140372 75812
rect 142528 75760 142580 75812
rect 142712 75760 142764 75812
rect 144000 75760 144052 75812
rect 144552 75760 144604 75812
rect 148048 75760 148100 75812
rect 148600 75760 148652 75812
rect 126980 75692 127032 75744
rect 134984 75692 135036 75744
rect 135996 75692 136048 75744
rect 136548 75692 136600 75744
rect 139584 75692 139636 75744
rect 140136 75692 140188 75744
rect 158996 75692 159048 75744
rect 164792 75692 164844 75744
rect 130016 75624 130068 75676
rect 130660 75624 130712 75676
rect 132684 75624 132736 75676
rect 133604 75624 133656 75676
rect 158260 75624 158312 75676
rect 122196 75556 122248 75608
rect 130476 75556 130528 75608
rect 159548 75556 159600 75608
rect 121460 75420 121512 75472
rect 126980 75420 127032 75472
rect 396080 75556 396132 75608
rect 164792 75488 164844 75540
rect 431960 75488 432012 75540
rect 438860 75420 438912 75472
rect 51080 75352 51132 75404
rect 128728 75352 128780 75404
rect 138020 75352 138072 75404
rect 138572 75352 138624 75404
rect 146760 75352 146812 75404
rect 147220 75352 147272 75404
rect 161848 75352 161900 75404
rect 467840 75352 467892 75404
rect 107660 75284 107712 75336
rect 132500 75284 132552 75336
rect 157340 75284 157392 75336
rect 157984 75284 158036 75336
rect 167828 75284 167880 75336
rect 490012 75284 490064 75336
rect 42800 75216 42852 75268
rect 6920 75148 6972 75200
rect 125692 75148 125744 75200
rect 125968 75148 126020 75200
rect 126244 75148 126296 75200
rect 127256 75148 127308 75200
rect 128176 75148 128228 75200
rect 128544 75216 128596 75268
rect 129280 75216 129332 75268
rect 130292 75216 130344 75268
rect 131028 75216 131080 75268
rect 138388 75216 138440 75268
rect 138572 75216 138624 75268
rect 140872 75216 140924 75268
rect 141792 75216 141844 75268
rect 146484 75216 146536 75268
rect 146760 75216 146812 75268
rect 149336 75216 149388 75268
rect 149704 75216 149756 75268
rect 166448 75216 166500 75268
rect 499580 75216 499632 75268
rect 128912 75148 128964 75200
rect 131304 75148 131356 75200
rect 132040 75148 132092 75200
rect 146576 75148 146628 75200
rect 146852 75148 146904 75200
rect 160192 75148 160244 75200
rect 160836 75148 160888 75200
rect 169300 75148 169352 75200
rect 564440 75148 564492 75200
rect 125876 75080 125928 75132
rect 126612 75080 126664 75132
rect 127348 75080 127400 75132
rect 128268 75080 128320 75132
rect 128728 75080 128780 75132
rect 129648 75080 129700 75132
rect 138204 75080 138256 75132
rect 138388 75080 138440 75132
rect 142528 75080 142580 75132
rect 142896 75080 142948 75132
rect 170220 75080 170272 75132
rect 170772 75080 170824 75132
rect 125968 75012 126020 75064
rect 126888 75012 126940 75064
rect 128360 75012 128412 75064
rect 133420 75012 133472 75064
rect 125692 74944 125744 74996
rect 126796 74944 126848 74996
rect 128452 74944 128504 74996
rect 129556 74944 129608 74996
rect 138204 74944 138256 74996
rect 138664 74944 138716 74996
rect 164700 74944 164752 74996
rect 164976 74944 165028 74996
rect 146484 74876 146536 74928
rect 147128 74876 147180 74928
rect 155868 74808 155920 74860
rect 159640 74808 159692 74860
rect 146300 74740 146352 74792
rect 147312 74740 147364 74792
rect 161848 74740 161900 74792
rect 162308 74740 162360 74792
rect 147680 74604 147732 74656
rect 148508 74604 148560 74656
rect 154580 74536 154632 74588
rect 155500 74536 155552 74588
rect 168564 74468 168616 74520
rect 173348 74468 173400 74520
rect 153292 74400 153344 74452
rect 153844 74400 153896 74452
rect 150440 74332 150492 74384
rect 156880 74332 156932 74384
rect 145472 74196 145524 74248
rect 209780 74196 209832 74248
rect 145840 74128 145892 74180
rect 216680 74128 216732 74180
rect 118700 74060 118752 74112
rect 134708 74060 134760 74112
rect 142988 74060 143040 74112
rect 223580 74060 223632 74112
rect 93952 73992 94004 74044
rect 133144 73992 133196 74044
rect 145012 73992 145064 74044
rect 145472 73992 145524 74044
rect 147404 73992 147456 74044
rect 251180 73992 251232 74044
rect 64880 73924 64932 73976
rect 129740 73924 129792 73976
rect 142252 73924 142304 73976
rect 143080 73924 143132 73976
rect 157708 73924 157760 73976
rect 158168 73924 158220 73976
rect 158444 73924 158496 73976
rect 318800 73924 318852 73976
rect 27620 73856 27672 73908
rect 127808 73856 127860 73908
rect 135720 73856 135772 73908
rect 136364 73856 136416 73908
rect 145012 73856 145064 73908
rect 146024 73856 146076 73908
rect 152004 73856 152056 73908
rect 152648 73856 152700 73908
rect 153108 73856 153160 73908
rect 354680 73856 354732 73908
rect 26240 73788 26292 73840
rect 127900 73788 127952 73840
rect 143540 73788 143592 73840
rect 144368 73788 144420 73840
rect 164792 73788 164844 73840
rect 165068 73788 165120 73840
rect 165160 73788 165212 73840
rect 375380 73788 375432 73840
rect 150532 73720 150584 73772
rect 151268 73720 151320 73772
rect 158996 73720 159048 73772
rect 159824 73720 159876 73772
rect 161664 73584 161716 73636
rect 162124 73584 162176 73636
rect 137468 73448 137520 73500
rect 138940 73448 138992 73500
rect 155960 73448 156012 73500
rect 156512 73448 156564 73500
rect 154764 73244 154816 73296
rect 155408 73244 155460 73296
rect 137376 73176 137428 73228
rect 142988 73176 143040 73228
rect 177304 73108 177356 73160
rect 580172 73108 580224 73160
rect 158720 72904 158772 72956
rect 158996 72904 159048 72956
rect 148324 72632 148376 72684
rect 291200 72632 291252 72684
rect 149888 72564 149940 72616
rect 311900 72564 311952 72616
rect 152740 72496 152792 72548
rect 340880 72496 340932 72548
rect 153200 72428 153252 72480
rect 357440 72428 357492 72480
rect 165252 72360 165304 72412
rect 171876 72360 171928 72412
rect 168564 72292 168616 72344
rect 169116 72292 169168 72344
rect 167092 72088 167144 72140
rect 168012 72088 168064 72140
rect 3424 71680 3476 71732
rect 179604 71680 179656 71732
rect 78680 71000 78732 71052
rect 131764 71000 131816 71052
rect 138848 71000 138900 71052
rect 152556 71000 152608 71052
rect 157340 71000 157392 71052
rect 284392 71000 284444 71052
rect 138664 70320 138716 70372
rect 142804 70320 142856 70372
rect 141516 70048 141568 70100
rect 209872 70048 209924 70100
rect 155316 69980 155368 70032
rect 382280 69980 382332 70032
rect 156788 69912 156840 69964
rect 390560 69912 390612 69964
rect 171692 69844 171744 69896
rect 426440 69844 426492 69896
rect 164884 69776 164936 69828
rect 505100 69776 505152 69828
rect 166632 69708 166684 69760
rect 518900 69708 518952 69760
rect 170312 69640 170364 69692
rect 568580 69640 568632 69692
rect 170220 68960 170272 69012
rect 171692 68960 171744 69012
rect 140044 68620 140096 68672
rect 184940 68620 184992 68672
rect 142712 68552 142764 68604
rect 218060 68552 218112 68604
rect 156880 68484 156932 68536
rect 320180 68484 320232 68536
rect 153752 68416 153804 68468
rect 362960 68416 363012 68468
rect 159272 68348 159324 68400
rect 427820 68348 427872 68400
rect 169484 68280 169536 68332
rect 564532 68280 564584 68332
rect 139952 67396 140004 67448
rect 189080 67396 189132 67448
rect 147128 67328 147180 67380
rect 270500 67328 270552 67380
rect 149704 67260 149756 67312
rect 306380 67260 306432 67312
rect 161020 67192 161072 67244
rect 347780 67192 347832 67244
rect 152464 67124 152516 67176
rect 340972 67124 341024 67176
rect 159180 67056 159232 67108
rect 437480 67056 437532 67108
rect 162032 66988 162084 67040
rect 462320 66988 462372 67040
rect 167736 66920 167788 66972
rect 539600 66920 539652 66972
rect 167644 66852 167696 66904
rect 543740 66852 543792 66904
rect 137284 66172 137336 66224
rect 140044 66172 140096 66224
rect 138572 66104 138624 66156
rect 141516 66104 141568 66156
rect 141424 65900 141476 65952
rect 202880 65900 202932 65952
rect 141332 65832 141384 65884
rect 207020 65832 207072 65884
rect 142620 65764 142672 65816
rect 220820 65764 220872 65816
rect 145472 65696 145524 65748
rect 251272 65696 251324 65748
rect 145564 65628 145616 65680
rect 256700 65628 256752 65680
rect 153660 65560 153712 65612
rect 358820 65560 358872 65612
rect 102232 65492 102284 65544
rect 125324 65492 125376 65544
rect 155224 65492 155276 65544
rect 376760 65492 376812 65544
rect 144276 64472 144328 64524
rect 234620 64472 234672 64524
rect 144184 64404 144236 64456
rect 238760 64404 238812 64456
rect 148232 64336 148284 64388
rect 292580 64336 292632 64388
rect 152372 64268 152424 64320
rect 338120 64268 338172 64320
rect 162216 64200 162268 64252
rect 368480 64200 368532 64252
rect 169024 64132 169076 64184
rect 561680 64132 561732 64184
rect 147036 63112 147088 63164
rect 274640 63112 274692 63164
rect 149612 63044 149664 63096
rect 309140 63044 309192 63096
rect 155132 62976 155184 63028
rect 374000 62976 374052 63028
rect 157984 62908 158036 62960
rect 408500 62908 408552 62960
rect 163596 62840 163648 62892
rect 488540 62840 488592 62892
rect 168932 62772 168984 62824
rect 557540 62772 557592 62824
rect 139860 61480 139912 61532
rect 185032 61480 185084 61532
rect 157892 61412 157944 61464
rect 412640 61412 412692 61464
rect 166356 61344 166408 61396
rect 525800 61344 525852 61396
rect 118516 60664 118568 60716
rect 580172 60664 580224 60716
rect 137192 59984 137244 60036
rect 138664 59984 138716 60036
rect 159088 59984 159140 60036
rect 433340 59984 433392 60036
rect 156512 58624 156564 58676
rect 401600 58624 401652 58676
rect 163504 57264 163556 57316
rect 481640 57264 481692 57316
rect 164792 57196 164844 57248
rect 507860 57196 507912 57248
rect 95240 53048 95292 53100
rect 125232 53048 125284 53100
rect 182824 46860 182876 46912
rect 580172 46860 580224 46912
rect 139768 46180 139820 46232
rect 180800 46180 180852 46232
rect 3424 45500 3476 45552
rect 174084 45500 174136 45552
rect 135996 44956 136048 45008
rect 142620 44956 142672 45008
rect 70400 44888 70452 44940
rect 130292 44888 130344 44940
rect 34520 44820 34572 44872
rect 127348 44820 127400 44872
rect 138480 44820 138532 44872
rect 147036 44820 147088 44872
rect 171600 43392 171652 43444
rect 411260 43392 411312 43444
rect 19340 42032 19392 42084
rect 125140 42032 125192 42084
rect 162492 42032 162544 42084
rect 390652 42032 390704 42084
rect 172428 40672 172480 40724
rect 418160 40672 418212 40724
rect 120080 40264 120132 40316
rect 123484 40264 123536 40316
rect 172336 39312 172388 39364
rect 404360 39312 404412 39364
rect 172152 37884 172204 37936
rect 397460 37884 397512 37936
rect 88340 36524 88392 36576
rect 125048 36524 125100 36576
rect 145380 35572 145432 35624
rect 259460 35572 259512 35624
rect 146944 35504 146996 35556
rect 276020 35504 276072 35556
rect 148140 35436 148192 35488
rect 287060 35436 287112 35488
rect 148048 35368 148100 35420
rect 293960 35368 294012 35420
rect 149428 35300 149480 35352
rect 305000 35300 305052 35352
rect 149520 35232 149572 35284
rect 307760 35232 307812 35284
rect 159732 35164 159784 35216
rect 382372 35164 382424 35216
rect 139676 34076 139728 34128
rect 187700 34076 187752 34128
rect 141056 34008 141108 34060
rect 198740 34008 198792 34060
rect 141240 33940 141292 33992
rect 201500 33940 201552 33992
rect 141148 33872 141200 33924
rect 205640 33872 205692 33924
rect 144092 33804 144144 33856
rect 234712 33804 234764 33856
rect 146852 33736 146904 33788
rect 269120 33736 269172 33788
rect 171692 33056 171744 33108
rect 580172 33056 580224 33108
rect 3424 32988 3476 33040
rect 181260 32988 181312 33040
rect 156420 32716 156472 32768
rect 391940 32716 391992 32768
rect 160008 32648 160060 32700
rect 434720 32648 434772 32700
rect 161940 32580 161992 32632
rect 463700 32580 463752 32632
rect 163412 32512 163464 32564
rect 481732 32512 481784 32564
rect 167552 32444 167604 32496
rect 539692 32444 539744 32496
rect 170128 32376 170180 32428
rect 574100 32376 574152 32428
rect 144000 31424 144052 31476
rect 242900 31424 242952 31476
rect 146760 31356 146812 31408
rect 267832 31356 267884 31408
rect 147956 31288 148008 31340
rect 289820 31288 289872 31340
rect 154120 31220 154172 31272
rect 332600 31220 332652 31272
rect 153568 31152 153620 31204
rect 357532 31152 357584 31204
rect 156972 31084 157024 31136
rect 389180 31084 389232 31136
rect 166264 31016 166316 31068
rect 524420 31016 524472 31068
rect 140964 30064 141016 30116
rect 204260 30064 204312 30116
rect 140872 29996 140924 30048
rect 208400 29996 208452 30048
rect 143908 29928 143960 29980
rect 233240 29928 233292 29980
rect 143816 29860 143868 29912
rect 236000 29860 236052 29912
rect 145196 29792 145248 29844
rect 253940 29792 253992 29844
rect 145288 29724 145340 29776
rect 258080 29724 258132 29776
rect 166172 29656 166224 29708
rect 521660 29656 521712 29708
rect 167460 29588 167512 29640
rect 542360 29588 542412 29640
rect 148692 28500 148744 28552
rect 190460 28500 190512 28552
rect 139584 28432 139636 28484
rect 186320 28432 186372 28484
rect 140780 28364 140832 28416
rect 201592 28364 201644 28416
rect 146668 28296 146720 28348
rect 271880 28296 271932 28348
rect 147864 28228 147916 28280
rect 285680 28228 285732 28280
rect 322204 28228 322256 28280
rect 581000 28228 581052 28280
rect 140504 27276 140556 27328
rect 176752 27276 176804 27328
rect 139492 27208 139544 27260
rect 179420 27208 179472 27260
rect 139400 27140 139452 27192
rect 183560 27140 183612 27192
rect 146576 27072 146628 27124
rect 276112 27072 276164 27124
rect 149336 27004 149388 27056
rect 310520 27004 310572 27056
rect 152280 26936 152332 26988
rect 339500 26936 339552 26988
rect 164700 26868 164752 26920
rect 506480 26868 506532 26920
rect 142528 25984 142580 26036
rect 222200 25984 222252 26036
rect 146484 25916 146536 25968
rect 278780 25916 278832 25968
rect 149244 25848 149296 25900
rect 307852 25848 307904 25900
rect 152188 25780 152240 25832
rect 346400 25780 346452 25832
rect 166080 25712 166132 25764
rect 517520 25712 517572 25764
rect 170680 25644 170732 25696
rect 558920 25644 558972 25696
rect 168840 25576 168892 25628
rect 563060 25576 563112 25628
rect 170036 25508 170088 25560
rect 572720 25508 572772 25560
rect 142344 24556 142396 24608
rect 215300 24556 215352 24608
rect 142436 24488 142488 24540
rect 218152 24488 218204 24540
rect 147772 24420 147824 24472
rect 292672 24420 292724 24472
rect 155040 24352 155092 24404
rect 374092 24352 374144 24404
rect 167184 24284 167236 24336
rect 467104 24284 467156 24336
rect 167276 24216 167328 24268
rect 535460 24216 535512 24268
rect 167368 24148 167420 24200
rect 538220 24148 538272 24200
rect 168748 24080 168800 24132
rect 552020 24080 552072 24132
rect 149152 23332 149204 23384
rect 303620 23332 303672 23384
rect 3424 23264 3476 23316
rect 173992 23264 174044 23316
rect 153476 23196 153528 23248
rect 360200 23196 360252 23248
rect 154948 23128 155000 23180
rect 379520 23128 379572 23180
rect 164608 23060 164660 23112
rect 498292 23060 498344 23112
rect 164516 22992 164568 23044
rect 509240 22992 509292 23044
rect 165896 22924 165948 22976
rect 516140 22924 516192 22976
rect 165988 22856 166040 22908
rect 520280 22856 520332 22908
rect 74540 22788 74592 22840
rect 129188 22788 129240 22840
rect 168656 22788 168708 22840
rect 556160 22788 556212 22840
rect 118424 22720 118476 22772
rect 580172 22720 580224 22772
rect 152096 21632 152148 21684
rect 343640 21632 343692 21684
rect 160652 21564 160704 21616
rect 447140 21564 447192 21616
rect 161848 21496 161900 21548
rect 473360 21496 473412 21548
rect 163320 21428 163372 21480
rect 484400 21428 484452 21480
rect 124312 21360 124364 21412
rect 134340 21360 134392 21412
rect 164424 21360 164476 21412
rect 506572 21360 506624 21412
rect 145104 20340 145156 20392
rect 255320 20340 255372 20392
rect 145012 20272 145064 20324
rect 262220 20272 262272 20324
rect 146392 20204 146444 20256
rect 273260 20204 273312 20256
rect 247684 20136 247736 20188
rect 456800 20136 456852 20188
rect 138388 20068 138440 20120
rect 162860 20068 162912 20120
rect 253204 20068 253256 20120
rect 465080 20068 465132 20120
rect 85580 20000 85632 20052
rect 131672 20000 131724 20052
rect 160560 20000 160612 20052
rect 455420 20000 455472 20052
rect 45560 19932 45612 19984
rect 120816 19932 120868 19984
rect 161756 19932 161808 19984
rect 465172 19932 465224 19984
rect 160468 18844 160520 18896
rect 448520 18844 448572 18896
rect 160376 18776 160428 18828
rect 451280 18776 451332 18828
rect 117320 18708 117372 18760
rect 134248 18708 134300 18760
rect 168472 18708 168524 18760
rect 553400 18708 553452 18760
rect 31760 18640 31812 18692
rect 122288 18640 122340 18692
rect 168380 18640 168432 18692
rect 556252 18640 556304 18692
rect 4160 18572 4212 18624
rect 126244 18572 126296 18624
rect 168564 18572 168616 18624
rect 560300 18572 560352 18624
rect 157800 17552 157852 17604
rect 415400 17552 415452 17604
rect 157708 17484 157760 17536
rect 419540 17484 419592 17536
rect 171968 17416 172020 17468
rect 440240 17416 440292 17468
rect 160284 17348 160336 17400
rect 448612 17348 448664 17400
rect 163228 17280 163280 17332
rect 492680 17280 492732 17332
rect 167092 17212 167144 17264
rect 545120 17212 545172 17264
rect 154856 16124 154908 16176
rect 378416 16124 378468 16176
rect 156236 16056 156288 16108
rect 395344 16056 395396 16108
rect 156328 15988 156380 16040
rect 398840 15988 398892 16040
rect 174544 15920 174596 15972
rect 425704 15920 425756 15972
rect 14280 15852 14332 15904
rect 124956 15852 125008 15904
rect 167000 15852 167052 15904
rect 541992 15852 542044 15904
rect 143724 14764 143776 14816
rect 241704 14764 241756 14816
rect 154672 14696 154724 14748
rect 381176 14696 381228 14748
rect 154764 14628 154816 14680
rect 384304 14628 384356 14680
rect 154580 14560 154632 14612
rect 385960 14560 386012 14612
rect 114008 14492 114060 14544
rect 134156 14492 134208 14544
rect 158904 14492 158956 14544
rect 436744 14492 436796 14544
rect 39120 14424 39172 14476
rect 120724 14424 120776 14476
rect 164332 14424 164384 14476
rect 502984 14424 503036 14476
rect 151912 13404 151964 13456
rect 345296 13404 345348 13456
rect 152004 13336 152056 13388
rect 349160 13336 349212 13388
rect 153384 13268 153436 13320
rect 365720 13268 365772 13320
rect 157616 13200 157668 13252
rect 417424 13200 417476 13252
rect 158812 13132 158864 13184
rect 429200 13132 429252 13184
rect 160192 13064 160244 13116
rect 453304 13064 453356 13116
rect 143632 11976 143684 12028
rect 237656 11976 237708 12028
rect 150348 11908 150400 11960
rect 313832 11908 313884 11960
rect 157524 11840 157576 11892
rect 414296 11840 414348 11892
rect 157432 11772 157484 11824
rect 415492 11772 415544 11824
rect 165804 11704 165856 11756
rect 523776 11704 523828 11756
rect 176660 11636 176712 11688
rect 177856 11636 177908 11688
rect 184940 11636 184992 11688
rect 186136 11636 186188 11688
rect 201500 11636 201552 11688
rect 202696 11636 202748 11688
rect 234620 11636 234672 11688
rect 235816 11636 235868 11688
rect 106464 10616 106516 10668
rect 133052 10616 133104 10668
rect 99840 10548 99892 10600
rect 132960 10548 133012 10600
rect 147680 10548 147732 10600
rect 295616 10548 295668 10600
rect 81624 10480 81676 10532
rect 131580 10480 131632 10532
rect 153292 10480 153344 10532
rect 364616 10480 364668 10532
rect 35992 10412 36044 10464
rect 127256 10412 127308 10464
rect 156052 10412 156104 10464
rect 394240 10412 394292 10464
rect 28448 10344 28500 10396
rect 127164 10344 127216 10396
rect 156144 10344 156196 10396
rect 398932 10344 398984 10396
rect 11152 10276 11204 10328
rect 126152 10276 126204 10328
rect 163136 10276 163188 10328
rect 486424 10276 486476 10328
rect 67916 9324 67968 9376
rect 130200 9324 130252 9376
rect 64328 9256 64380 9308
rect 126336 9256 126388 9308
rect 144920 9256 144972 9308
rect 260656 9256 260708 9308
rect 63224 9188 63276 9240
rect 130108 9188 130160 9240
rect 146300 9188 146352 9240
rect 278320 9188 278372 9240
rect 60832 9120 60884 9172
rect 129096 9120 129148 9172
rect 151820 9120 151872 9172
rect 343364 9120 343416 9172
rect 53748 9052 53800 9104
rect 128728 9052 128780 9104
rect 161664 9052 161716 9104
rect 471060 9052 471112 9104
rect 50160 8984 50212 9036
rect 127716 8984 127768 9036
rect 163044 8984 163096 9036
rect 492312 8984 492364 9036
rect 572 8916 624 8968
rect 124220 8916 124272 8968
rect 169944 8916 169996 8968
rect 571524 8916 571576 8968
rect 116400 7896 116452 7948
rect 134064 7896 134116 7948
rect 142252 7896 142304 7948
rect 225144 7896 225196 7948
rect 105728 7828 105780 7880
rect 132776 7828 132828 7880
rect 143540 7828 143592 7880
rect 242992 7828 243044 7880
rect 98644 7760 98696 7812
rect 132868 7760 132920 7812
rect 155960 7760 156012 7812
rect 401324 7760 401376 7812
rect 48964 7692 49016 7744
rect 128544 7692 128596 7744
rect 160100 7692 160152 7744
rect 446220 7692 446272 7744
rect 44272 7624 44324 7676
rect 128636 7624 128688 7676
rect 161572 7624 161624 7676
rect 469864 7624 469916 7676
rect 9956 7556 10008 7608
rect 126060 7556 126112 7608
rect 164240 7556 164292 7608
rect 504180 7556 504232 7608
rect 555424 6808 555476 6860
rect 580172 6808 580224 6860
rect 150808 6740 150860 6792
rect 323308 6740 323360 6792
rect 150992 6672 151044 6724
rect 326804 6672 326856 6724
rect 115204 6604 115256 6656
rect 134708 6604 134760 6656
rect 150900 6604 150952 6656
rect 329196 6604 329248 6656
rect 104532 6536 104584 6588
rect 132684 6536 132736 6588
rect 151084 6536 151136 6588
rect 330392 6536 330444 6588
rect 84476 6468 84528 6520
rect 131304 6468 131356 6520
rect 158536 6468 158588 6520
rect 410800 6468 410852 6520
rect 80888 6400 80940 6452
rect 131396 6400 131448 6452
rect 175924 6400 175976 6452
rect 433248 6400 433300 6452
rect 77392 6332 77444 6384
rect 131488 6332 131540 6384
rect 158720 6332 158772 6384
rect 441528 6332 441580 6384
rect 25320 6264 25372 6316
rect 57244 6264 57296 6316
rect 66720 6264 66772 6316
rect 130016 6264 130068 6316
rect 161480 6264 161532 6316
rect 467472 6264 467524 6316
rect 33600 6196 33652 6248
rect 127532 6196 127584 6248
rect 140412 6196 140464 6248
rect 156604 6196 156656 6248
rect 169760 6196 169812 6248
rect 572720 6196 572772 6248
rect 18236 6128 18288 6180
rect 125968 6128 126020 6180
rect 138296 6128 138348 6180
rect 162492 6128 162544 6180
rect 169852 6128 169904 6180
rect 576308 6128 576360 6180
rect 101036 5312 101088 5364
rect 133144 5312 133196 5364
rect 97448 5244 97500 5296
rect 132592 5244 132644 5296
rect 86868 5176 86920 5228
rect 132408 5176 132460 5228
rect 138020 5176 138072 5228
rect 169576 5176 169628 5228
rect 15936 5040 15988 5092
rect 59636 5108 59688 5160
rect 129924 5108 129976 5160
rect 142160 5108 142212 5160
rect 220452 5108 220504 5160
rect 46204 5040 46256 5092
rect 52552 5040 52604 5092
rect 128452 5040 128504 5092
rect 136916 5040 136968 5092
rect 148324 5040 148376 5092
rect 154488 5040 154540 5092
rect 365812 5040 365864 5092
rect 33232 4972 33284 5024
rect 127440 4972 127492 5024
rect 138204 4972 138256 5024
rect 171968 4972 172020 5024
rect 180064 4972 180116 5024
rect 450912 4972 450964 5024
rect 6460 4904 6512 4956
rect 22744 4904 22796 4956
rect 24216 4904 24268 4956
rect 122104 4904 122156 4956
rect 137008 4904 137060 4956
rect 150624 4904 150676 4956
rect 162952 4904 163004 4956
rect 487620 4904 487672 4956
rect 13544 4836 13596 4888
rect 125876 4836 125928 4888
rect 137100 4836 137152 4888
rect 157800 4836 157852 4888
rect 165620 4836 165672 4888
rect 523040 4836 523092 4888
rect 8760 4768 8812 4820
rect 125784 4768 125836 4820
rect 138112 4768 138164 4820
rect 164884 4768 164936 4820
rect 165712 4768 165764 4820
rect 527824 4768 527876 4820
rect 138940 4360 138992 4412
rect 143540 4360 143592 4412
rect 242900 4156 242952 4208
rect 244096 4156 244148 4208
rect 251180 4156 251232 4208
rect 252376 4156 252428 4208
rect 276020 4156 276072 4208
rect 276756 4156 276808 4208
rect 119896 4088 119948 4140
rect 124864 4088 124916 4140
rect 125876 4088 125928 4140
rect 134524 4088 134576 4140
rect 151544 4088 151596 4140
rect 325608 4088 325660 4140
rect 138664 4020 138716 4072
rect 145932 4020 145984 4072
rect 150900 4020 150952 4072
rect 328000 4020 328052 4072
rect 12348 3952 12400 4004
rect 126428 3952 126480 4004
rect 150532 3952 150584 4004
rect 331588 3952 331640 4004
rect 136824 3884 136876 3936
rect 144736 3884 144788 3936
rect 172060 3884 172112 3936
rect 356336 3884 356388 3936
rect 467104 3884 467156 3936
rect 534908 3884 534960 3936
rect 83280 3816 83332 3868
rect 131856 3816 131908 3868
rect 142988 3816 143040 3868
rect 151820 3816 151872 3868
rect 172244 3816 172296 3868
rect 303160 3816 303212 3868
rect 319444 3816 319496 3868
rect 583392 3816 583444 3868
rect 76196 3748 76248 3800
rect 129004 3748 129056 3800
rect 140044 3748 140096 3800
rect 149520 3748 149572 3800
rect 152556 3748 152608 3800
rect 168380 3748 168432 3800
rect 178684 3748 178736 3800
rect 475752 3748 475804 3800
rect 69112 3680 69164 3732
rect 130660 3680 130712 3732
rect 137744 3680 137796 3732
rect 154212 3680 154264 3732
rect 163964 3680 164016 3732
rect 491116 3680 491168 3732
rect 62028 3612 62080 3664
rect 122196 3612 122248 3664
rect 47860 3544 47912 3596
rect 127624 3612 127676 3664
rect 136732 3612 136784 3664
rect 155408 3612 155460 3664
rect 171876 3612 171928 3664
rect 501788 3612 501840 3664
rect 126980 3544 127032 3596
rect 130384 3544 130436 3596
rect 133788 3544 133840 3596
rect 147128 3544 147180 3596
rect 147220 3544 147272 3596
rect 167184 3544 167236 3596
rect 171784 3544 171836 3596
rect 515956 3544 516008 3596
rect 17040 3476 17092 3528
rect 125692 3476 125744 3528
rect 131764 3476 131816 3528
rect 135628 3476 135680 3528
rect 141516 3476 141568 3528
rect 166080 3476 166132 3528
rect 173164 3476 173216 3528
rect 93860 3408 93912 3460
rect 94780 3408 94832 3460
rect 142804 3408 142856 3460
rect 170772 3408 170824 3460
rect 173348 3408 173400 3460
rect 531320 3476 531372 3528
rect 532148 3476 532200 3528
rect 539600 3476 539652 3528
rect 540428 3476 540480 3528
rect 150808 3340 150860 3392
rect 322112 3340 322164 3392
rect 340972 3340 341024 3392
rect 342168 3340 342220 3392
rect 349252 3340 349304 3392
rect 350448 3340 350500 3392
rect 357440 3340 357492 3392
rect 358728 3340 358780 3392
rect 365720 3340 365772 3392
rect 367008 3340 367060 3392
rect 374092 3340 374144 3392
rect 375288 3340 375340 3392
rect 382372 3340 382424 3392
rect 383568 3340 383620 3392
rect 398932 3340 398984 3392
rect 400128 3340 400180 3392
rect 415400 3340 415452 3392
rect 416688 3340 416740 3392
rect 423772 3340 423824 3392
rect 424968 3340 425020 3392
rect 448612 3340 448664 3392
rect 449808 3340 449860 3392
rect 456800 3340 456852 3392
rect 458088 3340 458140 3392
rect 506480 3340 506532 3392
rect 507308 3340 507360 3392
rect 533712 3408 533764 3460
rect 537208 3340 537260 3392
rect 135720 3272 135772 3324
rect 138848 3272 138900 3324
rect 144460 3272 144512 3324
rect 153016 3272 153068 3324
rect 173256 3272 173308 3324
rect 212172 3272 212224 3324
rect 211804 3204 211856 3256
rect 362316 3272 362368 3324
rect 307760 3204 307812 3256
rect 309048 3204 309100 3256
rect 316040 3204 316092 3256
rect 317328 3204 317380 3256
rect 135536 3136 135588 3188
rect 140044 3136 140096 3188
rect 132960 3068 133012 3120
rect 135444 3068 135496 3120
rect 135812 3068 135864 3120
rect 137652 3068 137704 3120
rect 135904 3000 135956 3052
rect 141240 3000 141292 3052
rect 390560 1232 390612 1284
rect 391848 1232 391900 1284
rect 30104 1096 30156 1148
rect 33232 1096 33284 1148
<< metal2 >>
rect 6932 703582 7972 703610
rect 2778 684312 2834 684321
rect 2778 684247 2834 684256
rect 2792 683738 2820 684247
rect 2780 683732 2832 683738
rect 2780 683674 2832 683680
rect 4804 683732 4856 683738
rect 4804 683674 4856 683680
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 2780 632120 2832 632126
rect 2778 632088 2780 632097
rect 2832 632088 2834 632097
rect 2778 632023 2834 632032
rect 3054 566944 3110 566953
rect 3054 566879 3110 566888
rect 3068 565894 3096 566879
rect 3056 565888 3108 565894
rect 3056 565830 3108 565836
rect 3330 514856 3386 514865
rect 3330 514791 3332 514800
rect 3384 514791 3386 514800
rect 3332 514762 3384 514768
rect 2778 462632 2834 462641
rect 2778 462567 2780 462576
rect 2832 462567 2834 462576
rect 2780 462538 2832 462544
rect 3146 423600 3202 423609
rect 3146 423535 3202 423544
rect 3160 422958 3188 423535
rect 3148 422952 3200 422958
rect 3148 422894 3200 422900
rect 3330 410544 3386 410553
rect 3330 410479 3386 410488
rect 3344 409970 3372 410479
rect 3332 409964 3384 409970
rect 3332 409906 3384 409912
rect 3330 371376 3386 371385
rect 3330 371311 3386 371320
rect 3344 371278 3372 371311
rect 3332 371272 3384 371278
rect 3332 371214 3384 371220
rect 3330 358456 3386 358465
rect 3330 358391 3386 358400
rect 3344 357474 3372 358391
rect 3332 357468 3384 357474
rect 3332 357410 3384 357416
rect 2778 345400 2834 345409
rect 2778 345335 2834 345344
rect 2792 345234 2820 345335
rect 2780 345228 2832 345234
rect 2780 345170 2832 345176
rect 3146 319288 3202 319297
rect 3146 319223 3202 319232
rect 3160 318850 3188 319223
rect 3148 318844 3200 318850
rect 3148 318786 3200 318792
rect 3238 306232 3294 306241
rect 3238 306167 3294 306176
rect 3146 267200 3202 267209
rect 3146 267135 3202 267144
rect 3160 266762 3188 267135
rect 3148 266756 3200 266762
rect 3148 266698 3200 266704
rect 3146 254144 3202 254153
rect 3146 254079 3202 254088
rect 3160 253978 3188 254079
rect 3148 253972 3200 253978
rect 3148 253914 3200 253920
rect 2778 241088 2834 241097
rect 2778 241023 2834 241032
rect 2792 240242 2820 241023
rect 2780 240236 2832 240242
rect 2780 240178 2832 240184
rect 3146 228032 3202 228041
rect 3146 227967 3202 227976
rect 3160 227798 3188 227967
rect 3148 227792 3200 227798
rect 3148 227734 3200 227740
rect 3146 214976 3202 214985
rect 3146 214911 3202 214920
rect 3160 213994 3188 214911
rect 3148 213988 3200 213994
rect 3148 213930 3200 213936
rect 3146 201920 3202 201929
rect 3146 201855 3148 201864
rect 3200 201855 3202 201864
rect 3148 201826 3200 201832
rect 2778 188864 2834 188873
rect 2778 188799 2834 188808
rect 2792 187746 2820 188799
rect 2780 187740 2832 187746
rect 2780 187682 2832 187688
rect 3148 162920 3200 162926
rect 3146 162888 3148 162897
rect 3200 162888 3202 162897
rect 3146 162823 3202 162832
rect 3252 149734 3280 306167
rect 3330 293176 3386 293185
rect 3330 293111 3386 293120
rect 3240 149728 3292 149734
rect 3240 149670 3292 149676
rect 3238 136776 3294 136785
rect 3238 136711 3240 136720
rect 3292 136711 3294 136720
rect 3240 136682 3292 136688
rect 3240 133952 3292 133958
rect 3240 133894 3292 133900
rect 3148 111784 3200 111790
rect 3148 111726 3200 111732
rect 3160 110673 3188 111726
rect 3146 110664 3202 110673
rect 3146 110599 3202 110608
rect 3252 97617 3280 133894
rect 3238 97608 3294 97617
rect 3238 97543 3294 97552
rect 3344 93854 3372 293111
rect 3160 93826 3372 93854
rect 3160 84862 3188 93826
rect 3436 84946 3464 658135
rect 3514 619168 3570 619177
rect 3514 619103 3570 619112
rect 3528 618322 3556 619103
rect 3516 618316 3568 618322
rect 3516 618258 3568 618264
rect 3606 606112 3662 606121
rect 3606 606047 3662 606056
rect 3514 580000 3570 580009
rect 3514 579935 3570 579944
rect 3528 579698 3556 579935
rect 3516 579692 3568 579698
rect 3516 579634 3568 579640
rect 3514 553888 3570 553897
rect 3514 553823 3570 553832
rect 3252 84918 3464 84946
rect 3148 84856 3200 84862
rect 3148 84798 3200 84804
rect 3252 78985 3280 84918
rect 3332 84856 3384 84862
rect 3332 84798 3384 84804
rect 3424 84856 3476 84862
rect 3424 84798 3476 84804
rect 3344 79354 3372 84798
rect 3332 79348 3384 79354
rect 3332 79290 3384 79296
rect 3436 79121 3464 84798
rect 3528 81161 3556 553823
rect 3620 84862 3648 606047
rect 3882 527912 3938 527921
rect 3882 527847 3938 527856
rect 3790 501800 3846 501809
rect 3790 501735 3846 501744
rect 3698 449576 3754 449585
rect 3698 449511 3754 449520
rect 3608 84856 3660 84862
rect 3608 84798 3660 84804
rect 3608 84720 3660 84726
rect 3608 84662 3660 84668
rect 3514 81152 3570 81161
rect 3514 81087 3570 81096
rect 3620 79257 3648 84662
rect 3712 81297 3740 449511
rect 3804 84726 3832 501735
rect 3896 229770 3924 527847
rect 4066 475688 4122 475697
rect 4066 475623 4122 475632
rect 3974 397488 4030 397497
rect 3974 397423 4030 397432
rect 3884 229764 3936 229770
rect 3884 229706 3936 229712
rect 3882 149832 3938 149841
rect 3882 149767 3938 149776
rect 3896 138718 3924 149767
rect 3884 138712 3936 138718
rect 3884 138654 3936 138660
rect 3884 136672 3936 136678
rect 3884 136614 3936 136620
rect 3792 84720 3844 84726
rect 3792 84662 3844 84668
rect 3792 84584 3844 84590
rect 3792 84526 3844 84532
rect 3698 81288 3754 81297
rect 3698 81223 3754 81232
rect 3804 79393 3832 84526
rect 3790 79384 3846 79393
rect 3790 79319 3846 79328
rect 3606 79248 3662 79257
rect 3606 79183 3662 79192
rect 3422 79112 3478 79121
rect 3422 79047 3478 79056
rect 3238 78976 3294 78985
rect 3238 78911 3294 78920
rect 1398 76528 1454 76537
rect 1398 76463 1454 76472
rect 572 8968 624 8974
rect 572 8910 624 8916
rect 584 480 612 8910
rect 542 -960 654 480
rect 1412 354 1440 76463
rect 2778 75168 2834 75177
rect 2778 75103 2834 75112
rect 2792 16574 2820 75103
rect 3424 71732 3476 71738
rect 3424 71674 3476 71680
rect 3436 71641 3464 71674
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 3424 33040 3476 33046
rect 3424 32982 3476 32988
rect 3436 32473 3464 32982
rect 3422 32464 3478 32473
rect 3422 32399 3478 32408
rect 3424 23316 3476 23322
rect 3424 23258 3476 23264
rect 2792 16546 2912 16574
rect 2884 480 2912 16546
rect 3436 6497 3464 23258
rect 3896 19417 3924 136614
rect 3988 84794 4016 397423
rect 4080 231130 4108 475623
rect 4068 231124 4120 231130
rect 4068 231066 4120 231072
rect 4816 140078 4844 683674
rect 4896 632120 4948 632126
rect 4896 632062 4948 632068
rect 4908 141710 4936 632062
rect 4988 462596 5040 462602
rect 4988 462538 5040 462544
rect 4896 141704 4948 141710
rect 4896 141646 4948 141652
rect 4804 140072 4856 140078
rect 4804 140014 4856 140020
rect 4068 135312 4120 135318
rect 4068 135254 4120 135260
rect 3976 84788 4028 84794
rect 3976 84730 4028 84736
rect 3974 84688 4030 84697
rect 3974 84623 4030 84632
rect 3988 84250 4016 84623
rect 3976 84244 4028 84250
rect 3976 84186 4028 84192
rect 4080 58585 4108 135254
rect 5000 124166 5028 462538
rect 6184 422952 6236 422958
rect 6184 422894 6236 422900
rect 5080 345228 5132 345234
rect 5080 345170 5132 345176
rect 4988 124160 5040 124166
rect 4988 124102 5040 124108
rect 5092 78878 5120 345170
rect 5172 240236 5224 240242
rect 5172 240178 5224 240184
rect 5184 79626 5212 240178
rect 5264 187740 5316 187746
rect 5264 187682 5316 187688
rect 5276 80714 5304 187682
rect 6196 144362 6224 422894
rect 6184 144356 6236 144362
rect 6184 144298 6236 144304
rect 5264 80708 5316 80714
rect 5264 80650 5316 80656
rect 5172 79620 5224 79626
rect 5172 79562 5224 79568
rect 6932 79529 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 23492 703582 24164 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 15844 670744 15896 670750
rect 15844 670686 15896 670692
rect 10324 579692 10376 579698
rect 10324 579634 10376 579640
rect 8944 409964 8996 409970
rect 8944 409906 8996 409912
rect 7564 201884 7616 201890
rect 7564 201826 7616 201832
rect 7576 131102 7604 201826
rect 7564 131096 7616 131102
rect 7564 131038 7616 131044
rect 8956 125594 8984 409906
rect 9036 266756 9088 266762
rect 9036 266698 9088 266704
rect 9048 162178 9076 266698
rect 9036 162172 9088 162178
rect 9036 162114 9088 162120
rect 10336 140146 10364 579634
rect 10416 371272 10468 371278
rect 10416 371214 10468 371220
rect 10428 144430 10456 371214
rect 10416 144424 10468 144430
rect 10416 144366 10468 144372
rect 10324 140140 10376 140146
rect 10324 140082 10376 140088
rect 8944 125588 8996 125594
rect 8944 125530 8996 125536
rect 15856 118658 15884 670686
rect 19984 618316 20036 618322
rect 19984 618258 20036 618264
rect 19996 120086 20024 618258
rect 22744 253972 22796 253978
rect 22744 253914 22796 253920
rect 22756 129742 22784 253914
rect 22836 149728 22888 149734
rect 22836 149670 22888 149676
rect 22744 129736 22796 129742
rect 22744 129678 22796 129684
rect 22848 128314 22876 149670
rect 22836 128308 22888 128314
rect 22836 128250 22888 128256
rect 19984 120080 20036 120086
rect 19984 120022 20036 120028
rect 15844 118652 15896 118658
rect 15844 118594 15896 118600
rect 23492 117298 23520 703582
rect 24136 703474 24164 703582
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 24320 703474 24348 703520
rect 24136 703446 24348 703474
rect 37924 565888 37976 565894
rect 37924 565830 37976 565836
rect 24124 357468 24176 357474
rect 24124 357410 24176 357416
rect 24136 126954 24164 357410
rect 33784 318844 33836 318850
rect 33784 318786 33836 318792
rect 33796 144498 33824 318786
rect 33784 144492 33836 144498
rect 33784 144434 33836 144440
rect 25504 138712 25556 138718
rect 25504 138654 25556 138660
rect 25516 132462 25544 138654
rect 25504 132456 25556 132462
rect 25504 132398 25556 132404
rect 24124 126948 24176 126954
rect 24124 126890 24176 126896
rect 37936 121446 37964 565830
rect 40052 141778 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 104912 703582 105308 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 43444 514820 43496 514826
rect 43444 514762 43496 514768
rect 40040 141772 40092 141778
rect 40040 141714 40092 141720
rect 43456 122806 43484 514762
rect 69664 396772 69716 396778
rect 69664 396714 69716 396720
rect 69676 385014 69704 396714
rect 68284 385008 68336 385014
rect 68284 384950 68336 384956
rect 69664 385008 69716 385014
rect 69664 384950 69716 384956
rect 68296 359106 68324 384950
rect 65708 359100 65760 359106
rect 65708 359042 65760 359048
rect 68284 359100 68336 359106
rect 68284 359042 68336 359048
rect 65720 358222 65748 359042
rect 64144 358216 64196 358222
rect 64144 358158 64196 358164
rect 65708 358216 65760 358222
rect 65708 358158 65760 358164
rect 54484 358080 54536 358086
rect 54484 358022 54536 358028
rect 54496 349518 54524 358022
rect 51724 349512 51776 349518
rect 51724 349454 51776 349460
rect 54484 349512 54536 349518
rect 54484 349454 54536 349460
rect 46388 334008 46440 334014
rect 46388 333950 46440 333956
rect 46400 331566 46428 333950
rect 44916 331560 44968 331566
rect 44916 331502 44968 331508
rect 46388 331560 46440 331566
rect 46388 331502 46440 331508
rect 44824 244996 44876 245002
rect 44824 244938 44876 244944
rect 44836 231062 44864 244938
rect 44824 231056 44876 231062
rect 44824 230998 44876 231004
rect 44928 230586 44956 331502
rect 51736 330546 51764 349454
rect 62120 340196 62172 340202
rect 62120 340138 62172 340144
rect 62132 337414 62160 340138
rect 53840 337408 53892 337414
rect 53840 337350 53892 337356
rect 62120 337408 62172 337414
rect 62120 337350 62172 337356
rect 53852 334014 53880 337350
rect 53840 334008 53892 334014
rect 53840 333950 53892 333956
rect 62856 331900 62908 331906
rect 62856 331842 62908 331848
rect 45008 330540 45060 330546
rect 45008 330482 45060 330488
rect 51724 330540 51776 330546
rect 51724 330482 51776 330488
rect 44916 230580 44968 230586
rect 44916 230522 44968 230528
rect 45020 228410 45048 330482
rect 62764 319456 62816 319462
rect 62764 319398 62816 319404
rect 61476 318436 61528 318442
rect 61476 318378 61528 318384
rect 61488 311234 61516 318378
rect 62120 312180 62172 312186
rect 62120 312122 62172 312128
rect 60004 311228 60056 311234
rect 60004 311170 60056 311176
rect 61476 311228 61528 311234
rect 61476 311170 61528 311176
rect 60016 291174 60044 311170
rect 62132 307290 62160 312122
rect 60096 307284 60148 307290
rect 60096 307226 60148 307232
rect 62120 307284 62172 307290
rect 62120 307226 62172 307232
rect 58624 291168 58676 291174
rect 58624 291110 58676 291116
rect 60004 291168 60056 291174
rect 60004 291110 60056 291116
rect 55220 289808 55272 289814
rect 55220 289750 55272 289756
rect 55232 282962 55260 289750
rect 55864 289128 55916 289134
rect 55864 289070 55916 289076
rect 55140 282934 55260 282962
rect 54208 281444 54260 281450
rect 54208 281386 54260 281392
rect 53288 280832 53340 280838
rect 53288 280774 53340 280780
rect 53104 279472 53156 279478
rect 53104 279414 53156 279420
rect 50344 274916 50396 274922
rect 50344 274858 50396 274864
rect 50356 268394 50384 274858
rect 50436 274780 50488 274786
rect 50436 274722 50488 274728
rect 45284 268388 45336 268394
rect 45284 268330 45336 268336
rect 50344 268388 50396 268394
rect 50344 268330 50396 268336
rect 45192 256760 45244 256766
rect 45192 256702 45244 256708
rect 45100 240848 45152 240854
rect 45100 240790 45152 240796
rect 45112 233170 45140 240790
rect 45100 233164 45152 233170
rect 45100 233106 45152 233112
rect 45008 228404 45060 228410
rect 45008 228346 45060 228352
rect 45204 226302 45232 256702
rect 45192 226296 45244 226302
rect 45192 226238 45244 226244
rect 45296 217666 45324 268330
rect 50448 266422 50476 274722
rect 53116 272066 53144 279414
rect 53196 274712 53248 274718
rect 53196 274654 53248 274660
rect 51724 272060 51776 272066
rect 51724 272002 51776 272008
rect 53104 272060 53156 272066
rect 53104 272002 53156 272008
rect 51080 270496 51132 270502
rect 51080 270438 51132 270444
rect 51092 266422 51120 270438
rect 50436 266416 50488 266422
rect 50436 266358 50488 266364
rect 51080 266416 51132 266422
rect 51080 266358 51132 266364
rect 46204 266348 46256 266354
rect 46204 266290 46256 266296
rect 48320 266348 48372 266354
rect 48320 266290 48372 266296
rect 45744 259140 45796 259146
rect 45744 259082 45796 259088
rect 45652 255332 45704 255338
rect 45652 255274 45704 255280
rect 45664 248414 45692 255274
rect 45572 248386 45692 248414
rect 45468 240780 45520 240786
rect 45468 240722 45520 240728
rect 45376 238808 45428 238814
rect 45376 238750 45428 238756
rect 45388 233238 45416 238750
rect 45376 233232 45428 233238
rect 45376 233174 45428 233180
rect 45480 232830 45508 240722
rect 45572 233306 45600 248386
rect 45652 240576 45704 240582
rect 45652 240518 45704 240524
rect 45560 233300 45612 233306
rect 45560 233242 45612 233248
rect 45560 232892 45612 232898
rect 45560 232834 45612 232840
rect 45468 232824 45520 232830
rect 45468 232766 45520 232772
rect 45572 230382 45600 232834
rect 45560 230376 45612 230382
rect 45560 230318 45612 230324
rect 45664 219434 45692 240518
rect 45756 233374 45784 259082
rect 46216 256766 46244 266290
rect 48332 262290 48360 266290
rect 51736 263634 51764 272002
rect 53208 267734 53236 274654
rect 53300 270502 53328 280774
rect 53380 280220 53432 280226
rect 53380 280162 53432 280168
rect 53392 274786 53420 280162
rect 54220 279478 54248 281386
rect 55140 280226 55168 282934
rect 55128 280220 55180 280226
rect 55128 280162 55180 280168
rect 54208 279472 54260 279478
rect 54208 279414 54260 279420
rect 54484 278792 54536 278798
rect 54484 278734 54536 278740
rect 53840 277364 53892 277370
rect 53840 277306 53892 277312
rect 53380 274780 53432 274786
rect 53380 274722 53432 274728
rect 53852 274718 53880 277306
rect 53840 274712 53892 274718
rect 53840 274654 53892 274660
rect 53288 270496 53340 270502
rect 53288 270438 53340 270444
rect 53116 267706 53236 267734
rect 49700 263628 49752 263634
rect 49700 263570 49752 263576
rect 51724 263628 51776 263634
rect 51724 263570 51776 263576
rect 48240 262262 48360 262290
rect 48240 259146 48268 262262
rect 48228 259140 48280 259146
rect 48228 259082 48280 259088
rect 49712 258602 49740 263570
rect 46940 258596 46992 258602
rect 46940 258538 46992 258544
rect 49700 258596 49752 258602
rect 49700 258538 49752 258544
rect 46204 256760 46256 256766
rect 46204 256702 46256 256708
rect 46952 255338 46980 258538
rect 50436 256692 50488 256698
rect 50436 256634 50488 256640
rect 46940 255332 46992 255338
rect 46940 255274 46992 255280
rect 50448 253978 50476 256634
rect 47584 253972 47636 253978
rect 47584 253914 47636 253920
rect 50436 253972 50488 253978
rect 50436 253914 50488 253920
rect 46204 253904 46256 253910
rect 46204 253846 46256 253852
rect 45836 245676 45888 245682
rect 45836 245618 45888 245624
rect 45848 238814 45876 245618
rect 46216 245002 46244 253846
rect 47596 245682 47624 253914
rect 53116 252890 53144 267706
rect 54496 266490 54524 278734
rect 55876 274922 55904 289070
rect 57244 287700 57296 287706
rect 57244 287642 57296 287648
rect 56508 284300 56560 284306
rect 56508 284242 56560 284248
rect 56520 281450 56548 284242
rect 56508 281444 56560 281450
rect 56508 281386 56560 281392
rect 57256 277438 57284 287642
rect 58636 284374 58664 291110
rect 60108 289882 60136 307226
rect 62776 299130 62804 319398
rect 62868 318442 62896 331842
rect 64156 319462 64184 358158
rect 70308 332580 70360 332586
rect 70308 332522 70360 332528
rect 70320 328098 70348 332522
rect 68192 328092 68244 328098
rect 68192 328034 68244 328040
rect 70308 328092 70360 328098
rect 70308 328034 70360 328040
rect 68204 320142 68232 328034
rect 66904 320136 66956 320142
rect 66904 320078 66956 320084
rect 68192 320136 68244 320142
rect 68192 320078 68244 320084
rect 64144 319456 64196 319462
rect 64144 319398 64196 319404
rect 62856 318436 62908 318442
rect 62856 318378 62908 318384
rect 66916 312186 66944 320078
rect 66904 312180 66956 312186
rect 66904 312122 66956 312128
rect 61568 299124 61620 299130
rect 61568 299066 61620 299072
rect 62764 299124 62816 299130
rect 62764 299066 62816 299072
rect 61580 294030 61608 299066
rect 60188 294024 60240 294030
rect 60188 293966 60240 293972
rect 61568 294024 61620 294030
rect 61568 293966 61620 293972
rect 60096 289876 60148 289882
rect 60096 289818 60148 289824
rect 58624 284368 58676 284374
rect 58624 284310 58676 284316
rect 60200 282946 60228 293966
rect 66996 291236 67048 291242
rect 66996 291178 67048 291184
rect 67008 289134 67036 291178
rect 66996 289128 67048 289134
rect 66996 289070 67048 289076
rect 71792 287706 71820 702986
rect 89180 702434 89208 703520
rect 88352 702406 89208 702434
rect 86868 382968 86920 382974
rect 86868 382910 86920 382916
rect 86880 379098 86908 382910
rect 79324 379092 79376 379098
rect 79324 379034 79376 379040
rect 86868 379092 86920 379098
rect 86868 379034 86920 379040
rect 73804 359508 73856 359514
rect 73804 359450 73856 359456
rect 73816 340202 73844 359450
rect 79336 358086 79364 379034
rect 87512 364540 87564 364546
rect 87512 364482 87564 364488
rect 87524 358970 87552 364482
rect 86224 358964 86276 358970
rect 86224 358906 86276 358912
rect 87512 358964 87564 358970
rect 87512 358906 87564 358912
rect 79324 358080 79376 358086
rect 79324 358022 79376 358028
rect 86236 353326 86264 358906
rect 85028 353320 85080 353326
rect 85028 353262 85080 353268
rect 86224 353320 86276 353326
rect 86224 353262 86276 353268
rect 85040 351354 85068 353262
rect 82820 351348 82872 351354
rect 82820 351290 82872 351296
rect 85028 351348 85080 351354
rect 85028 351290 85080 351296
rect 82832 346458 82860 351290
rect 82820 346452 82872 346458
rect 82820 346394 82872 346400
rect 78680 346384 78732 346390
rect 78680 346326 78732 346332
rect 78692 345014 78720 346326
rect 78600 344986 78720 345014
rect 78600 340950 78628 344986
rect 75920 340944 75972 340950
rect 75920 340886 75972 340892
rect 78588 340944 78640 340950
rect 78588 340886 78640 340892
rect 73804 340196 73856 340202
rect 73804 340138 73856 340144
rect 75932 338178 75960 340886
rect 75840 338150 75960 338178
rect 75840 336802 75868 338150
rect 73160 336796 73212 336802
rect 73160 336738 73212 336744
rect 75828 336796 75880 336802
rect 75828 336738 75880 336744
rect 73172 335354 73200 336738
rect 73080 335326 73200 335354
rect 73080 332654 73108 335326
rect 73068 332648 73120 332654
rect 73068 332590 73120 332596
rect 88352 331906 88380 702406
rect 101404 519580 101456 519586
rect 101404 519522 101456 519528
rect 101416 511970 101444 519522
rect 98644 511964 98696 511970
rect 98644 511906 98696 511912
rect 101404 511964 101456 511970
rect 101404 511906 101456 511912
rect 98656 466478 98684 511906
rect 102784 499588 102836 499594
rect 102784 499530 102836 499536
rect 102796 477562 102824 499530
rect 101404 477556 101456 477562
rect 101404 477498 101456 477504
rect 102784 477556 102836 477562
rect 102784 477498 102836 477504
rect 95884 466472 95936 466478
rect 95884 466414 95936 466420
rect 98644 466472 98696 466478
rect 98644 466414 98696 466420
rect 95896 429758 95924 466414
rect 101416 452674 101444 477498
rect 101404 452668 101456 452674
rect 101404 452610 101456 452616
rect 97264 452600 97316 452606
rect 97264 452542 97316 452548
rect 93124 429752 93176 429758
rect 93124 429694 93176 429700
rect 95884 429752 95936 429758
rect 95884 429694 95936 429700
rect 88984 384464 89036 384470
rect 88984 384406 89036 384412
rect 88996 359514 89024 384406
rect 91928 379568 91980 379574
rect 91928 379510 91980 379516
rect 91940 377874 91968 379510
rect 90364 377868 90416 377874
rect 90364 377810 90416 377816
rect 91928 377868 91980 377874
rect 91928 377810 91980 377816
rect 90376 364546 90404 377810
rect 90364 364540 90416 364546
rect 90364 364482 90416 364488
rect 88984 359508 89036 359514
rect 88984 359450 89036 359456
rect 88340 331900 88392 331906
rect 88340 331842 88392 331848
rect 84844 315308 84896 315314
rect 84844 315250 84896 315256
rect 73160 294636 73212 294642
rect 73160 294578 73212 294584
rect 73172 291242 73200 294578
rect 73160 291236 73212 291242
rect 73160 291178 73212 291184
rect 71780 287700 71832 287706
rect 71780 287642 71832 287648
rect 84856 284374 84884 315250
rect 93136 311914 93164 429694
rect 97276 415070 97304 452542
rect 100024 424380 100076 424386
rect 100024 424322 100076 424328
rect 95884 415064 95936 415070
rect 95884 415006 95936 415012
rect 97264 415064 97316 415070
rect 97264 415006 97316 415012
rect 93216 406428 93268 406434
rect 93216 406370 93268 406376
rect 93228 384470 93256 406370
rect 95896 393378 95924 415006
rect 100036 406434 100064 424322
rect 100024 406428 100076 406434
rect 100024 406370 100076 406376
rect 93308 393372 93360 393378
rect 93308 393314 93360 393320
rect 95884 393372 95936 393378
rect 95884 393314 95936 393320
rect 93216 384464 93268 384470
rect 93216 384406 93268 384412
rect 93320 379574 93348 393314
rect 97540 385076 97592 385082
rect 97540 385018 97592 385024
rect 97552 382974 97580 385018
rect 97540 382968 97592 382974
rect 97540 382910 97592 382916
rect 93308 379568 93360 379574
rect 93308 379510 93360 379516
rect 104912 315314 104940 703582
rect 105280 703474 105308 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 136652 703582 137692 703610
rect 105464 703474 105492 703520
rect 105280 703446 105492 703474
rect 135904 641776 135956 641782
rect 135904 641718 135956 641724
rect 135916 603158 135944 641718
rect 134524 603152 134576 603158
rect 134524 603094 134576 603100
rect 135904 603152 135956 603158
rect 135904 603094 135956 603100
rect 134536 583778 134564 603094
rect 134524 583772 134576 583778
rect 134524 583714 134576 583720
rect 130384 583704 130436 583710
rect 130384 583646 130436 583652
rect 127624 567860 127676 567866
rect 127624 567802 127676 567808
rect 127636 558890 127664 567802
rect 124864 558884 124916 558890
rect 124864 558826 124916 558832
rect 127624 558884 127676 558890
rect 127624 558826 127676 558832
rect 124876 545630 124904 558826
rect 130396 550254 130424 583646
rect 129004 550248 129056 550254
rect 129004 550190 129056 550196
rect 130384 550248 130436 550254
rect 130384 550190 130436 550196
rect 122104 545624 122156 545630
rect 122104 545566 122156 545572
rect 124864 545624 124916 545630
rect 124864 545566 124916 545572
rect 122116 527202 122144 545566
rect 123484 536104 123536 536110
rect 123484 536046 123536 536052
rect 117136 527196 117188 527202
rect 117136 527138 117188 527144
rect 122104 527196 122156 527202
rect 122104 527138 122156 527144
rect 106924 525088 106976 525094
rect 106924 525030 106976 525036
rect 106936 514078 106964 525030
rect 117148 519586 117176 527138
rect 117136 519580 117188 519586
rect 117136 519522 117188 519528
rect 105544 514072 105596 514078
rect 105544 514014 105596 514020
rect 106924 514072 106976 514078
rect 106924 514014 106976 514020
rect 105556 499594 105584 514014
rect 123496 508570 123524 536046
rect 129016 525094 129044 550190
rect 133144 544400 133196 544406
rect 133144 544342 133196 544348
rect 133156 536110 133184 544342
rect 133144 536104 133196 536110
rect 133144 536046 133196 536052
rect 129004 525088 129056 525094
rect 129004 525030 129056 525036
rect 127624 516792 127676 516798
rect 127624 516734 127676 516740
rect 113824 508564 113876 508570
rect 113824 508506 113876 508512
rect 123484 508564 123536 508570
rect 123484 508506 123536 508512
rect 105544 499588 105596 499594
rect 105544 499530 105596 499536
rect 113836 447778 113864 508506
rect 127636 482322 127664 516734
rect 119344 482316 119396 482322
rect 119344 482258 119396 482264
rect 127624 482316 127676 482322
rect 127624 482258 127676 482264
rect 119356 469266 119384 482258
rect 116584 469260 116636 469266
rect 116584 469202 116636 469208
rect 119344 469260 119396 469266
rect 119344 469202 119396 469208
rect 108304 447772 108356 447778
rect 108304 447714 108356 447720
rect 113824 447772 113876 447778
rect 113824 447714 113876 447720
rect 108316 424386 108344 447714
rect 108304 424380 108356 424386
rect 108304 424322 108356 424328
rect 116596 411942 116624 469202
rect 108304 411936 108356 411942
rect 108304 411878 108356 411884
rect 116584 411936 116636 411942
rect 116584 411878 116636 411884
rect 108316 394670 108344 411878
rect 136652 396778 136680 703582
rect 137664 703474 137692 703582
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 234632 703582 235028 703610
rect 137848 703474 137876 703520
rect 137664 703446 137876 703474
rect 154132 699718 154160 703520
rect 170324 702434 170352 703520
rect 169772 702406 170352 702434
rect 152464 699712 152516 699718
rect 152464 699654 152516 699660
rect 154120 699712 154172 699718
rect 154120 699654 154172 699660
rect 152476 689314 152504 699654
rect 150440 689308 150492 689314
rect 150440 689250 150492 689256
rect 152464 689308 152516 689314
rect 152464 689250 152516 689256
rect 150452 683738 150480 689250
rect 149060 683732 149112 683738
rect 149060 683674 149112 683680
rect 150440 683732 150492 683738
rect 150440 683674 150492 683680
rect 149072 680354 149100 683674
rect 148980 680326 149100 680354
rect 148980 676394 149008 680326
rect 146208 676388 146260 676394
rect 146208 676330 146260 676336
rect 148968 676388 149020 676394
rect 148968 676330 149020 676336
rect 146220 674490 146248 676330
rect 143540 674484 143592 674490
rect 143540 674426 143592 674432
rect 146208 674484 146260 674490
rect 146208 674426 146260 674432
rect 143552 667962 143580 674426
rect 143540 667956 143592 667962
rect 143540 667898 143592 667904
rect 140044 667888 140096 667894
rect 140044 667830 140096 667836
rect 140056 651438 140084 667830
rect 138664 651432 138716 651438
rect 138664 651374 138716 651380
rect 140044 651432 140096 651438
rect 140044 651374 140096 651380
rect 138676 641782 138704 651374
rect 138664 641776 138716 641782
rect 138664 641718 138716 641724
rect 153844 605124 153896 605130
rect 153844 605066 153896 605072
rect 153856 575278 153884 605066
rect 149060 575272 149112 575278
rect 149060 575214 149112 575220
rect 153844 575272 153896 575278
rect 153844 575214 153896 575220
rect 149072 572014 149100 575214
rect 137284 572008 137336 572014
rect 137284 571950 137336 571956
rect 149060 572008 149112 572014
rect 149060 571950 149112 571956
rect 137296 567866 137324 571950
rect 137284 567860 137336 567866
rect 137284 567802 137336 567808
rect 163504 554056 163556 554062
rect 163504 553998 163556 554004
rect 163516 547194 163544 553998
rect 146116 547188 146168 547194
rect 146116 547130 146168 547136
rect 163504 547188 163556 547194
rect 163504 547130 163556 547136
rect 146128 544406 146156 547130
rect 146116 544400 146168 544406
rect 146116 544342 146168 544348
rect 156604 537532 156656 537538
rect 156604 537474 156656 537480
rect 156616 516798 156644 537474
rect 156604 516792 156656 516798
rect 156604 516734 156656 516740
rect 167644 478848 167696 478854
rect 167644 478790 167696 478796
rect 167656 423638 167684 478790
rect 166264 423632 166316 423638
rect 166264 423574 166316 423580
rect 167644 423632 167696 423638
rect 167644 423574 167696 423580
rect 166276 415138 166304 423574
rect 164792 415132 164844 415138
rect 164792 415074 164844 415080
rect 166264 415132 166316 415138
rect 166264 415074 166316 415080
rect 164804 407182 164832 415074
rect 161848 407176 161900 407182
rect 161848 407118 161900 407124
rect 164792 407176 164844 407182
rect 164792 407118 164844 407124
rect 161860 406434 161888 407118
rect 160100 406428 160152 406434
rect 160100 406370 160152 406376
rect 161848 406428 161900 406434
rect 161848 406370 161900 406376
rect 160112 404394 160140 406370
rect 160100 404388 160152 404394
rect 160100 404330 160152 404336
rect 157340 404320 157392 404326
rect 157340 404262 157392 404268
rect 157352 400246 157380 404262
rect 157340 400240 157392 400246
rect 157340 400182 157392 400188
rect 153844 400172 153896 400178
rect 153844 400114 153896 400120
rect 136640 396772 136692 396778
rect 136640 396714 136692 396720
rect 105544 394664 105596 394670
rect 105544 394606 105596 394612
rect 108304 394664 108356 394670
rect 108304 394606 108356 394612
rect 105556 385082 105584 394606
rect 153856 392018 153884 400114
rect 153844 392012 153896 392018
rect 153844 391954 153896 391960
rect 146944 391944 146996 391950
rect 146944 391886 146996 391892
rect 105544 385076 105596 385082
rect 105544 385018 105596 385024
rect 146956 358834 146984 391886
rect 146944 358828 146996 358834
rect 146944 358770 146996 358776
rect 142804 358760 142856 358766
rect 142804 358702 142856 358708
rect 142816 353326 142844 358702
rect 140780 353320 140832 353326
rect 140780 353262 140832 353268
rect 142804 353320 142856 353326
rect 142804 353262 142856 353268
rect 140792 350606 140820 353262
rect 137284 350600 137336 350606
rect 137284 350542 137336 350548
rect 140780 350600 140832 350606
rect 140780 350542 140832 350548
rect 137296 329594 137324 350542
rect 134524 329588 134576 329594
rect 134524 329530 134576 329536
rect 137284 329588 137336 329594
rect 137284 329530 137336 329536
rect 134536 320210 134564 329530
rect 134524 320204 134576 320210
rect 134524 320146 134576 320152
rect 126244 320136 126296 320142
rect 126244 320078 126296 320084
rect 104900 315308 104952 315314
rect 104900 315250 104952 315256
rect 90364 311908 90416 311914
rect 90364 311850 90416 311856
rect 93124 311908 93176 311914
rect 93124 311850 93176 311856
rect 90376 294642 90404 311850
rect 90364 294636 90416 294642
rect 90364 294578 90416 294584
rect 126256 292602 126284 320078
rect 124864 292596 124916 292602
rect 124864 292538 124916 292544
rect 126244 292596 126296 292602
rect 126244 292538 126296 292544
rect 84844 284368 84896 284374
rect 84844 284310 84896 284316
rect 82084 284300 82136 284306
rect 82084 284242 82136 284248
rect 57980 282940 58032 282946
rect 57980 282882 58032 282888
rect 60188 282940 60240 282946
rect 60188 282882 60240 282888
rect 57992 280242 58020 282882
rect 57900 280214 58020 280242
rect 57900 278798 57928 280214
rect 57888 278792 57940 278798
rect 57888 278734 57940 278740
rect 57244 277432 57296 277438
rect 57244 277374 57296 277380
rect 82096 276690 82124 284242
rect 55956 276684 56008 276690
rect 55956 276626 56008 276632
rect 82084 276684 82136 276690
rect 82084 276626 82136 276632
rect 55864 274916 55916 274922
rect 55864 274858 55916 274864
rect 53196 266484 53248 266490
rect 53196 266426 53248 266432
rect 54484 266484 54536 266490
rect 54484 266426 54536 266432
rect 53208 254046 53236 266426
rect 55968 266422 55996 276626
rect 124876 273290 124904 292538
rect 169772 280838 169800 702406
rect 202800 699718 202828 703520
rect 218992 699718 219020 703520
rect 196624 699712 196676 699718
rect 196624 699654 196676 699660
rect 202788 699712 202840 699718
rect 202788 699654 202840 699660
rect 217324 699712 217376 699718
rect 217324 699654 217376 699660
rect 218980 699712 219032 699718
rect 218980 699654 219032 699660
rect 189724 645176 189776 645182
rect 189724 645118 189776 645124
rect 189736 636886 189764 645118
rect 179420 636880 179472 636886
rect 179420 636822 179472 636828
rect 189724 636880 189776 636886
rect 189724 636822 189776 636828
rect 179432 630698 179460 636822
rect 174452 630692 174504 630698
rect 174452 630634 174504 630640
rect 179420 630692 179472 630698
rect 179420 630634 179472 630640
rect 174464 629066 174492 630634
rect 171784 629060 171836 629066
rect 171784 629002 171836 629008
rect 174452 629060 174504 629066
rect 174452 629002 174504 629008
rect 171796 605130 171824 629002
rect 196636 623830 196664 699654
rect 217336 688702 217364 699654
rect 217324 688696 217376 688702
rect 217324 688638 217376 688644
rect 213184 688628 213236 688634
rect 213184 688570 213236 688576
rect 213196 672110 213224 688570
rect 224224 685160 224276 685166
rect 224224 685102 224276 685108
rect 224236 673810 224264 685102
rect 220820 673804 220872 673810
rect 220820 673746 220872 673752
rect 224224 673804 224276 673810
rect 224224 673746 224276 673752
rect 211528 672104 211580 672110
rect 211528 672046 211580 672052
rect 213184 672104 213236 672110
rect 213184 672046 213236 672052
rect 211540 670750 211568 672046
rect 208400 670744 208452 670750
rect 208400 670686 208452 670692
rect 211528 670744 211580 670750
rect 211528 670686 211580 670692
rect 208412 667978 208440 670686
rect 208320 667950 208440 667978
rect 208320 665922 208348 667950
rect 220832 667690 220860 673746
rect 218704 667684 218756 667690
rect 218704 667626 218756 667632
rect 220820 667684 220872 667690
rect 220820 667626 220872 667632
rect 206284 665916 206336 665922
rect 206284 665858 206336 665864
rect 208308 665916 208360 665922
rect 208308 665858 208360 665864
rect 201408 647896 201460 647902
rect 201408 647838 201460 647844
rect 201420 645182 201448 647838
rect 206296 647222 206324 665858
rect 218716 662454 218744 667626
rect 215300 662448 215352 662454
rect 215300 662390 215352 662396
rect 218704 662448 218756 662454
rect 218704 662390 218756 662396
rect 215312 657626 215340 662390
rect 211804 657620 211856 657626
rect 211804 657562 211856 657568
rect 215300 657620 215352 657626
rect 215300 657562 215352 657568
rect 211816 647902 211844 657562
rect 211804 647896 211856 647902
rect 211804 647838 211856 647844
rect 204904 647216 204956 647222
rect 204904 647158 204956 647164
rect 206284 647216 206336 647222
rect 206284 647158 206336 647164
rect 201408 645176 201460 645182
rect 201408 645118 201460 645124
rect 193864 623824 193916 623830
rect 193864 623766 193916 623772
rect 196624 623824 196676 623830
rect 196624 623766 196676 623772
rect 193876 610706 193904 623766
rect 191104 610700 191156 610706
rect 191104 610642 191156 610648
rect 193864 610700 193916 610706
rect 193864 610642 193916 610648
rect 171784 605124 171836 605130
rect 171784 605066 171836 605072
rect 191116 599894 191144 610642
rect 204916 601730 204944 647158
rect 233884 616820 233936 616826
rect 233884 616762 233936 616768
rect 232596 610292 232648 610298
rect 232596 610234 232648 610240
rect 232504 603152 232556 603158
rect 232504 603094 232556 603100
rect 203616 601724 203668 601730
rect 203616 601666 203668 601672
rect 204904 601724 204956 601730
rect 204904 601666 204956 601672
rect 184204 599888 184256 599894
rect 184204 599830 184256 599836
rect 191104 599888 191156 599894
rect 191104 599830 191156 599836
rect 184216 592074 184244 599830
rect 203628 599690 203656 601666
rect 224408 600976 224460 600982
rect 224408 600918 224460 600924
rect 202144 599684 202196 599690
rect 202144 599626 202196 599632
rect 203616 599684 203668 599690
rect 203616 599626 203668 599632
rect 181444 592068 181496 592074
rect 181444 592010 181496 592016
rect 184204 592068 184256 592074
rect 184204 592010 184256 592016
rect 181456 554062 181484 592010
rect 202156 560998 202184 599626
rect 224420 598194 224448 600918
rect 220820 598188 220872 598194
rect 220820 598130 220872 598136
rect 224408 598188 224460 598194
rect 224408 598130 224460 598136
rect 220832 594862 220860 598130
rect 214564 594856 214616 594862
rect 214564 594798 214616 594804
rect 220820 594856 220872 594862
rect 220820 594798 220872 594804
rect 214576 578202 214604 594798
rect 211804 578196 211856 578202
rect 211804 578138 211856 578144
rect 214564 578196 214616 578202
rect 214564 578138 214616 578144
rect 211816 565010 211844 578138
rect 232516 572762 232544 603094
rect 232608 600982 232636 610234
rect 233896 603158 233924 616762
rect 234632 610298 234660 703582
rect 235000 703474 235028 703582
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 412652 703582 413508 703610
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 267660 700330 267688 703520
rect 254584 700324 254636 700330
rect 254584 700266 254636 700272
rect 267648 700324 267700 700330
rect 267648 700266 267700 700272
rect 254596 689314 254624 700266
rect 283852 697610 283880 703520
rect 300136 700398 300164 703520
rect 332520 703050 332548 703520
rect 331220 703044 331272 703050
rect 331220 702986 331272 702992
rect 332508 703044 332560 703050
rect 332508 702986 332560 702992
rect 300124 700392 300176 700398
rect 300124 700334 300176 700340
rect 303252 700392 303304 700398
rect 303252 700334 303304 700340
rect 282184 697604 282236 697610
rect 282184 697546 282236 697552
rect 283840 697604 283892 697610
rect 283840 697546 283892 697552
rect 239036 689308 239088 689314
rect 239036 689250 239088 689256
rect 254584 689308 254636 689314
rect 254584 689250 254636 689256
rect 239048 685166 239076 689250
rect 239036 685160 239088 685166
rect 239036 685102 239088 685108
rect 282196 681018 282224 697546
rect 303264 693462 303292 700334
rect 303252 693456 303304 693462
rect 303252 693398 303304 693404
rect 316040 693456 316092 693462
rect 316040 693398 316092 693404
rect 316052 688226 316080 693398
rect 331232 688906 331260 702986
rect 348804 699854 348832 703520
rect 364996 702434 365024 703520
rect 364352 702406 365024 702434
rect 348792 699848 348844 699854
rect 348792 699790 348844 699796
rect 351184 699848 351236 699854
rect 351184 699790 351236 699796
rect 351196 692102 351224 699790
rect 351184 692096 351236 692102
rect 351184 692038 351236 692044
rect 358084 692096 358136 692102
rect 358084 692038 358136 692044
rect 331220 688900 331272 688906
rect 331220 688842 331272 688848
rect 334624 688900 334676 688906
rect 334624 688842 334676 688848
rect 316040 688220 316092 688226
rect 316040 688162 316092 688168
rect 323584 688220 323636 688226
rect 323584 688162 323636 688168
rect 261484 681012 261536 681018
rect 261484 680954 261536 680960
rect 282184 681012 282236 681018
rect 282184 680954 282236 680960
rect 261496 666602 261524 680954
rect 261484 666596 261536 666602
rect 261484 666538 261536 666544
rect 258724 666528 258776 666534
rect 258724 666470 258776 666476
rect 258736 654158 258764 666470
rect 323596 662386 323624 688162
rect 323584 662380 323636 662386
rect 323584 662322 323636 662328
rect 326620 662380 326672 662386
rect 326620 662322 326672 662328
rect 326632 659258 326660 662322
rect 326620 659252 326672 659258
rect 326620 659194 326672 659200
rect 330024 659252 330076 659258
rect 330024 659194 330076 659200
rect 330036 656198 330064 659194
rect 330024 656192 330076 656198
rect 330024 656134 330076 656140
rect 257436 654152 257488 654158
rect 257436 654094 257488 654100
rect 258724 654152 258776 654158
rect 258724 654094 258776 654100
rect 257448 651438 257476 654094
rect 255320 651432 255372 651438
rect 255320 651374 255372 651380
rect 257436 651432 257488 651438
rect 257436 651374 257488 651380
rect 255332 645182 255360 651374
rect 334636 646542 334664 688842
rect 358096 681086 358124 692038
rect 364352 690470 364380 702406
rect 364340 690464 364392 690470
rect 364340 690406 364392 690412
rect 369860 690464 369912 690470
rect 369860 690406 369912 690412
rect 369872 688226 369900 690406
rect 369860 688220 369912 688226
rect 369860 688162 369912 688168
rect 372620 688220 372672 688226
rect 372620 688162 372672 688168
rect 372632 683670 372660 688162
rect 372620 683664 372672 683670
rect 372620 683606 372672 683612
rect 375380 683664 375432 683670
rect 375380 683606 375432 683612
rect 358084 681080 358136 681086
rect 358084 681022 358136 681028
rect 360476 681080 360528 681086
rect 360476 681022 360528 681028
rect 360488 678298 360516 681022
rect 375392 681018 375420 683606
rect 375380 681012 375432 681018
rect 375380 680954 375432 680960
rect 389180 681012 389232 681018
rect 389180 680954 389232 680960
rect 360476 678292 360528 678298
rect 360476 678234 360528 678240
rect 369124 678292 369176 678298
rect 369124 678234 369176 678240
rect 369136 675510 369164 678234
rect 369124 675504 369176 675510
rect 369124 675446 369176 675452
rect 378784 675504 378836 675510
rect 378784 675446 378836 675452
rect 378796 664494 378824 675446
rect 389192 675238 389220 680954
rect 389180 675232 389232 675238
rect 389180 675174 389232 675180
rect 393320 675232 393372 675238
rect 393320 675174 393372 675180
rect 393332 673266 393360 675174
rect 393320 673260 393372 673266
rect 393320 673202 393372 673208
rect 396448 673260 396500 673266
rect 396448 673202 396500 673208
rect 378784 664488 378836 664494
rect 378784 664430 378836 664436
rect 387064 664488 387116 664494
rect 387064 664430 387116 664436
rect 336740 656192 336792 656198
rect 336740 656134 336792 656140
rect 336752 649330 336780 656134
rect 387076 652322 387104 664430
rect 387064 652316 387116 652322
rect 387064 652258 387116 652264
rect 395344 652316 395396 652322
rect 395344 652258 395396 652264
rect 336740 649324 336792 649330
rect 336740 649266 336792 649272
rect 345664 649324 345716 649330
rect 345664 649266 345716 649272
rect 334624 646536 334676 646542
rect 334624 646478 334676 646484
rect 342904 646536 342956 646542
rect 342904 646478 342956 646484
rect 245568 645176 245620 645182
rect 245568 645118 245620 645124
rect 255320 645176 255372 645182
rect 255320 645118 255372 645124
rect 245580 640354 245608 645118
rect 243544 640348 243596 640354
rect 243544 640290 243596 640296
rect 245568 640348 245620 640354
rect 245568 640290 245620 640296
rect 243556 623830 243584 640290
rect 243544 623824 243596 623830
rect 243544 623766 243596 623772
rect 239956 623756 240008 623762
rect 239956 623698 240008 623704
rect 239968 621042 239996 623698
rect 237380 621036 237432 621042
rect 237380 620978 237432 620984
rect 239956 621036 240008 621042
rect 239956 620978 240008 620984
rect 237392 616894 237420 620978
rect 237380 616888 237432 616894
rect 237380 616830 237432 616836
rect 342916 616146 342944 646478
rect 345676 644366 345704 649266
rect 345664 644360 345716 644366
rect 345664 644302 345716 644308
rect 353944 644360 353996 644366
rect 353944 644302 353996 644308
rect 353956 622402 353984 644302
rect 353944 622396 353996 622402
rect 353944 622338 353996 622344
rect 356704 622396 356756 622402
rect 356704 622338 356756 622344
rect 342904 616140 342956 616146
rect 342904 616082 342956 616088
rect 234620 610292 234672 610298
rect 234620 610234 234672 610240
rect 356716 607918 356744 622338
rect 360844 616140 360896 616146
rect 360844 616082 360896 616088
rect 356704 607912 356756 607918
rect 356704 607854 356756 607860
rect 233884 603152 233936 603158
rect 233884 603094 233936 603100
rect 232596 600976 232648 600982
rect 232596 600918 232648 600924
rect 360856 594454 360884 616082
rect 369124 607912 369176 607918
rect 369124 607854 369176 607860
rect 360844 594448 360896 594454
rect 360844 594390 360896 594396
rect 366364 594448 366416 594454
rect 366364 594390 366416 594396
rect 366376 574122 366404 594390
rect 369136 590646 369164 607854
rect 369124 590640 369176 590646
rect 369124 590582 369176 590588
rect 371884 590640 371936 590646
rect 371884 590582 371936 590588
rect 371896 585818 371924 590582
rect 371884 585812 371936 585818
rect 371884 585754 371936 585760
rect 380164 585812 380216 585818
rect 380164 585754 380216 585760
rect 366364 574116 366416 574122
rect 366364 574058 366416 574064
rect 369124 574116 369176 574122
rect 369124 574058 369176 574064
rect 231124 572756 231176 572762
rect 231124 572698 231176 572704
rect 232504 572756 232556 572762
rect 232504 572698 232556 572704
rect 209044 565004 209096 565010
rect 209044 564946 209096 564952
rect 211804 565004 211856 565010
rect 211804 564946 211856 564952
rect 189080 560992 189132 560998
rect 189080 560934 189132 560940
rect 202144 560992 202196 560998
rect 202144 560934 202196 560940
rect 189092 559026 189120 560934
rect 184940 559020 184992 559026
rect 184940 558962 184992 558968
rect 189080 559020 189132 559026
rect 189080 558962 189132 558968
rect 184952 554826 184980 558962
rect 209056 556238 209084 564946
rect 231136 564738 231164 572698
rect 229928 564732 229980 564738
rect 229928 564674 229980 564680
rect 231124 564732 231176 564738
rect 231124 564674 231176 564680
rect 229940 562698 229968 564674
rect 228364 562692 228416 562698
rect 228364 562634 228416 562640
rect 229928 562692 229980 562698
rect 229928 562634 229980 562640
rect 201224 556232 201276 556238
rect 201224 556174 201276 556180
rect 209044 556232 209096 556238
rect 209044 556174 209096 556180
rect 184860 554798 184980 554826
rect 181444 554056 181496 554062
rect 181444 553998 181496 554004
rect 184860 552702 184888 554798
rect 201236 552906 201264 556174
rect 193864 552900 193916 552906
rect 193864 552842 193916 552848
rect 201224 552900 201276 552906
rect 201224 552842 201276 552848
rect 183192 552696 183244 552702
rect 183192 552638 183244 552644
rect 184848 552696 184900 552702
rect 184848 552638 184900 552644
rect 183204 550458 183232 552638
rect 181444 550452 181496 550458
rect 181444 550394 181496 550400
rect 183192 550452 183244 550458
rect 183192 550394 183244 550400
rect 170404 545760 170456 545766
rect 170404 545702 170456 545708
rect 170416 537538 170444 545702
rect 170404 537532 170456 537538
rect 170404 537474 170456 537480
rect 181456 534070 181484 550394
rect 193876 545766 193904 552842
rect 228376 552702 228404 562634
rect 226984 552696 227036 552702
rect 226984 552638 227036 552644
rect 228364 552696 228416 552702
rect 228364 552638 228416 552644
rect 226996 546514 227024 552638
rect 224960 546508 225012 546514
rect 224960 546450 225012 546456
rect 226984 546508 227036 546514
rect 226984 546450 227036 546456
rect 193864 545760 193916 545766
rect 193864 545702 193916 545708
rect 224972 542450 225000 546450
rect 224880 542422 225000 542450
rect 224880 540122 224908 542422
rect 223028 540116 223080 540122
rect 223028 540058 223080 540064
rect 224868 540116 224920 540122
rect 224868 540058 224920 540064
rect 223040 535498 223068 540058
rect 220360 535492 220412 535498
rect 220360 535434 220412 535440
rect 223028 535492 223080 535498
rect 223028 535434 223080 535440
rect 180064 534064 180116 534070
rect 180064 534006 180116 534012
rect 181444 534064 181496 534070
rect 181444 534006 181496 534012
rect 180076 505170 180104 534006
rect 220372 532370 220400 535434
rect 218704 532364 218756 532370
rect 218704 532306 218756 532312
rect 220360 532364 220412 532370
rect 220360 532306 220412 532312
rect 178684 505164 178736 505170
rect 178684 505106 178736 505112
rect 180064 505164 180116 505170
rect 180064 505106 180116 505112
rect 178696 498234 178724 505106
rect 175280 498228 175332 498234
rect 175280 498170 175332 498176
rect 178684 498228 178736 498234
rect 178684 498170 178736 498176
rect 175292 495530 175320 498170
rect 175200 495502 175320 495530
rect 175200 493338 175228 495502
rect 218716 493338 218744 532306
rect 173164 493332 173216 493338
rect 173164 493274 173216 493280
rect 175188 493332 175240 493338
rect 175188 493274 175240 493280
rect 217324 493332 217376 493338
rect 217324 493274 217376 493280
rect 218704 493332 218756 493338
rect 218704 493274 218756 493280
rect 173176 482866 173204 493274
rect 171140 482860 171192 482866
rect 171140 482802 171192 482808
rect 173164 482860 173216 482866
rect 173164 482802 173216 482808
rect 171152 478922 171180 482802
rect 217336 482730 217364 493274
rect 369136 490414 369164 574058
rect 380176 570654 380204 585754
rect 380164 570648 380216 570654
rect 380164 570590 380216 570596
rect 392584 570648 392636 570654
rect 392584 570590 392636 570596
rect 392596 564398 392624 570590
rect 392584 564392 392636 564398
rect 392584 564334 392636 564340
rect 369124 490408 369176 490414
rect 369124 490350 369176 490356
rect 376024 490408 376076 490414
rect 376024 490350 376076 490356
rect 215944 482724 215996 482730
rect 215944 482666 215996 482672
rect 217324 482724 217376 482730
rect 217324 482666 217376 482672
rect 171140 478916 171192 478922
rect 171140 478858 171192 478864
rect 215956 469266 215984 482666
rect 213184 469260 213236 469266
rect 213184 469202 213236 469208
rect 215944 469260 215996 469266
rect 215944 469202 215996 469208
rect 213196 454102 213224 469202
rect 376036 456074 376064 490350
rect 376024 456068 376076 456074
rect 376024 456010 376076 456016
rect 385684 456068 385736 456074
rect 385684 456010 385736 456016
rect 213184 454096 213236 454102
rect 213184 454038 213236 454044
rect 210516 454028 210568 454034
rect 210516 453970 210568 453976
rect 210528 446418 210556 453970
rect 209044 446412 209096 446418
rect 209044 446354 209096 446360
rect 210516 446412 210568 446418
rect 210516 446354 210568 446360
rect 209056 438938 209084 446354
rect 207664 438932 207716 438938
rect 207664 438874 207716 438880
rect 209044 438932 209096 438938
rect 209044 438874 209096 438880
rect 207676 430642 207704 438874
rect 204904 430636 204956 430642
rect 204904 430578 204956 430584
rect 207664 430636 207716 430642
rect 207664 430578 207716 430584
rect 204916 388482 204944 430578
rect 385696 388550 385724 456010
rect 385684 388544 385736 388550
rect 385684 388486 385736 388492
rect 389272 388544 389324 388550
rect 389272 388486 389324 388492
rect 199384 388476 199436 388482
rect 199384 388418 199436 388424
rect 204904 388476 204956 388482
rect 204904 388418 204956 388424
rect 199396 372638 199424 388418
rect 389284 385014 389312 388486
rect 389272 385008 389324 385014
rect 389272 384950 389324 384956
rect 392768 385008 392820 385014
rect 392768 384950 392820 384956
rect 392780 382226 392808 384950
rect 392768 382220 392820 382226
rect 392768 382162 392820 382168
rect 197360 372632 197412 372638
rect 197360 372574 197412 372580
rect 199384 372632 199436 372638
rect 199384 372574 199436 372580
rect 197372 369918 197400 372574
rect 197360 369912 197412 369918
rect 197360 369854 197412 369860
rect 192484 369844 192536 369850
rect 192484 369786 192536 369792
rect 192496 345098 192524 369786
rect 189724 345092 189776 345098
rect 189724 345034 189776 345040
rect 192484 345092 192536 345098
rect 192484 345034 192536 345040
rect 189736 336802 189764 345034
rect 189724 336796 189776 336802
rect 189724 336738 189776 336744
rect 186228 336728 186280 336734
rect 186228 336670 186280 336676
rect 186240 330070 186268 336670
rect 183560 330064 183612 330070
rect 183560 330006 183612 330012
rect 186228 330064 186280 330070
rect 186228 330006 186280 330012
rect 183572 326466 183600 330006
rect 182824 326460 182876 326466
rect 182824 326402 182876 326408
rect 183560 326460 183612 326466
rect 183560 326402 183612 326408
rect 182836 306406 182864 326402
rect 179604 306400 179656 306406
rect 179604 306342 179656 306348
rect 182824 306400 182876 306406
rect 182824 306342 182876 306348
rect 179616 301442 179644 306342
rect 178684 301436 178736 301442
rect 178684 301378 178736 301384
rect 179604 301436 179656 301442
rect 179604 301378 179656 301384
rect 178696 294030 178724 301378
rect 175280 294024 175332 294030
rect 175280 293966 175332 293972
rect 178684 294024 178736 294030
rect 178684 293966 178736 293972
rect 175292 289762 175320 293966
rect 174924 289734 175320 289762
rect 174924 281858 174952 289734
rect 173164 281852 173216 281858
rect 173164 281794 173216 281800
rect 174912 281852 174964 281858
rect 174912 281794 174964 281800
rect 169760 280832 169812 280838
rect 169760 280774 169812 280780
rect 124864 273284 124916 273290
rect 124864 273226 124916 273232
rect 118700 273216 118752 273222
rect 118700 273158 118752 273164
rect 118712 270570 118740 273158
rect 173176 271862 173204 281794
rect 167644 271856 167696 271862
rect 167644 271798 167696 271804
rect 173164 271856 173216 271862
rect 173164 271798 173216 271804
rect 116768 270564 116820 270570
rect 116768 270506 116820 270512
rect 118700 270564 118752 270570
rect 118700 270506 118752 270512
rect 116780 268394 116808 270506
rect 112168 268388 112220 268394
rect 112168 268330 112220 268336
rect 116768 268388 116820 268394
rect 116768 268330 116820 268336
rect 112180 266422 112208 268330
rect 167656 266626 167684 271798
rect 165620 266620 165672 266626
rect 165620 266562 165672 266568
rect 167644 266620 167696 266626
rect 167644 266562 167696 266568
rect 54208 266416 54260 266422
rect 54208 266358 54260 266364
rect 55956 266416 56008 266422
rect 55956 266358 56008 266364
rect 109040 266416 109092 266422
rect 109040 266358 109092 266364
rect 112168 266416 112220 266422
rect 112168 266358 112220 266364
rect 54220 263634 54248 266358
rect 53288 263628 53340 263634
rect 53288 263570 53340 263576
rect 54208 263628 54260 263634
rect 54208 263570 54260 263576
rect 53300 256766 53328 263570
rect 109052 262290 109080 266358
rect 165632 265674 165660 266562
rect 158720 265668 158772 265674
rect 158720 265610 158772 265616
rect 165620 265668 165672 265674
rect 165620 265610 165672 265616
rect 108960 262262 109080 262290
rect 108960 260506 108988 262262
rect 107016 260500 107068 260506
rect 107016 260442 107068 260448
rect 108948 260500 109000 260506
rect 108948 260442 109000 260448
rect 107028 256766 107056 260442
rect 158732 259282 158760 265610
rect 151820 259276 151872 259282
rect 151820 259218 151872 259224
rect 158720 259276 158772 259282
rect 158720 259218 158772 259224
rect 53288 256760 53340 256766
rect 53288 256702 53340 256708
rect 104900 256760 104952 256766
rect 104900 256702 104952 256708
rect 107016 256760 107068 256766
rect 151832 256714 151860 259218
rect 107016 256702 107068 256708
rect 104912 255338 104940 256702
rect 151740 256686 151860 256714
rect 104900 255332 104952 255338
rect 104900 255274 104952 255280
rect 101404 255264 101456 255270
rect 101404 255206 101456 255212
rect 53196 254040 53248 254046
rect 53196 253982 53248 253988
rect 51080 252884 51132 252890
rect 51080 252826 51132 252832
rect 53104 252884 53156 252890
rect 53104 252826 53156 252832
rect 51092 250442 51120 252826
rect 50344 250436 50396 250442
rect 50344 250378 50396 250384
rect 51080 250436 51132 250442
rect 51080 250378 51132 250384
rect 47584 245676 47636 245682
rect 47584 245618 47636 245624
rect 46204 244996 46256 245002
rect 46204 244938 46256 244944
rect 50356 240582 50384 250378
rect 101416 240854 101444 255206
rect 151740 253978 151768 256686
rect 151728 253972 151780 253978
rect 151728 253914 151780 253920
rect 146944 253904 146996 253910
rect 146944 253846 146996 253852
rect 146956 247110 146984 253846
rect 143264 247104 143316 247110
rect 143264 247046 143316 247052
rect 146944 247104 146996 247110
rect 146944 247046 146996 247052
rect 101404 240848 101456 240854
rect 101404 240790 101456 240796
rect 143276 240786 143304 247046
rect 143264 240780 143316 240786
rect 143264 240722 143316 240728
rect 50344 240576 50396 240582
rect 50344 240518 50396 240524
rect 395356 239834 395384 652258
rect 395436 564392 395488 564398
rect 395436 564334 395488 564340
rect 395448 240106 395476 564334
rect 395528 382220 395580 382226
rect 395528 382162 395580 382168
rect 395540 343670 395568 382162
rect 395528 343664 395580 343670
rect 395528 343606 395580 343612
rect 395436 240100 395488 240106
rect 395436 240042 395488 240048
rect 395344 239828 395396 239834
rect 395344 239770 395396 239776
rect 45836 238808 45888 238814
rect 45836 238750 45888 238756
rect 45744 233368 45796 233374
rect 45744 233310 45796 233316
rect 45836 233164 45888 233170
rect 45836 233106 45888 233112
rect 45744 232824 45796 232830
rect 45744 232766 45796 232772
rect 45756 230450 45784 232766
rect 45848 231198 45876 233106
rect 62764 232416 62816 232422
rect 62764 232358 62816 232364
rect 82084 232416 82136 232422
rect 82084 232358 82136 232364
rect 395436 232416 395488 232422
rect 395436 232358 395488 232364
rect 45836 231192 45888 231198
rect 45836 231134 45888 231140
rect 47676 230580 47728 230586
rect 47676 230522 47728 230528
rect 45744 230444 45796 230450
rect 45744 230386 45796 230392
rect 47584 230444 47636 230450
rect 47584 230386 47636 230392
rect 47596 222154 47624 230386
rect 47584 222148 47636 222154
rect 47584 222090 47636 222096
rect 45572 219406 45692 219434
rect 45284 217660 45336 217666
rect 45284 217602 45336 217608
rect 45572 207670 45600 219406
rect 47584 217660 47636 217666
rect 47584 217602 47636 217608
rect 45560 207664 45612 207670
rect 45560 207606 45612 207612
rect 47596 194546 47624 217602
rect 47688 216782 47716 230522
rect 55128 230376 55180 230382
rect 55128 230318 55180 230324
rect 55140 228970 55168 230318
rect 55140 228942 55260 228970
rect 49976 228404 50028 228410
rect 49976 228346 50028 228352
rect 48228 226296 48280 226302
rect 48228 226238 48280 226244
rect 48240 222222 48268 226238
rect 49988 225010 50016 228346
rect 49976 225004 50028 225010
rect 49976 224946 50028 224952
rect 53840 225004 53892 225010
rect 53840 224946 53892 224952
rect 48228 222216 48280 222222
rect 48228 222158 48280 222164
rect 48320 222148 48372 222154
rect 48320 222090 48372 222096
rect 53196 222148 53248 222154
rect 53196 222090 53248 222096
rect 48332 219502 48360 222090
rect 48320 219496 48372 219502
rect 48320 219438 48372 219444
rect 47676 216776 47728 216782
rect 47676 216718 47728 216724
rect 50344 216776 50396 216782
rect 50344 216718 50396 216724
rect 50356 205766 50384 216718
rect 53208 215286 53236 222090
rect 53852 221474 53880 224946
rect 55232 224194 55260 228942
rect 55220 224188 55272 224194
rect 55220 224130 55272 224136
rect 53840 221468 53892 221474
rect 53840 221410 53892 221416
rect 55128 219428 55180 219434
rect 55128 219370 55180 219376
rect 53196 215280 53248 215286
rect 53196 215222 53248 215228
rect 53840 215280 53892 215286
rect 53840 215222 53892 215228
rect 55140 215234 55168 219370
rect 53852 211750 53880 215222
rect 55140 215206 55260 215234
rect 55232 213246 55260 215206
rect 55220 213240 55272 213246
rect 55220 213182 55272 213188
rect 53840 211744 53892 211750
rect 53840 211686 53892 211692
rect 55220 211744 55272 211750
rect 55220 211686 55272 211692
rect 55232 208894 55260 211686
rect 55220 208888 55272 208894
rect 55220 208830 55272 208836
rect 50436 207664 50488 207670
rect 50436 207606 50488 207612
rect 50344 205760 50396 205766
rect 50344 205702 50396 205708
rect 50448 201958 50476 207606
rect 54484 205760 54536 205766
rect 54484 205702 54536 205708
rect 50436 201952 50488 201958
rect 50436 201894 50488 201900
rect 47584 194540 47636 194546
rect 47584 194482 47636 194488
rect 54496 192506 54524 205702
rect 56612 195974 56640 230588
rect 62776 227186 62804 232358
rect 82096 227730 82124 232358
rect 395344 232348 395396 232354
rect 395344 232290 395396 232296
rect 391204 232280 391256 232286
rect 391204 232222 391256 232228
rect 134156 231192 134208 231198
rect 134156 231134 134208 231140
rect 84844 231056 84896 231062
rect 84844 230998 84896 231004
rect 82084 227724 82136 227730
rect 82084 227666 82136 227672
rect 62764 227180 62816 227186
rect 62764 227122 62816 227128
rect 65800 227180 65852 227186
rect 65800 227122 65852 227128
rect 59360 224188 59412 224194
rect 59360 224130 59412 224136
rect 59268 221468 59320 221474
rect 59268 221410 59320 221416
rect 59280 215762 59308 221410
rect 59372 220794 59400 224130
rect 65812 222154 65840 227122
rect 65800 222148 65852 222154
rect 65800 222090 65852 222096
rect 69664 222148 69716 222154
rect 69664 222090 69716 222096
rect 59360 220788 59412 220794
rect 59360 220730 59412 220736
rect 62764 220788 62816 220794
rect 62764 220730 62816 220736
rect 59268 215756 59320 215762
rect 59268 215698 59320 215704
rect 61384 215756 61436 215762
rect 61384 215698 61436 215704
rect 56876 208888 56928 208894
rect 56876 208830 56928 208836
rect 56888 205698 56916 208830
rect 56876 205692 56928 205698
rect 56876 205634 56928 205640
rect 60004 205624 60056 205630
rect 60004 205566 60056 205572
rect 57244 201952 57296 201958
rect 57244 201894 57296 201900
rect 56600 195968 56652 195974
rect 56600 195910 56652 195916
rect 54576 194540 54628 194546
rect 54576 194482 54628 194488
rect 54484 192500 54536 192506
rect 54484 192442 54536 192448
rect 54588 189786 54616 194482
rect 54576 189780 54628 189786
rect 54576 189722 54628 189728
rect 57256 184210 57284 201894
rect 60016 197334 60044 205566
rect 61396 204950 61424 215698
rect 61384 204944 61436 204950
rect 61384 204886 61436 204892
rect 60004 197328 60056 197334
rect 60004 197270 60056 197276
rect 58624 192500 58676 192506
rect 58624 192442 58676 192448
rect 57244 184204 57296 184210
rect 57244 184146 57296 184152
rect 58636 182510 58664 192442
rect 60740 189780 60792 189786
rect 60740 189722 60792 189728
rect 60752 184890 60780 189722
rect 62776 186114 62804 220730
rect 68284 213240 68336 213246
rect 68284 213182 68336 213188
rect 68296 204270 68324 213182
rect 69676 209574 69704 222090
rect 84856 220794 84884 230998
rect 85488 227724 85540 227730
rect 85488 227666 85540 227672
rect 85500 224262 85528 227666
rect 85488 224256 85540 224262
rect 85488 224198 85540 224204
rect 84844 220788 84896 220794
rect 84844 220730 84896 220736
rect 85764 220788 85816 220794
rect 85764 220730 85816 220736
rect 85776 218074 85804 220730
rect 85764 218068 85816 218074
rect 85764 218010 85816 218016
rect 69664 209568 69716 209574
rect 69664 209510 69716 209516
rect 77024 209568 77076 209574
rect 77024 209510 77076 209516
rect 77036 205834 77064 209510
rect 77024 205828 77076 205834
rect 77024 205770 77076 205776
rect 78680 205828 78732 205834
rect 78680 205770 78732 205776
rect 75184 204944 75236 204950
rect 75184 204886 75236 204892
rect 68284 204264 68336 204270
rect 68284 204206 68336 204212
rect 69664 204264 69716 204270
rect 69664 204206 69716 204212
rect 65524 197328 65576 197334
rect 65524 197270 65576 197276
rect 62764 186108 62816 186114
rect 62764 186050 62816 186056
rect 64144 186108 64196 186114
rect 64144 186050 64196 186056
rect 60740 184884 60792 184890
rect 60740 184826 60792 184832
rect 58624 182504 58676 182510
rect 58624 182446 58676 182452
rect 64156 159390 64184 186050
rect 64880 182504 64932 182510
rect 64880 182446 64932 182452
rect 64892 177206 64920 182446
rect 65536 179926 65564 197270
rect 69676 186386 69704 204206
rect 75196 187814 75224 204886
rect 78692 202162 78720 205770
rect 78680 202156 78732 202162
rect 78680 202098 78732 202104
rect 86972 195906 87000 230588
rect 115952 230574 116518 230602
rect 100024 224256 100076 224262
rect 100024 224198 100076 224204
rect 87604 218068 87656 218074
rect 87604 218010 87656 218016
rect 87616 202842 87644 218010
rect 100036 215966 100064 224198
rect 100024 215960 100076 215966
rect 100024 215902 100076 215908
rect 111064 215960 111116 215966
rect 111064 215902 111116 215908
rect 87604 202836 87656 202842
rect 87604 202778 87656 202784
rect 93124 202836 93176 202842
rect 93124 202778 93176 202784
rect 88064 202156 88116 202162
rect 88064 202098 88116 202104
rect 88076 198762 88104 202098
rect 88064 198756 88116 198762
rect 88064 198698 88116 198704
rect 90364 198756 90416 198762
rect 90364 198698 90416 198704
rect 86960 195900 87012 195906
rect 86960 195842 87012 195848
rect 75184 187808 75236 187814
rect 75184 187750 75236 187756
rect 80060 187808 80112 187814
rect 80060 187750 80112 187756
rect 69664 186380 69716 186386
rect 69664 186322 69716 186328
rect 71136 186380 71188 186386
rect 71136 186322 71188 186328
rect 65616 184884 65668 184890
rect 65616 184826 65668 184832
rect 65524 179920 65576 179926
rect 65524 179862 65576 179868
rect 64880 177200 64932 177206
rect 64880 177142 64932 177148
rect 65628 172446 65656 184826
rect 65800 184204 65852 184210
rect 65800 184146 65852 184152
rect 65812 180606 65840 184146
rect 71148 183530 71176 186322
rect 71136 183524 71188 183530
rect 71136 183466 71188 183472
rect 72516 183524 72568 183530
rect 72516 183466 72568 183472
rect 65800 180600 65852 180606
rect 65800 180542 65852 180548
rect 68376 180600 68428 180606
rect 68376 180542 68428 180548
rect 66996 179920 67048 179926
rect 66996 179862 67048 179868
rect 67008 172514 67036 179862
rect 66996 172508 67048 172514
rect 66996 172450 67048 172456
rect 68284 172508 68336 172514
rect 68284 172450 68336 172456
rect 65616 172440 65668 172446
rect 65616 172382 65668 172388
rect 64144 159384 64196 159390
rect 64144 159326 64196 159332
rect 66168 159384 66220 159390
rect 66168 159326 66220 159332
rect 66180 151814 66208 159326
rect 66180 151786 66300 151814
rect 66272 151502 66300 151786
rect 66260 151496 66312 151502
rect 66260 151438 66312 151444
rect 62764 139528 62816 139534
rect 62764 139470 62816 139476
rect 43444 122800 43496 122806
rect 43444 122742 43496 122748
rect 37924 121440 37976 121446
rect 37924 121382 37976 121388
rect 23480 117292 23532 117298
rect 23480 117234 23532 117240
rect 62776 111790 62804 139470
rect 68296 132190 68324 172450
rect 68388 167006 68416 180542
rect 72528 178090 72556 183466
rect 80072 182850 80100 187750
rect 80060 182844 80112 182850
rect 80060 182786 80112 182792
rect 88984 182844 89036 182850
rect 88984 182786 89036 182792
rect 72516 178084 72568 178090
rect 72516 178026 72568 178032
rect 73804 178084 73856 178090
rect 73804 178026 73856 178032
rect 68468 177200 68520 177206
rect 68468 177142 68520 177148
rect 68480 168094 68508 177142
rect 71044 172440 71096 172446
rect 71044 172382 71096 172388
rect 68468 168088 68520 168094
rect 68468 168030 68520 168036
rect 68376 167000 68428 167006
rect 68376 166942 68428 166948
rect 71056 154562 71084 172382
rect 71504 168088 71556 168094
rect 71504 168030 71556 168036
rect 71516 163606 71544 168030
rect 71780 167000 71832 167006
rect 71780 166942 71832 166948
rect 71504 163600 71556 163606
rect 71504 163542 71556 163548
rect 71792 163538 71820 166942
rect 71780 163532 71832 163538
rect 71780 163474 71832 163480
rect 73816 160138 73844 178026
rect 82820 163600 82872 163606
rect 82820 163542 82872 163548
rect 73804 160132 73856 160138
rect 73804 160074 73856 160080
rect 76564 160064 76616 160070
rect 76564 160006 76616 160012
rect 71044 154556 71096 154562
rect 71044 154498 71096 154504
rect 74172 154556 74224 154562
rect 74172 154498 74224 154504
rect 68376 151496 68428 151502
rect 68376 151438 68428 151444
rect 68284 132184 68336 132190
rect 68284 132126 68336 132132
rect 68388 129062 68416 151438
rect 74184 145586 74212 154498
rect 76576 147626 76604 160006
rect 82832 159118 82860 163542
rect 86224 163532 86276 163538
rect 86224 163474 86276 163480
rect 82820 159112 82872 159118
rect 82820 159054 82872 159060
rect 86236 147966 86264 163474
rect 86592 159112 86644 159118
rect 86592 159054 86644 159060
rect 86604 153202 86632 159054
rect 88996 158710 89024 182786
rect 90376 181490 90404 198698
rect 93136 189310 93164 202778
rect 111076 202162 111104 215902
rect 111064 202156 111116 202162
rect 111064 202098 111116 202104
rect 115952 194614 115980 230574
rect 134168 230110 134196 231134
rect 180800 231124 180852 231130
rect 180800 231066 180852 231072
rect 146312 230574 146510 230602
rect 134156 230104 134208 230110
rect 134156 230046 134208 230052
rect 136364 230104 136416 230110
rect 136364 230046 136416 230052
rect 136376 225214 136404 230046
rect 138664 227792 138716 227798
rect 138664 227734 138716 227740
rect 136364 225208 136416 225214
rect 136364 225150 136416 225156
rect 118700 222896 118752 222902
rect 118700 222838 118752 222844
rect 118608 218068 118660 218074
rect 118608 218010 118660 218016
rect 115940 194608 115992 194614
rect 115940 194550 115992 194556
rect 93124 189304 93176 189310
rect 93124 189246 93176 189252
rect 94504 189304 94556 189310
rect 94504 189246 94556 189252
rect 94516 184890 94544 189246
rect 94504 184884 94556 184890
rect 94504 184826 94556 184832
rect 97264 184884 97316 184890
rect 97264 184826 97316 184832
rect 90364 181484 90416 181490
rect 90364 181426 90416 181432
rect 97276 165578 97304 184826
rect 100024 181484 100076 181490
rect 100024 181426 100076 181432
rect 97264 165572 97316 165578
rect 97264 165514 97316 165520
rect 98644 165572 98696 165578
rect 98644 165514 98696 165520
rect 88984 158704 89036 158710
rect 88984 158646 89036 158652
rect 96528 158704 96580 158710
rect 96528 158646 96580 158652
rect 96540 153882 96568 158646
rect 96528 153876 96580 153882
rect 96528 153818 96580 153824
rect 86592 153196 86644 153202
rect 86592 153138 86644 153144
rect 89628 153196 89680 153202
rect 89628 153138 89680 153144
rect 86224 147960 86276 147966
rect 86224 147902 86276 147908
rect 88984 147960 89036 147966
rect 88984 147902 89036 147908
rect 76564 147620 76616 147626
rect 76564 147562 76616 147568
rect 79968 147620 80020 147626
rect 79968 147562 80020 147568
rect 74172 145580 74224 145586
rect 74172 145522 74224 145528
rect 78680 145580 78732 145586
rect 78680 145522 78732 145528
rect 78692 143546 78720 145522
rect 79980 143614 80008 147562
rect 79968 143608 80020 143614
rect 79968 143550 80020 143556
rect 78680 143540 78732 143546
rect 78680 143482 78732 143488
rect 82084 143540 82136 143546
rect 82084 143482 82136 143488
rect 84200 143540 84252 143546
rect 84200 143482 84252 143488
rect 69020 132184 69072 132190
rect 69020 132126 69072 132132
rect 69032 131034 69060 132126
rect 69020 131028 69072 131034
rect 69020 130970 69072 130976
rect 74908 131028 74960 131034
rect 74908 130970 74960 130976
rect 74920 129062 74948 130970
rect 68376 129056 68428 129062
rect 68376 128998 68428 129004
rect 69664 129056 69716 129062
rect 69664 128998 69716 129004
rect 74908 129056 74960 129062
rect 74908 128998 74960 129004
rect 69676 120902 69704 128998
rect 82096 123486 82124 143482
rect 84212 137358 84240 143482
rect 88996 138718 89024 147902
rect 89640 146946 89668 153138
rect 89628 146940 89680 146946
rect 89628 146882 89680 146888
rect 98656 139670 98684 165514
rect 98644 139664 98696 139670
rect 98644 139606 98696 139612
rect 88984 138712 89036 138718
rect 88984 138654 89036 138660
rect 97264 138712 97316 138718
rect 97264 138654 97316 138660
rect 84200 137352 84252 137358
rect 84200 137294 84252 137300
rect 87604 137352 87656 137358
rect 87604 137294 87656 137300
rect 87616 129810 87644 137294
rect 87604 129804 87656 129810
rect 87604 129746 87656 129752
rect 90364 129804 90416 129810
rect 90364 129746 90416 129752
rect 84844 129056 84896 129062
rect 84844 128998 84896 129004
rect 82084 123480 82136 123486
rect 82084 123422 82136 123428
rect 69664 120896 69716 120902
rect 69664 120838 69716 120844
rect 71688 120896 71740 120902
rect 71688 120838 71740 120844
rect 71700 119950 71728 120838
rect 71688 119944 71740 119950
rect 71688 119886 71740 119892
rect 73160 119944 73212 119950
rect 73160 119886 73212 119892
rect 73172 114918 73200 119886
rect 73160 114912 73212 114918
rect 73160 114854 73212 114860
rect 74908 114912 74960 114918
rect 74908 114854 74960 114860
rect 74920 111858 74948 114854
rect 84856 113150 84884 128998
rect 84844 113144 84896 113150
rect 84844 113086 84896 113092
rect 90376 112198 90404 129746
rect 97276 124098 97304 138654
rect 97264 124092 97316 124098
rect 97264 124034 97316 124040
rect 90456 123480 90508 123486
rect 90456 123422 90508 123428
rect 90364 112192 90416 112198
rect 90364 112134 90416 112140
rect 74908 111852 74960 111858
rect 74908 111794 74960 111800
rect 62764 111784 62816 111790
rect 62764 111726 62816 111732
rect 90468 110566 90496 123422
rect 100036 122126 100064 181426
rect 118424 169040 118476 169046
rect 118424 168982 118476 168988
rect 109684 153876 109736 153882
rect 109684 153818 109736 153824
rect 106004 146940 106056 146946
rect 106004 146882 106056 146888
rect 106016 144634 106044 146882
rect 106004 144628 106056 144634
rect 106004 144570 106056 144576
rect 109696 140214 109724 153818
rect 109776 144628 109828 144634
rect 109776 144570 109828 144576
rect 109684 140208 109736 140214
rect 109684 140150 109736 140156
rect 100852 139664 100904 139670
rect 100852 139606 100904 139612
rect 100864 135250 100892 139606
rect 100852 135244 100904 135250
rect 100852 135186 100904 135192
rect 102876 135244 102928 135250
rect 102876 135186 102928 135192
rect 102888 129674 102916 135186
rect 109788 131782 109816 144570
rect 118056 144288 118108 144294
rect 118056 144230 118108 144236
rect 117318 136912 117374 136921
rect 117318 136847 117374 136856
rect 116584 136740 116636 136746
rect 116584 136682 116636 136688
rect 109776 131776 109828 131782
rect 109776 131718 109828 131724
rect 102876 129668 102928 129674
rect 102876 129610 102928 129616
rect 104164 129668 104216 129674
rect 104164 129610 104216 129616
rect 100116 124092 100168 124098
rect 100116 124034 100168 124040
rect 100024 122120 100076 122126
rect 100024 122062 100076 122068
rect 100128 113830 100156 124034
rect 104176 118590 104204 129610
rect 110420 122120 110472 122126
rect 110420 122062 110472 122068
rect 110432 120018 110460 122062
rect 110420 120012 110472 120018
rect 110420 119954 110472 119960
rect 114468 120012 114520 120018
rect 114468 119954 114520 119960
rect 104164 118584 104216 118590
rect 104164 118526 104216 118532
rect 108304 118584 108356 118590
rect 108304 118526 108356 118532
rect 100116 113824 100168 113830
rect 100116 113766 100168 113772
rect 91836 112192 91888 112198
rect 91836 112134 91888 112140
rect 91848 111110 91876 112134
rect 91836 111104 91888 111110
rect 91836 111046 91888 111052
rect 97908 111104 97960 111110
rect 97908 111046 97960 111052
rect 90456 110560 90508 110566
rect 90456 110502 90508 110508
rect 93124 110560 93176 110566
rect 93124 110502 93176 110508
rect 93136 101454 93164 110502
rect 97920 110430 97948 111046
rect 97908 110424 97960 110430
rect 97908 110366 97960 110372
rect 108316 108322 108344 118526
rect 114480 114510 114508 119954
rect 114468 114504 114520 114510
rect 114468 114446 114520 114452
rect 111800 113824 111852 113830
rect 111800 113766 111852 113772
rect 108304 108316 108356 108322
rect 108304 108258 108356 108264
rect 109776 108316 109828 108322
rect 109776 108258 109828 108264
rect 109788 104854 109816 108258
rect 111812 106962 111840 113766
rect 111800 106956 111852 106962
rect 111800 106898 111852 106904
rect 109776 104848 109828 104854
rect 109776 104790 109828 104796
rect 111156 104848 111208 104854
rect 111156 104790 111208 104796
rect 93124 101448 93176 101454
rect 93124 101390 93176 101396
rect 102140 101448 102192 101454
rect 102140 101390 102192 101396
rect 102152 99346 102180 101390
rect 102140 99340 102192 99346
rect 102140 99282 102192 99288
rect 105544 99340 105596 99346
rect 105544 99282 105596 99288
rect 105556 86290 105584 99282
rect 111168 97986 111196 104790
rect 111156 97980 111208 97986
rect 111156 97922 111208 97928
rect 112444 97980 112496 97986
rect 112444 97922 112496 97928
rect 112456 92274 112484 97922
rect 112444 92268 112496 92274
rect 112444 92210 112496 92216
rect 113916 92268 113968 92274
rect 113916 92210 113968 92216
rect 113928 86970 113956 92210
rect 113916 86964 113968 86970
rect 113916 86906 113968 86912
rect 105544 86284 105596 86290
rect 105544 86226 105596 86232
rect 6918 79520 6974 79529
rect 116596 79490 116624 136682
rect 117332 136678 117360 136847
rect 117320 136672 117372 136678
rect 117320 136614 117372 136620
rect 117318 135416 117374 135425
rect 117318 135351 117374 135360
rect 117332 135318 117360 135351
rect 117320 135312 117372 135318
rect 117320 135254 117372 135260
rect 117320 133952 117372 133958
rect 117318 133920 117320 133929
rect 117372 133920 117374 133929
rect 117318 133855 117374 133864
rect 117320 132456 117372 132462
rect 117318 132424 117320 132433
rect 117372 132424 117374 132433
rect 117318 132359 117374 132368
rect 117964 131776 118016 131782
rect 117964 131718 118016 131724
rect 117320 131096 117372 131102
rect 117320 131038 117372 131044
rect 117332 130937 117360 131038
rect 117318 130928 117374 130937
rect 117318 130863 117374 130872
rect 117320 129736 117372 129742
rect 117320 129678 117372 129684
rect 117332 129441 117360 129678
rect 117318 129432 117374 129441
rect 117318 129367 117374 129376
rect 117320 128308 117372 128314
rect 117320 128250 117372 128256
rect 117332 127945 117360 128250
rect 117318 127936 117374 127945
rect 117318 127871 117374 127880
rect 117320 126948 117372 126954
rect 117320 126890 117372 126896
rect 117332 126449 117360 126890
rect 117318 126440 117374 126449
rect 117318 126375 117374 126384
rect 117320 125588 117372 125594
rect 117320 125530 117372 125536
rect 117332 124953 117360 125530
rect 117318 124944 117374 124953
rect 117318 124879 117374 124888
rect 117320 124160 117372 124166
rect 117320 124102 117372 124108
rect 117332 123457 117360 124102
rect 117318 123448 117374 123457
rect 117318 123383 117374 123392
rect 117320 122800 117372 122806
rect 117320 122742 117372 122748
rect 117332 121961 117360 122742
rect 117318 121952 117374 121961
rect 117318 121887 117374 121896
rect 117320 121440 117372 121446
rect 117320 121382 117372 121388
rect 117332 120465 117360 121382
rect 117318 120456 117374 120465
rect 117318 120391 117374 120400
rect 117320 120080 117372 120086
rect 117320 120022 117372 120028
rect 117332 118969 117360 120022
rect 117318 118960 117374 118969
rect 117318 118895 117374 118904
rect 117320 118652 117372 118658
rect 117320 118594 117372 118600
rect 117332 117473 117360 118594
rect 117318 117464 117374 117473
rect 117318 117399 117374 117408
rect 117320 117292 117372 117298
rect 117320 117234 117372 117240
rect 117332 115977 117360 117234
rect 117318 115968 117374 115977
rect 117318 115903 117374 115912
rect 117320 114504 117372 114510
rect 117318 114472 117320 114481
rect 117372 114472 117374 114481
rect 117318 114407 117374 114416
rect 117320 113144 117372 113150
rect 117320 113086 117372 113092
rect 117332 112985 117360 113086
rect 117318 112976 117374 112985
rect 117318 112911 117374 112920
rect 117320 111784 117372 111790
rect 117320 111726 117372 111732
rect 117332 111489 117360 111726
rect 117318 111480 117374 111489
rect 117318 111415 117374 111424
rect 117320 110424 117372 110430
rect 117320 110366 117372 110372
rect 117332 109993 117360 110366
rect 117318 109984 117374 109993
rect 117318 109919 117374 109928
rect 117976 99414 118004 131718
rect 117964 99408 118016 99414
rect 117964 99350 118016 99356
rect 118068 95033 118096 144230
rect 118148 142928 118200 142934
rect 118148 142870 118200 142876
rect 118054 95024 118110 95033
rect 118054 94959 118110 94968
rect 118160 92041 118188 142870
rect 118240 142860 118292 142866
rect 118240 142802 118292 142808
rect 118146 92032 118202 92041
rect 118146 91967 118202 91976
rect 118252 90545 118280 142802
rect 118332 139460 118384 139466
rect 118332 139402 118384 139408
rect 118238 90536 118294 90545
rect 118238 90471 118294 90480
rect 116676 86964 116728 86970
rect 116676 86906 116728 86912
rect 116688 82414 116716 86906
rect 118344 86057 118372 139402
rect 118436 108497 118464 168982
rect 118516 148368 118568 148374
rect 118516 148310 118568 148316
rect 118422 108488 118478 108497
rect 118422 108423 118478 108432
rect 118528 87553 118556 148310
rect 118620 89049 118648 218010
rect 118712 93537 118740 222838
rect 126888 202156 126940 202162
rect 126888 202098 126940 202104
rect 126900 196382 126928 202098
rect 138676 196790 138704 227734
rect 138756 225208 138808 225214
rect 138756 225150 138808 225156
rect 138768 218754 138796 225150
rect 138756 218748 138808 218754
rect 138756 218690 138808 218696
rect 146312 197418 146340 230574
rect 157984 228404 158036 228410
rect 157984 228346 158036 228352
rect 147772 202156 147824 202162
rect 147772 202098 147824 202104
rect 146142 197390 146340 197418
rect 147784 197404 147812 202098
rect 155960 199436 156012 199442
rect 155960 199378 156012 199384
rect 148968 198008 149020 198014
rect 148968 197950 149020 197956
rect 148980 197404 149008 197950
rect 155972 197470 156000 199378
rect 154488 197464 154540 197470
rect 154146 197412 154488 197418
rect 154146 197406 154540 197412
rect 155960 197464 156012 197470
rect 155960 197406 156012 197412
rect 154146 197390 154528 197406
rect 157996 197334 158024 228346
rect 158720 218748 158772 218754
rect 158720 218690 158772 218696
rect 158732 216034 158760 218690
rect 158720 216028 158772 216034
rect 158720 215970 158772 215976
rect 162768 216028 162820 216034
rect 162768 215970 162820 215976
rect 162780 212906 162808 215970
rect 162768 212900 162820 212906
rect 162768 212842 162820 212848
rect 164884 212900 164936 212906
rect 164884 212842 164936 212848
rect 164896 208418 164924 212842
rect 164884 208412 164936 208418
rect 164884 208354 164936 208360
rect 166264 208412 166316 208418
rect 166264 208354 166316 208360
rect 166276 197402 166304 208354
rect 176672 202162 176700 230588
rect 179420 229764 179472 229770
rect 179420 229706 179472 229712
rect 176660 202156 176712 202162
rect 176660 202098 176712 202104
rect 166264 197396 166316 197402
rect 166264 197338 166316 197344
rect 167644 197396 167696 197402
rect 167644 197338 167696 197344
rect 152740 197328 152792 197334
rect 152582 197276 152740 197282
rect 152582 197270 152792 197276
rect 157984 197328 158036 197334
rect 157984 197270 158036 197276
rect 152582 197254 152780 197270
rect 138664 196784 138716 196790
rect 164240 196784 164292 196790
rect 138664 196726 138716 196732
rect 150926 196722 151216 196738
rect 164240 196726 164292 196732
rect 150926 196716 151228 196722
rect 150926 196710 151176 196716
rect 151176 196658 151228 196664
rect 155960 196648 156012 196654
rect 155802 196596 155960 196602
rect 155802 196590 156012 196596
rect 155802 196574 156000 196590
rect 126888 196376 126940 196382
rect 126888 196318 126940 196324
rect 129004 196376 129056 196382
rect 129004 196318 129056 196324
rect 129016 185638 129044 196318
rect 140424 196030 140530 196058
rect 157366 196030 157656 196058
rect 138112 195968 138164 195974
rect 138110 195936 138112 195945
rect 140424 195945 140452 196030
rect 138164 195936 138166 195945
rect 140410 195936 140466 195945
rect 138110 195871 138166 195880
rect 139400 195900 139452 195906
rect 157628 195906 157656 196030
rect 158824 195937 158852 196044
rect 160100 195968 160152 195974
rect 158810 195928 158866 195937
rect 140410 195871 140466 195880
rect 157616 195900 157668 195906
rect 139400 195842 139452 195848
rect 158810 195863 158866 195872
rect 160098 195936 160100 195945
rect 160152 195936 160154 195945
rect 160098 195871 160154 195880
rect 157616 195842 157668 195848
rect 139412 195537 139440 195842
rect 140778 195664 140834 195673
rect 140778 195599 140834 195608
rect 139398 195528 139454 195537
rect 139398 195463 139454 195472
rect 140792 194614 140820 195599
rect 140780 194608 140832 194614
rect 140780 194550 140832 194556
rect 140870 191856 140926 191865
rect 140870 191791 140926 191800
rect 140778 190904 140834 190913
rect 140778 190839 140834 190848
rect 129004 185632 129056 185638
rect 129004 185574 129056 185580
rect 132408 185632 132460 185638
rect 132408 185574 132460 185580
rect 132420 183326 132448 185574
rect 140792 184249 140820 190839
rect 140884 184385 140912 191791
rect 140962 191584 141018 191593
rect 140962 191519 141018 191528
rect 140870 184376 140926 184385
rect 140870 184311 140926 184320
rect 140778 184240 140834 184249
rect 140778 184175 140834 184184
rect 140976 184113 141004 191519
rect 144458 191040 144514 191049
rect 144302 190998 144458 191026
rect 144458 190975 144514 190984
rect 144736 190528 144788 190534
rect 144394 190476 144736 190482
rect 144394 190470 144788 190476
rect 144394 190454 144776 190470
rect 145012 190324 145064 190330
rect 145012 190266 145064 190272
rect 145024 188970 145052 190266
rect 145852 189774 145958 189802
rect 145852 189009 145880 189774
rect 164252 189652 164280 196726
rect 166172 193860 166224 193866
rect 166172 193802 166224 193808
rect 145838 189000 145894 189009
rect 144736 188964 144788 188970
rect 144736 188906 144788 188912
rect 145012 188964 145064 188970
rect 145838 188935 145894 188944
rect 145012 188906 145064 188912
rect 140962 184104 141018 184113
rect 140962 184039 141018 184048
rect 132408 183320 132460 183326
rect 132408 183262 132460 183268
rect 135904 183320 135956 183326
rect 135904 183262 135956 183268
rect 121460 180124 121512 180130
rect 121460 180066 121512 180072
rect 118792 167680 118844 167686
rect 118792 167622 118844 167628
rect 118804 102513 118832 167622
rect 118884 160744 118936 160750
rect 118884 160686 118936 160692
rect 118790 102504 118846 102513
rect 118790 102439 118846 102448
rect 118896 101017 118924 160686
rect 118976 153876 119028 153882
rect 118976 153818 119028 153824
rect 118882 101008 118938 101017
rect 118882 100943 118938 100952
rect 118988 99521 119016 153818
rect 119252 144220 119304 144226
rect 119252 144162 119304 144168
rect 119160 141500 119212 141506
rect 119160 141442 119212 141448
rect 119068 141432 119120 141438
rect 119068 141374 119120 141380
rect 118974 99512 119030 99521
rect 118974 99447 119030 99456
rect 119080 96529 119108 141374
rect 119172 98025 119200 141442
rect 119264 105505 119292 144162
rect 119344 141636 119396 141642
rect 119344 141578 119396 141584
rect 119356 107001 119384 141578
rect 120724 141568 120776 141574
rect 120724 141510 120776 141516
rect 120736 113174 120764 141510
rect 121472 139890 121500 180066
rect 122840 178696 122892 178702
rect 122840 178638 122892 178644
rect 122852 151814 122880 178638
rect 124220 177336 124272 177342
rect 124220 177278 124272 177284
rect 124232 151814 124260 177278
rect 126980 176112 127032 176118
rect 126980 176054 127032 176060
rect 125600 175976 125652 175982
rect 125600 175918 125652 175924
rect 125612 151814 125640 175918
rect 126992 151814 127020 176054
rect 128360 175228 128412 175234
rect 128360 175170 128412 175176
rect 128372 151814 128400 175170
rect 133880 173936 133932 173942
rect 133880 173878 133932 173884
rect 131120 172576 131172 172582
rect 131120 172518 131172 172524
rect 122852 151786 122972 151814
rect 124232 151786 124536 151814
rect 125612 151786 126100 151814
rect 126992 151786 127664 151814
rect 128372 151786 129228 151814
rect 122944 139890 122972 151786
rect 124508 139890 124536 151786
rect 126072 139890 126100 151786
rect 127636 139890 127664 151786
rect 129200 139890 129228 151786
rect 131132 139890 131160 172518
rect 132500 171148 132552 171154
rect 132500 171090 132552 171096
rect 132512 139890 132540 171090
rect 133892 139890 133920 173878
rect 135916 173194 135944 183262
rect 136376 182158 136758 182186
rect 136376 180130 136404 182158
rect 144642 181112 144698 181121
rect 144578 181070 144642 181098
rect 144642 181047 144698 181056
rect 144748 180985 144776 188906
rect 166184 188034 166212 193802
rect 165646 188020 166212 188034
rect 165632 188006 166212 188020
rect 144920 181008 144972 181014
rect 144734 180976 144790 180985
rect 136468 180934 136758 180962
rect 136364 180124 136416 180130
rect 136364 180066 136416 180072
rect 135996 178900 136048 178906
rect 135996 178842 136048 178848
rect 136008 177342 136036 178842
rect 136468 178702 136496 180934
rect 144734 180911 144790 180920
rect 144872 180976 144920 180985
rect 144928 180950 144972 180956
rect 144928 180934 144960 180950
rect 144872 180911 144928 180920
rect 153936 180804 153988 180810
rect 153936 180746 153988 180752
rect 153948 180690 153976 180746
rect 153948 180674 154436 180690
rect 153948 180668 154448 180674
rect 153948 180662 154396 180668
rect 154396 180610 154448 180616
rect 165632 180130 165660 188006
rect 167656 183530 167684 197338
rect 167644 183524 167696 183530
rect 167644 183466 167696 183472
rect 169116 183524 169168 183530
rect 169116 183466 169168 183472
rect 157800 180124 157852 180130
rect 157800 180066 157852 180072
rect 158628 180124 158680 180130
rect 158628 180066 158680 180072
rect 165620 180124 165672 180130
rect 165620 180066 165672 180072
rect 157812 180033 157840 180066
rect 157798 180024 157854 180033
rect 136560 179982 136758 180010
rect 136560 178906 136588 179982
rect 157798 179959 157854 179968
rect 136548 178900 136600 178906
rect 136548 178842 136600 178848
rect 136744 178786 136772 179044
rect 144090 178936 144146 178945
rect 144090 178871 144146 178880
rect 136560 178758 136772 178786
rect 141606 178800 141662 178809
rect 136456 178696 136508 178702
rect 136456 178638 136508 178644
rect 136560 178514 136588 178758
rect 141606 178735 141662 178744
rect 143078 178800 143134 178809
rect 143078 178735 143134 178744
rect 136192 178486 136588 178514
rect 135996 177336 136048 177342
rect 135996 177278 136048 177284
rect 136192 175982 136220 178486
rect 136284 177942 136758 177970
rect 136284 176118 136312 177942
rect 136376 177126 136758 177154
rect 136272 176112 136324 176118
rect 136272 176054 136324 176060
rect 136180 175976 136232 175982
rect 136180 175918 136232 175924
rect 136376 175234 136404 177126
rect 136744 175794 136772 175916
rect 136560 175766 136772 175794
rect 136364 175228 136416 175234
rect 136364 175170 136416 175176
rect 135904 173188 135956 173194
rect 135904 173130 135956 173136
rect 136560 172582 136588 175766
rect 136548 172576 136600 172582
rect 136548 172518 136600 172524
rect 135260 171692 135312 171698
rect 135260 171634 135312 171640
rect 135272 151814 135300 171634
rect 136744 171154 136772 174964
rect 141620 174758 141648 178735
rect 143092 174758 143120 178735
rect 144104 175982 144132 178871
rect 149336 176520 149388 176526
rect 158640 176497 158668 180066
rect 159454 180024 159510 180033
rect 159454 179959 159510 179968
rect 159468 177886 159496 179959
rect 166540 178084 166592 178090
rect 166540 178026 166592 178032
rect 159456 177880 159508 177886
rect 159456 177822 159508 177828
rect 149336 176462 149388 176468
rect 158626 176488 158682 176497
rect 149348 175982 149376 176462
rect 153936 176452 153988 176458
rect 154396 176452 154448 176458
rect 153988 176412 154396 176440
rect 153936 176394 153988 176400
rect 158626 176423 158682 176432
rect 154396 176394 154448 176400
rect 144092 175976 144144 175982
rect 144092 175918 144144 175924
rect 149336 175976 149388 175982
rect 149336 175918 149388 175924
rect 162492 175976 162544 175982
rect 162492 175918 162544 175924
rect 144460 175568 144512 175574
rect 144460 175510 144512 175516
rect 149980 175568 150032 175574
rect 149980 175510 150032 175516
rect 141608 174752 141660 174758
rect 141608 174694 141660 174700
rect 143080 174752 143132 174758
rect 143080 174694 143132 174700
rect 137376 173936 137428 173942
rect 137428 173884 137586 173890
rect 137376 173878 137586 173884
rect 137388 173862 137586 173878
rect 138020 172168 138072 172174
rect 138020 172110 138072 172116
rect 136732 171148 136784 171154
rect 136732 171090 136784 171096
rect 138032 151814 138060 172110
rect 138676 171698 138704 173196
rect 139596 173182 139702 173210
rect 138664 171692 138716 171698
rect 138664 171634 138716 171640
rect 135272 151786 135484 151814
rect 138032 151786 138612 151814
rect 135456 139890 135484 151786
rect 137744 143472 137796 143478
rect 137744 143414 137796 143420
rect 137756 139890 137784 143414
rect 121472 139862 121808 139890
rect 122944 139862 123372 139890
rect 124508 139862 124936 139890
rect 126072 139862 126500 139890
rect 127636 139862 128064 139890
rect 129200 139862 129628 139890
rect 131132 139862 131192 139890
rect 132512 139862 132756 139890
rect 133892 139862 134320 139890
rect 135456 139862 135884 139890
rect 137448 139862 137784 139890
rect 138584 139890 138612 151786
rect 139492 146124 139544 146130
rect 139492 146066 139544 146072
rect 139504 140706 139532 146066
rect 139596 143478 139624 173182
rect 140792 172174 140820 173196
rect 140780 172168 140832 172174
rect 140780 172110 140832 172116
rect 141700 146260 141752 146266
rect 141700 146202 141752 146208
rect 139584 143472 139636 143478
rect 139584 143414 139636 143420
rect 139504 140678 140176 140706
rect 140148 139890 140176 140678
rect 141712 139890 141740 146202
rect 142264 146130 142292 173196
rect 142526 172952 142582 172961
rect 142526 172887 142582 172896
rect 142436 166320 142488 166326
rect 142436 166262 142488 166268
rect 142448 146266 142476 166262
rect 142436 146260 142488 146266
rect 142436 146202 142488 146208
rect 142252 146124 142304 146130
rect 142252 146066 142304 146072
rect 142540 143002 142568 172887
rect 142632 166326 142660 173196
rect 142620 166320 142672 166326
rect 142620 166262 142672 166268
rect 143644 161474 143672 173196
rect 143552 161446 143672 161474
rect 142528 142996 142580 143002
rect 142528 142938 142580 142944
rect 143552 139890 143580 161446
rect 144472 143070 144500 175510
rect 149992 175508 150020 175510
rect 154486 175400 154542 175409
rect 154486 175335 154542 175344
rect 152464 174684 152516 174690
rect 152464 174626 152516 174632
rect 152476 174570 152504 174626
rect 152398 174542 152504 174570
rect 144460 143064 144512 143070
rect 144460 143006 144512 143012
rect 144932 139890 144960 173196
rect 146312 151814 146340 173196
rect 146680 161474 146708 173196
rect 148336 172990 148364 173196
rect 149348 172990 149376 173196
rect 148324 172984 148376 172990
rect 148324 172926 148376 172932
rect 149060 172984 149112 172990
rect 149060 172926 149112 172932
rect 149336 172984 149388 172990
rect 149336 172926 149388 172932
rect 148968 172916 149020 172922
rect 148968 172858 149020 172864
rect 148980 170406 149008 172858
rect 148968 170400 149020 170406
rect 148968 170342 149020 170348
rect 146496 161446 146708 161474
rect 146312 151786 146432 151814
rect 146404 139890 146432 151786
rect 146496 143546 146524 161446
rect 146484 143540 146536 143546
rect 146484 143482 146536 143488
rect 148048 143540 148100 143546
rect 148048 143482 148100 143488
rect 148060 139890 148088 143482
rect 149072 142154 149100 172926
rect 149624 161474 149652 173196
rect 150636 161474 150664 173196
rect 151452 172984 151504 172990
rect 151452 172926 151504 172932
rect 149532 161446 149652 161474
rect 150544 161446 150664 161474
rect 149532 142254 149560 161446
rect 150544 143138 150572 161446
rect 150532 143132 150584 143138
rect 150532 143074 150584 143080
rect 149520 142248 149572 142254
rect 149520 142190 149572 142196
rect 149072 142126 149560 142154
rect 149532 139890 149560 142126
rect 151464 139890 151492 172926
rect 152660 161474 152688 173196
rect 152476 161446 152688 161474
rect 153488 173182 153686 173210
rect 152476 143478 152504 161446
rect 153488 143546 153516 173182
rect 154500 158030 154528 175335
rect 156512 174684 156564 174690
rect 156512 174626 156564 174632
rect 154488 158024 154540 158030
rect 154488 157966 154540 157972
rect 153476 143540 153528 143546
rect 153476 143482 153528 143488
rect 152464 143472 152516 143478
rect 152464 143414 152516 143420
rect 154580 143132 154632 143138
rect 154580 143074 154632 143080
rect 152740 142180 152792 142186
rect 152740 142122 152792 142128
rect 152752 139890 152780 142122
rect 154592 139890 154620 143074
rect 156524 139890 156552 174626
rect 161480 174548 161532 174554
rect 161480 174490 161532 174496
rect 157352 142186 157380 173196
rect 158442 172952 158498 172961
rect 158442 172887 158498 172896
rect 158456 169046 158484 172887
rect 158444 169040 158496 169046
rect 158444 168982 158496 168988
rect 161492 151814 161520 174490
rect 162504 172990 162532 175918
rect 162492 172984 162544 172990
rect 162492 172926 162544 172932
rect 162676 170400 162728 170406
rect 162676 170342 162728 170348
rect 162688 167754 162716 170342
rect 162676 167748 162728 167754
rect 162676 167690 162728 167696
rect 161492 151786 162072 151814
rect 158996 143540 159048 143546
rect 158996 143482 159048 143488
rect 157432 143472 157484 143478
rect 157432 143414 157484 143420
rect 157340 142180 157392 142186
rect 157340 142122 157392 142128
rect 138584 139862 139012 139890
rect 140148 139862 140576 139890
rect 141712 139862 142140 139890
rect 143552 139862 143704 139890
rect 144932 139862 145268 139890
rect 146404 139862 146832 139890
rect 148060 139862 148396 139890
rect 149532 139862 149960 139890
rect 151464 139862 151524 139890
rect 152752 139862 153088 139890
rect 154592 139862 154652 139890
rect 156216 139862 156552 139890
rect 157444 139890 157472 143414
rect 159008 139890 159036 143482
rect 160560 143064 160612 143070
rect 160560 143006 160612 143012
rect 160572 139890 160600 143006
rect 162044 139890 162072 151786
rect 163516 143070 163544 175100
rect 163608 143206 163636 173196
rect 164528 173182 164634 173210
rect 163596 143200 163648 143206
rect 163596 143142 163648 143148
rect 164528 143138 164556 173182
rect 165436 172984 165488 172990
rect 165436 172926 165488 172932
rect 164516 143132 164568 143138
rect 164516 143074 164568 143080
rect 163504 143064 163556 143070
rect 163504 143006 163556 143012
rect 163688 142180 163740 142186
rect 163688 142122 163740 142128
rect 163700 139890 163728 142122
rect 165448 139890 165476 172926
rect 166552 161474 166580 178026
rect 167644 177880 167696 177886
rect 167644 177822 167696 177828
rect 167000 174344 167052 174350
rect 167000 174286 167052 174292
rect 166460 161446 166580 161474
rect 165620 158024 165672 158030
rect 165620 157966 165672 157972
rect 165632 154562 165660 157966
rect 165620 154556 165672 154562
rect 165620 154498 165672 154504
rect 166460 148374 166488 161446
rect 166448 148368 166500 148374
rect 166448 148310 166500 148316
rect 167012 139890 167040 174286
rect 167656 143546 167684 177822
rect 169128 176390 169156 183466
rect 169116 176384 169168 176390
rect 169116 176326 169168 176332
rect 169760 176384 169812 176390
rect 169760 176326 169812 176332
rect 169772 171426 169800 176326
rect 169760 171420 169812 171426
rect 169760 171362 169812 171368
rect 171784 171420 171836 171426
rect 171784 171362 171836 171368
rect 168380 154556 168432 154562
rect 168380 154498 168432 154504
rect 167644 143540 167696 143546
rect 167644 143482 167696 143488
rect 168392 139890 168420 154498
rect 171796 147014 171824 171362
rect 172244 167748 172296 167754
rect 172244 167690 172296 167696
rect 172256 164218 172284 167690
rect 172244 164212 172296 164218
rect 172244 164154 172296 164160
rect 175188 164212 175240 164218
rect 175188 164154 175240 164160
rect 175200 158914 175228 164154
rect 175188 158908 175240 158914
rect 175188 158850 175240 158856
rect 177304 158908 177356 158914
rect 177304 158850 177356 158856
rect 171784 147008 171836 147014
rect 171784 146950 171836 146956
rect 172520 147008 172572 147014
rect 172520 146950 172572 146956
rect 172532 143546 172560 146950
rect 177316 144906 177344 158850
rect 177304 144900 177356 144906
rect 177304 144842 177356 144848
rect 169944 143540 169996 143546
rect 169944 143482 169996 143488
rect 172520 143540 172572 143546
rect 172520 143482 172572 143488
rect 176476 143540 176528 143546
rect 176476 143482 176528 143488
rect 169956 139890 169984 143482
rect 174636 143200 174688 143206
rect 174636 143142 174688 143148
rect 173072 142996 173124 143002
rect 173072 142938 173124 142944
rect 171506 142760 171562 142769
rect 171506 142695 171562 142704
rect 171520 139890 171548 142695
rect 173084 139890 173112 142938
rect 174648 139890 174676 143142
rect 176200 143132 176252 143138
rect 176200 143074 176252 143080
rect 176212 139890 176240 143074
rect 176488 141370 176516 143482
rect 178040 143064 178092 143070
rect 178040 143006 178092 143012
rect 176476 141364 176528 141370
rect 176476 141306 176528 141312
rect 178052 139890 178080 143006
rect 157444 139862 157780 139890
rect 159008 139862 159344 139890
rect 160572 139862 160908 139890
rect 162044 139862 162472 139890
rect 163700 139862 164036 139890
rect 165448 139862 165600 139890
rect 167012 139862 167164 139890
rect 168392 139862 168728 139890
rect 169956 139862 170292 139890
rect 171520 139862 171856 139890
rect 173084 139862 173420 139890
rect 174648 139862 174984 139890
rect 176212 139862 176548 139890
rect 178052 139862 178112 139890
rect 179432 122913 179460 229706
rect 179512 213988 179564 213994
rect 179512 213930 179564 213936
rect 179524 132025 179552 213930
rect 180064 191888 180116 191894
rect 180064 191830 180116 191836
rect 179602 135552 179658 135561
rect 179602 135487 179658 135496
rect 179510 132016 179566 132025
rect 179510 131951 179566 131960
rect 179418 122904 179474 122913
rect 179418 122839 179474 122848
rect 120644 113146 120764 113174
rect 119342 106992 119398 107001
rect 119342 106927 119398 106936
rect 119436 106956 119488 106962
rect 119436 106898 119488 106904
rect 119250 105496 119306 105505
rect 119250 105431 119306 105440
rect 119158 98016 119214 98025
rect 119158 97951 119214 97960
rect 119066 96520 119122 96529
rect 119066 96455 119122 96464
rect 118698 93528 118754 93537
rect 118698 93463 118754 93472
rect 118606 89040 118662 89049
rect 118606 88975 118662 88984
rect 118514 87544 118570 87553
rect 118514 87479 118570 87488
rect 118330 86048 118386 86057
rect 118330 85983 118386 85992
rect 118514 83056 118570 83065
rect 118514 82991 118570 83000
rect 116676 82408 116728 82414
rect 116676 82350 116728 82356
rect 118422 81560 118478 81569
rect 118422 81495 118478 81504
rect 6918 79455 6974 79464
rect 116584 79484 116636 79490
rect 116584 79426 116636 79432
rect 5080 78872 5132 78878
rect 5080 78814 5132 78820
rect 89720 78192 89772 78198
rect 89720 78134 89772 78140
rect 46204 78124 46256 78130
rect 46204 78066 46256 78072
rect 22744 77988 22796 77994
rect 22744 77930 22796 77936
rect 20718 76664 20774 76673
rect 20718 76599 20774 76608
rect 6920 75200 6972 75206
rect 6920 75142 6972 75148
rect 4066 58576 4122 58585
rect 4066 58511 4122 58520
rect 3882 19408 3938 19417
rect 3882 19343 3938 19352
rect 4160 18624 4212 18630
rect 4160 18566 4212 18572
rect 4172 16574 4200 18566
rect 6932 16574 6960 75142
rect 19340 42084 19392 42090
rect 19340 42026 19392 42032
rect 19352 16574 19380 42026
rect 20732 16574 20760 76599
rect 22098 43480 22154 43489
rect 22098 43415 22154 43424
rect 22112 16574 22140 43415
rect 4172 16546 5304 16574
rect 6932 16546 7696 16574
rect 19352 16546 19472 16574
rect 20732 16546 21864 16574
rect 22112 16546 22600 16574
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 4066 4856 4122 4865
rect 4066 4791 4122 4800
rect 4080 480 4108 4791
rect 5276 480 5304 16546
rect 6460 4956 6512 4962
rect 6460 4898 6512 4904
rect 6472 480 6500 4898
rect 7668 480 7696 16546
rect 14280 15904 14332 15910
rect 14280 15846 14332 15852
rect 11152 10328 11204 10334
rect 11152 10270 11204 10276
rect 9956 7608 10008 7614
rect 9956 7550 10008 7556
rect 8760 4820 8812 4826
rect 8760 4762 8812 4768
rect 8772 480 8800 4762
rect 9968 480 9996 7550
rect 11164 480 11192 10270
rect 13544 4888 13596 4894
rect 13544 4830 13596 4836
rect 12348 4004 12400 4010
rect 12348 3946 12400 3952
rect 12360 480 12388 3946
rect 13556 480 13584 4830
rect 1646 354 1758 480
rect 1412 326 1758 354
rect 1646 -960 1758 326
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14292 354 14320 15846
rect 18236 6180 18288 6186
rect 18236 6122 18288 6128
rect 15936 5092 15988 5098
rect 15936 5034 15988 5040
rect 15948 480 15976 5034
rect 17040 3528 17092 3534
rect 17040 3470 17092 3476
rect 17052 480 17080 3470
rect 18248 480 18276 6122
rect 19444 480 19472 16546
rect 20626 3360 20682 3369
rect 20626 3295 20682 3304
rect 20640 480 20668 3295
rect 21836 480 21864 16546
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22572 354 22600 16546
rect 22756 4962 22784 77930
rect 44180 76628 44232 76634
rect 44180 76570 44232 76576
rect 30380 76560 30432 76566
rect 30380 76502 30432 76508
rect 27620 73908 27672 73914
rect 27620 73850 27672 73856
rect 26240 73840 26292 73846
rect 26240 73782 26292 73788
rect 25320 6316 25372 6322
rect 25320 6258 25372 6264
rect 22744 4956 22796 4962
rect 22744 4898 22796 4904
rect 24216 4956 24268 4962
rect 24216 4898 24268 4904
rect 24228 480 24256 4898
rect 25332 480 25360 6258
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 73782
rect 27632 16574 27660 73850
rect 30392 16574 30420 76502
rect 35898 75304 35954 75313
rect 35898 75239 35954 75248
rect 42800 75268 42852 75274
rect 34520 44872 34572 44878
rect 34520 44814 34572 44820
rect 31760 18692 31812 18698
rect 31760 18634 31812 18640
rect 31772 16574 31800 18634
rect 27632 16546 27752 16574
rect 30392 16546 30880 16574
rect 31772 16546 31984 16574
rect 27724 480 27752 16546
rect 28448 10396 28500 10402
rect 28448 10338 28500 10344
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28460 354 28488 10338
rect 30104 1148 30156 1154
rect 30104 1090 30156 1096
rect 30116 480 30144 1090
rect 28878 354 28990 480
rect 28460 326 28990 354
rect 28878 -960 28990 326
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31956 354 31984 16546
rect 33600 6248 33652 6254
rect 33600 6190 33652 6196
rect 33232 5024 33284 5030
rect 33232 4966 33284 4972
rect 33244 1154 33272 4966
rect 33232 1148 33284 1154
rect 33232 1090 33284 1096
rect 33612 480 33640 6190
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 31270 -960 31382 326
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34532 354 34560 44814
rect 35912 12434 35940 75239
rect 42800 75210 42852 75216
rect 40038 73808 40094 73817
rect 40038 73743 40094 73752
rect 40052 16574 40080 73743
rect 40052 16546 40264 16574
rect 39120 14476 39172 14482
rect 39120 14418 39172 14424
rect 35912 12406 36860 12434
rect 35992 10464 36044 10470
rect 35992 10406 36044 10412
rect 36004 480 36032 10406
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36832 354 36860 12406
rect 38382 7576 38438 7585
rect 38382 7511 38438 7520
rect 38396 480 38424 7511
rect 37158 354 37270 480
rect 36832 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39132 354 39160 14418
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 40236 354 40264 16546
rect 41878 7712 41934 7721
rect 41878 7647 41934 7656
rect 41892 480 41920 7647
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 39550 -960 39662 326
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 42812 354 42840 75210
rect 44192 16574 44220 76570
rect 45560 19984 45612 19990
rect 45560 19926 45612 19932
rect 45572 16574 45600 19926
rect 44192 16546 45048 16574
rect 45572 16546 46152 16574
rect 44272 7676 44324 7682
rect 44272 7618 44324 7624
rect 44284 480 44312 7618
rect 43046 354 43158 480
rect 42812 326 43158 354
rect 43046 -960 43158 326
rect 44242 -960 44354 480
rect 45020 354 45048 16546
rect 46124 3482 46152 16546
rect 46216 5098 46244 78066
rect 57244 78056 57296 78062
rect 57244 77998 57296 78004
rect 53838 75440 53894 75449
rect 51080 75404 51132 75410
rect 53838 75375 53894 75384
rect 51080 75346 51132 75352
rect 50160 9036 50212 9042
rect 50160 8978 50212 8984
rect 48964 7744 49016 7750
rect 48964 7686 49016 7692
rect 46204 5092 46256 5098
rect 46204 5034 46256 5040
rect 47860 3596 47912 3602
rect 47860 3538 47912 3544
rect 46124 3454 46704 3482
rect 46676 480 46704 3454
rect 47872 480 47900 3538
rect 48976 480 49004 7686
rect 50172 480 50200 8978
rect 45438 354 45550 480
rect 45020 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51092 354 51120 75346
rect 53852 16574 53880 75375
rect 53852 16546 54984 16574
rect 53748 9104 53800 9110
rect 53748 9046 53800 9052
rect 52552 5092 52604 5098
rect 52552 5034 52604 5040
rect 52564 480 52592 5034
rect 53760 480 53788 9046
rect 54956 480 54984 16546
rect 57150 8936 57206 8945
rect 57150 8871 57206 8880
rect 56046 7848 56102 7857
rect 56046 7783 56102 7792
rect 56060 480 56088 7783
rect 57164 3482 57192 8871
rect 57256 6322 57284 77998
rect 86960 76764 87012 76770
rect 86960 76706 87012 76712
rect 69020 76696 69072 76702
rect 69020 76638 69072 76644
rect 57978 75576 58034 75585
rect 57978 75511 58034 75520
rect 57992 16574 58020 75511
rect 64880 73976 64932 73982
rect 64880 73918 64932 73924
rect 64892 16574 64920 73918
rect 69032 16574 69060 76638
rect 78680 71052 78732 71058
rect 78680 70994 78732 71000
rect 70400 44940 70452 44946
rect 70400 44882 70452 44888
rect 70412 16574 70440 44882
rect 74540 22840 74592 22846
rect 74540 22782 74592 22788
rect 74552 16574 74580 22782
rect 78692 16574 78720 70994
rect 85580 20052 85632 20058
rect 85580 19994 85632 20000
rect 85592 16574 85620 19994
rect 86972 16574 87000 76706
rect 88340 36576 88392 36582
rect 88340 36518 88392 36524
rect 88352 16574 88380 36518
rect 89732 16574 89760 78134
rect 111798 76936 111854 76945
rect 111798 76871 111854 76880
rect 102140 76832 102192 76838
rect 93858 76800 93914 76809
rect 102140 76774 102192 76780
rect 93858 76735 93914 76744
rect 91098 44840 91154 44849
rect 91098 44775 91154 44784
rect 91112 16574 91140 44775
rect 57992 16546 58480 16574
rect 64892 16546 65104 16574
rect 69032 16546 69888 16574
rect 70412 16546 71544 16574
rect 74552 16546 75040 16574
rect 78692 16546 79272 16574
rect 85592 16546 85712 16574
rect 86972 16546 87552 16574
rect 88352 16546 89208 16574
rect 89732 16546 89944 16574
rect 91112 16546 91600 16574
rect 57244 6316 57296 6322
rect 57244 6258 57296 6264
rect 57164 3454 57284 3482
rect 57256 480 57284 3454
rect 58452 480 58480 16546
rect 64328 9308 64380 9314
rect 64328 9250 64380 9256
rect 63224 9240 63276 9246
rect 63224 9182 63276 9188
rect 60832 9172 60884 9178
rect 60832 9114 60884 9120
rect 59636 5160 59688 5166
rect 59636 5102 59688 5108
rect 59648 480 59676 5102
rect 60844 480 60872 9114
rect 62028 3664 62080 3670
rect 62028 3606 62080 3612
rect 62040 480 62068 3606
rect 63236 480 63264 9182
rect 64340 480 64368 9250
rect 51326 354 51438 480
rect 51092 326 51438 354
rect 51326 -960 51438 326
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 354 65104 16546
rect 67916 9376 67968 9382
rect 67916 9318 67968 9324
rect 66720 6316 66772 6322
rect 66720 6258 66772 6264
rect 66732 480 66760 6258
rect 67928 480 67956 9318
rect 69112 3732 69164 3738
rect 69112 3674 69164 3680
rect 69124 480 69152 3674
rect 65494 354 65606 480
rect 65076 326 65606 354
rect 65494 -960 65606 326
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 69860 354 69888 16546
rect 71516 480 71544 16546
rect 73802 6216 73858 6225
rect 73802 6151 73858 6160
rect 72606 3496 72662 3505
rect 72606 3431 72662 3440
rect 72620 480 72648 3431
rect 73816 480 73844 6151
rect 75012 480 75040 16546
rect 78586 9072 78642 9081
rect 78586 9007 78642 9016
rect 77392 6384 77444 6390
rect 77392 6326 77444 6332
rect 76196 3800 76248 3806
rect 76196 3742 76248 3748
rect 76208 480 76236 3742
rect 77404 480 77432 6326
rect 78600 480 78628 9007
rect 70278 354 70390 480
rect 69860 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79244 354 79272 16546
rect 81624 10532 81676 10538
rect 81624 10474 81676 10480
rect 80888 6452 80940 6458
rect 80888 6394 80940 6400
rect 80900 480 80928 6394
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 81636 354 81664 10474
rect 84476 6520 84528 6526
rect 84476 6462 84528 6468
rect 83280 3868 83332 3874
rect 83280 3810 83332 3816
rect 83292 480 83320 3810
rect 84488 480 84516 6462
rect 85684 480 85712 16546
rect 86868 5228 86920 5234
rect 86868 5170 86920 5176
rect 86880 480 86908 5170
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87524 354 87552 16546
rect 89180 480 89208 16546
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91572 480 91600 16546
rect 92478 10296 92534 10305
rect 92478 10231 92534 10240
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 10231
rect 93872 3466 93900 76735
rect 93952 74044 94004 74050
rect 93952 73986 94004 73992
rect 93860 3460 93912 3466
rect 93860 3402 93912 3408
rect 93964 480 93992 73986
rect 95240 53100 95292 53106
rect 95240 53042 95292 53048
rect 95252 16574 95280 53042
rect 95252 16546 95832 16574
rect 94780 3460 94832 3466
rect 94780 3402 94832 3408
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 94792 354 94820 3402
rect 95118 354 95230 480
rect 94792 326 95230 354
rect 95804 354 95832 16546
rect 99840 10600 99892 10606
rect 99840 10542 99892 10548
rect 98644 7812 98696 7818
rect 98644 7754 98696 7760
rect 97448 5296 97500 5302
rect 97448 5238 97500 5244
rect 97460 480 97488 5238
rect 98656 480 98684 7754
rect 99852 480 99880 10542
rect 102152 6914 102180 76774
rect 107660 75336 107712 75342
rect 107660 75278 107712 75284
rect 102232 65544 102284 65550
rect 102232 65486 102284 65492
rect 102244 16574 102272 65486
rect 107672 16574 107700 75278
rect 111812 16574 111840 76871
rect 118436 22778 118464 81495
rect 118528 60722 118556 82991
rect 119448 80782 119476 106898
rect 120644 104553 120672 113146
rect 120630 104544 120686 104553
rect 120630 104479 120686 104488
rect 120908 99408 120960 99414
rect 120908 99350 120960 99356
rect 120724 86284 120776 86290
rect 120724 86226 120776 86232
rect 120630 84280 120686 84289
rect 120448 84244 120500 84250
rect 120630 84215 120686 84224
rect 120448 84186 120500 84192
rect 119988 82408 120040 82414
rect 119988 82350 120040 82356
rect 119436 80776 119488 80782
rect 119436 80718 119488 80724
rect 120000 80102 120028 82350
rect 119988 80096 120040 80102
rect 119988 80038 120040 80044
rect 120460 79218 120488 84186
rect 120644 81433 120672 84215
rect 120630 81424 120686 81433
rect 120630 81359 120686 81368
rect 120448 79212 120500 79218
rect 120448 79154 120500 79160
rect 120632 77648 120684 77654
rect 120632 77590 120684 77596
rect 118700 74112 118752 74118
rect 118700 74054 118752 74060
rect 118516 60716 118568 60722
rect 118516 60658 118568 60664
rect 118424 22772 118476 22778
rect 118424 22714 118476 22720
rect 117320 18760 117372 18766
rect 117320 18702 117372 18708
rect 102244 16546 103376 16574
rect 107672 16546 108160 16574
rect 111812 16546 112392 16574
rect 102152 6886 102272 6914
rect 101036 5364 101088 5370
rect 101036 5306 101088 5312
rect 101048 480 101076 5306
rect 102244 480 102272 6886
rect 103348 480 103376 16546
rect 106464 10668 106516 10674
rect 106464 10610 106516 10616
rect 105728 7880 105780 7886
rect 105728 7822 105780 7828
rect 104532 6588 104584 6594
rect 104532 6530 104584 6536
rect 104544 480 104572 6530
rect 105740 480 105768 7822
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 95118 -960 95230 326
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106476 354 106504 10610
rect 108132 480 108160 16546
rect 110510 10432 110566 10441
rect 110510 10367 110566 10376
rect 109314 7984 109370 7993
rect 109314 7919 109370 7928
rect 109328 480 109356 7919
rect 110524 480 110552 10367
rect 111614 6352 111670 6361
rect 111614 6287 111670 6296
rect 111628 480 111656 6287
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 16546
rect 114008 14544 114060 14550
rect 114008 14486 114060 14492
rect 114020 480 114048 14486
rect 116400 7948 116452 7954
rect 116400 7890 116452 7896
rect 115204 6656 115256 6662
rect 115204 6598 115256 6604
rect 115216 480 115244 6598
rect 116412 480 116440 7890
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117332 354 117360 18702
rect 118712 16574 118740 74054
rect 120644 70394 120672 77590
rect 120736 77314 120764 86226
rect 120816 77716 120868 77722
rect 120816 77658 120868 77664
rect 120724 77308 120776 77314
rect 120724 77250 120776 77256
rect 120644 70366 120764 70394
rect 120080 40316 120132 40322
rect 120080 40258 120132 40264
rect 120092 16574 120120 40258
rect 118712 16546 118832 16574
rect 120092 16546 120672 16574
rect 118804 480 118832 16546
rect 119896 4140 119948 4146
rect 119896 4082 119948 4088
rect 119908 480 119936 4082
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 16546
rect 120736 14482 120764 70366
rect 120828 19990 120856 77658
rect 120920 76362 120948 99350
rect 178498 81016 178554 81025
rect 178498 80951 178554 80960
rect 174820 80708 174872 80714
rect 174820 80650 174872 80656
rect 174912 80708 174964 80714
rect 174912 80650 174964 80656
rect 174728 80504 174780 80510
rect 174340 80430 174584 80458
rect 174728 80446 174780 80452
rect 174452 80300 174504 80306
rect 174452 80242 174504 80248
rect 124128 80028 124180 80034
rect 124128 79970 124180 79976
rect 124784 80022 125580 80050
rect 124140 78554 124168 79970
rect 124140 78526 124260 78554
rect 123576 77784 123628 77790
rect 123576 77726 123628 77732
rect 122288 77580 122340 77586
rect 122288 77522 122340 77528
rect 122104 77512 122156 77518
rect 122104 77454 122156 77460
rect 120908 76356 120960 76362
rect 120908 76298 120960 76304
rect 121460 75472 121512 75478
rect 121460 75414 121512 75420
rect 120816 19984 120868 19990
rect 120816 19926 120868 19932
rect 121472 16574 121500 75414
rect 121472 16546 122052 16574
rect 120724 14476 120776 14482
rect 120724 14418 120776 14424
rect 122024 3482 122052 16546
rect 122116 4962 122144 77454
rect 122196 75608 122248 75614
rect 122196 75550 122248 75556
rect 122104 4956 122156 4962
rect 122104 4898 122156 4904
rect 122208 3670 122236 75550
rect 122300 18698 122328 77522
rect 122840 76900 122892 76906
rect 122840 76842 122892 76848
rect 122288 18692 122340 18698
rect 122288 18634 122340 18640
rect 122852 16574 122880 76842
rect 123484 76764 123536 76770
rect 123484 76706 123536 76712
rect 123496 76430 123524 76706
rect 123484 76424 123536 76430
rect 123484 76366 123536 76372
rect 123588 70394 123616 77726
rect 124232 76498 124260 78526
rect 124220 76492 124272 76498
rect 124220 76434 124272 76440
rect 124784 70394 124812 80022
rect 125658 79880 125686 80036
rect 125750 79937 125778 80036
rect 125842 79966 125870 80036
rect 125934 79966 125962 80036
rect 126026 79966 126054 80036
rect 125830 79960 125882 79966
rect 125612 79852 125686 79880
rect 125736 79928 125792 79937
rect 125830 79902 125882 79908
rect 125922 79960 125974 79966
rect 125922 79902 125974 79908
rect 126014 79960 126066 79966
rect 126014 79902 126066 79908
rect 125736 79863 125792 79872
rect 125048 78260 125100 78266
rect 125048 78202 125100 78208
rect 124956 77376 125008 77382
rect 124956 77318 125008 77324
rect 124864 77036 124916 77042
rect 124864 76978 124916 76984
rect 123496 70366 123616 70394
rect 124232 70366 124812 70394
rect 123496 40322 123524 70366
rect 123484 40316 123536 40322
rect 123484 40258 123536 40264
rect 122852 16546 123064 16574
rect 122196 3664 122248 3670
rect 122196 3606 122248 3612
rect 122024 3454 122328 3482
rect 122300 480 122328 3454
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123036 354 123064 16546
rect 124232 8974 124260 70366
rect 124312 21412 124364 21418
rect 124312 21354 124364 21360
rect 124324 16574 124352 21354
rect 124324 16546 124720 16574
rect 124220 8968 124272 8974
rect 124220 8910 124272 8916
rect 124692 480 124720 16546
rect 124876 4146 124904 76978
rect 124968 15910 124996 77318
rect 125060 36582 125088 78202
rect 125324 77920 125376 77926
rect 125324 77862 125376 77868
rect 125232 77852 125284 77858
rect 125232 77794 125284 77800
rect 125140 77308 125192 77314
rect 125140 77250 125192 77256
rect 125152 42090 125180 77250
rect 125244 53106 125272 77794
rect 125336 65550 125364 77862
rect 125612 76537 125640 79852
rect 125876 79824 125928 79830
rect 126118 79812 126146 80036
rect 126210 79937 126238 80036
rect 126196 79928 126252 79937
rect 126196 79863 126252 79872
rect 126302 79812 126330 80036
rect 126394 79966 126422 80036
rect 126382 79960 126434 79966
rect 126382 79902 126434 79908
rect 126486 79898 126514 80036
rect 126578 79966 126606 80036
rect 126670 79971 126698 80036
rect 126566 79960 126618 79966
rect 126566 79902 126618 79908
rect 126656 79962 126712 79971
rect 126474 79892 126526 79898
rect 126656 79897 126712 79906
rect 126474 79834 126526 79840
rect 126118 79784 126192 79812
rect 126302 79784 126376 79812
rect 125876 79766 125928 79772
rect 126164 79778 126192 79784
rect 125692 79756 125744 79762
rect 125692 79698 125744 79704
rect 125704 77994 125732 79698
rect 125782 78840 125838 78849
rect 125782 78775 125838 78784
rect 125692 77988 125744 77994
rect 125692 77930 125744 77936
rect 125598 76528 125654 76537
rect 125598 76463 125654 76472
rect 125692 75880 125744 75886
rect 125692 75822 125744 75828
rect 125704 75206 125732 75822
rect 125692 75200 125744 75206
rect 125692 75142 125744 75148
rect 125692 74996 125744 75002
rect 125692 74938 125744 74944
rect 125324 65544 125376 65550
rect 125324 65486 125376 65492
rect 125232 53100 125284 53106
rect 125232 53042 125284 53048
rect 125140 42084 125192 42090
rect 125140 42026 125192 42032
rect 125048 36576 125100 36582
rect 125048 36518 125100 36524
rect 124956 15904 125008 15910
rect 124956 15846 125008 15852
rect 124864 4140 124916 4146
rect 124864 4082 124916 4088
rect 125704 3534 125732 74938
rect 125796 4826 125824 78775
rect 125888 78713 125916 79766
rect 126164 79750 126238 79778
rect 126210 79744 126238 79750
rect 126210 79716 126284 79744
rect 125968 79620 126020 79626
rect 125968 79562 126020 79568
rect 126152 79620 126204 79626
rect 126152 79562 126204 79568
rect 125874 78704 125930 78713
rect 125874 78639 125930 78648
rect 125874 77616 125930 77625
rect 125874 77551 125930 77560
rect 125888 77518 125916 77551
rect 125876 77512 125928 77518
rect 125876 77454 125928 77460
rect 125980 75206 126008 79562
rect 126060 78668 126112 78674
rect 126060 78610 126112 78616
rect 125968 75200 126020 75206
rect 125968 75142 126020 75148
rect 125876 75132 125928 75138
rect 125876 75074 125928 75080
rect 125888 4894 125916 75074
rect 125968 75064 126020 75070
rect 125968 75006 126020 75012
rect 125980 6186 126008 75006
rect 126072 7614 126100 78610
rect 126164 10334 126192 79562
rect 126256 75886 126284 79716
rect 126348 78674 126376 79784
rect 126612 79756 126664 79762
rect 126762 79744 126790 80036
rect 126612 79698 126664 79704
rect 126716 79716 126790 79744
rect 126518 79656 126574 79665
rect 126518 79591 126574 79600
rect 126428 79552 126480 79558
rect 126428 79494 126480 79500
rect 126336 78668 126388 78674
rect 126336 78610 126388 78616
rect 126336 78532 126388 78538
rect 126336 78474 126388 78480
rect 126244 75880 126296 75886
rect 126244 75822 126296 75828
rect 126244 75200 126296 75206
rect 126244 75142 126296 75148
rect 126256 18630 126284 75142
rect 126244 18624 126296 18630
rect 126244 18566 126296 18572
rect 126152 10328 126204 10334
rect 126152 10270 126204 10276
rect 126348 9314 126376 78474
rect 126336 9308 126388 9314
rect 126336 9250 126388 9256
rect 126060 7608 126112 7614
rect 126060 7550 126112 7556
rect 125968 6180 126020 6186
rect 125968 6122 126020 6128
rect 125876 4888 125928 4894
rect 125876 4830 125928 4836
rect 125784 4820 125836 4826
rect 125784 4762 125836 4768
rect 125876 4140 125928 4146
rect 125876 4082 125928 4088
rect 125692 3528 125744 3534
rect 125692 3470 125744 3476
rect 125888 480 125916 4082
rect 126440 4010 126468 79494
rect 126532 77382 126560 79591
rect 126520 77376 126572 77382
rect 126520 77318 126572 77324
rect 126624 75138 126652 79698
rect 126716 78130 126744 79716
rect 126854 79676 126882 80036
rect 126946 79898 126974 80036
rect 126934 79892 126986 79898
rect 126934 79834 126986 79840
rect 127038 79744 127066 80036
rect 127130 79898 127158 80036
rect 127222 79903 127250 80036
rect 127118 79892 127170 79898
rect 127118 79834 127170 79840
rect 127208 79894 127264 79903
rect 127314 79898 127342 80036
rect 127208 79829 127264 79838
rect 127302 79892 127354 79898
rect 127302 79834 127354 79840
rect 126808 79648 126882 79676
rect 126992 79716 127066 79744
rect 127164 79756 127216 79762
rect 126704 78124 126756 78130
rect 126704 78066 126756 78072
rect 126612 75132 126664 75138
rect 126612 75074 126664 75080
rect 126808 75002 126836 79648
rect 126888 79552 126940 79558
rect 126888 79494 126940 79500
rect 126900 75070 126928 79494
rect 126992 77314 127020 79716
rect 127164 79698 127216 79704
rect 127256 79756 127308 79762
rect 127256 79698 127308 79704
rect 127070 79656 127126 79665
rect 127070 79591 127126 79600
rect 126980 77308 127032 77314
rect 126980 77250 127032 77256
rect 127084 76673 127112 79591
rect 127176 77489 127204 79698
rect 127162 77480 127218 77489
rect 127162 77415 127218 77424
rect 127268 77353 127296 79698
rect 127406 79676 127434 80036
rect 127360 79665 127434 79676
rect 127346 79656 127434 79665
rect 127402 79648 127434 79656
rect 127498 79676 127526 80036
rect 127590 79744 127618 80036
rect 127682 79971 127710 80036
rect 127668 79962 127724 79971
rect 127774 79966 127802 80036
rect 127668 79897 127724 79906
rect 127762 79960 127814 79966
rect 127762 79902 127814 79908
rect 127866 79898 127894 80036
rect 127958 79898 127986 80036
rect 128050 79966 128078 80036
rect 128038 79960 128090 79966
rect 128142 79937 128170 80036
rect 128234 79966 128262 80036
rect 128222 79960 128274 79966
rect 128038 79902 128090 79908
rect 128128 79928 128184 79937
rect 127854 79892 127906 79898
rect 127854 79834 127906 79840
rect 127946 79892 127998 79898
rect 128222 79902 128274 79908
rect 128128 79863 128184 79872
rect 127946 79834 127998 79840
rect 128084 79824 128136 79830
rect 127806 79792 127862 79801
rect 127590 79716 127664 79744
rect 128326 79801 128354 80036
rect 128418 79898 128446 80036
rect 128406 79892 128458 79898
rect 128406 79834 128458 79840
rect 128084 79766 128136 79772
rect 128312 79792 128368 79801
rect 127806 79727 127862 79736
rect 127900 79756 127952 79762
rect 127498 79648 127572 79676
rect 127346 79591 127402 79600
rect 127348 79552 127400 79558
rect 127348 79494 127400 79500
rect 127254 77344 127310 77353
rect 127254 77279 127310 77288
rect 127360 77194 127388 79494
rect 127440 79416 127492 79422
rect 127440 79358 127492 79364
rect 127176 77166 127388 77194
rect 127070 76664 127126 76673
rect 127070 76599 127126 76608
rect 126980 75744 127032 75750
rect 126980 75686 127032 75692
rect 126992 75478 127020 75686
rect 126980 75472 127032 75478
rect 126980 75414 127032 75420
rect 126888 75064 126940 75070
rect 126888 75006 126940 75012
rect 126796 74996 126848 75002
rect 126796 74938 126848 74944
rect 127070 44976 127126 44985
rect 127070 44911 127126 44920
rect 127084 6914 127112 44911
rect 127176 10402 127204 77166
rect 127256 75200 127308 75206
rect 127256 75142 127308 75148
rect 127268 10470 127296 75142
rect 127348 75132 127400 75138
rect 127348 75074 127400 75080
rect 127360 44878 127388 75074
rect 127348 44872 127400 44878
rect 127348 44814 127400 44820
rect 127256 10464 127308 10470
rect 127256 10406 127308 10412
rect 127164 10396 127216 10402
rect 127164 10338 127216 10344
rect 127084 6886 127388 6914
rect 126428 4004 126480 4010
rect 126428 3946 126480 3952
rect 126980 3596 127032 3602
rect 126980 3538 127032 3544
rect 126992 480 127020 3538
rect 127360 3482 127388 6886
rect 127452 5030 127480 79358
rect 127544 79234 127572 79648
rect 127636 79354 127664 79716
rect 127714 79656 127770 79665
rect 127714 79591 127770 79600
rect 127624 79348 127676 79354
rect 127624 79290 127676 79296
rect 127544 79206 127664 79234
rect 127532 79076 127584 79082
rect 127532 79018 127584 79024
rect 127544 6254 127572 79018
rect 127636 78062 127664 79206
rect 127728 79082 127756 79591
rect 127716 79076 127768 79082
rect 127716 79018 127768 79024
rect 127716 78736 127768 78742
rect 127716 78678 127768 78684
rect 127624 78056 127676 78062
rect 127624 77998 127676 78004
rect 127624 77444 127676 77450
rect 127624 77386 127676 77392
rect 127532 6248 127584 6254
rect 127532 6190 127584 6196
rect 127440 5024 127492 5030
rect 127440 4966 127492 4972
rect 127636 3670 127664 77386
rect 127728 9042 127756 78678
rect 127820 73914 127848 79727
rect 127900 79698 127952 79704
rect 127992 79756 128044 79762
rect 127992 79698 128044 79704
rect 127912 79490 127940 79698
rect 127900 79484 127952 79490
rect 127900 79426 127952 79432
rect 127900 79348 127952 79354
rect 127900 79290 127952 79296
rect 127808 73908 127860 73914
rect 127808 73850 127860 73856
rect 127912 73846 127940 79290
rect 128004 76566 128032 79698
rect 128096 77586 128124 79766
rect 128312 79727 128368 79736
rect 128510 79744 128538 80036
rect 128602 79898 128630 80036
rect 128590 79892 128642 79898
rect 128590 79834 128642 79840
rect 128694 79830 128722 80036
rect 128786 79937 128814 80036
rect 128878 79966 128906 80036
rect 128970 79966 128998 80036
rect 128866 79960 128918 79966
rect 128772 79928 128828 79937
rect 128866 79902 128918 79908
rect 128958 79960 129010 79966
rect 129062 79937 129090 80036
rect 128958 79902 129010 79908
rect 129048 79928 129104 79937
rect 128772 79863 128828 79872
rect 129048 79863 129104 79872
rect 128682 79824 128734 79830
rect 129154 79812 129182 80036
rect 128682 79766 128734 79772
rect 129002 79792 129058 79801
rect 128820 79756 128872 79762
rect 128510 79716 128584 79744
rect 128268 79688 128320 79694
rect 128174 79656 128230 79665
rect 128268 79630 128320 79636
rect 128174 79591 128230 79600
rect 128084 77580 128136 77586
rect 128084 77522 128136 77528
rect 127992 76560 128044 76566
rect 127992 76502 128044 76508
rect 128188 75206 128216 79591
rect 128176 75200 128228 75206
rect 128176 75142 128228 75148
rect 128280 75138 128308 79630
rect 128360 79620 128412 79626
rect 128360 79562 128412 79568
rect 128452 79620 128504 79626
rect 128452 79562 128504 79568
rect 128372 75313 128400 79562
rect 128464 77654 128492 79562
rect 128556 78849 128584 79716
rect 129002 79727 129058 79736
rect 129108 79784 129182 79812
rect 128820 79698 128872 79704
rect 128728 79688 128780 79694
rect 128726 79656 128728 79665
rect 128780 79656 128782 79665
rect 128636 79620 128688 79626
rect 128726 79591 128782 79600
rect 128636 79562 128688 79568
rect 128542 78840 128598 78849
rect 128542 78775 128598 78784
rect 128452 77648 128504 77654
rect 128452 77590 128504 77596
rect 128358 75304 128414 75313
rect 128358 75239 128414 75248
rect 128544 75268 128596 75274
rect 128544 75210 128596 75216
rect 128268 75132 128320 75138
rect 128268 75074 128320 75080
rect 128360 75064 128412 75070
rect 128360 75006 128412 75012
rect 127900 73840 127952 73846
rect 127900 73782 127952 73788
rect 127716 9036 127768 9042
rect 127716 8978 127768 8984
rect 127624 3664 127676 3670
rect 127624 3606 127676 3612
rect 127360 3454 128216 3482
rect 128188 480 128216 3454
rect 128372 490 128400 75006
rect 128452 74996 128504 75002
rect 128452 74938 128504 74944
rect 128464 5098 128492 74938
rect 128556 7750 128584 75210
rect 128544 7744 128596 7750
rect 128544 7686 128596 7692
rect 128648 7682 128676 79562
rect 128832 79370 128860 79698
rect 128832 79342 128952 79370
rect 128728 78668 128780 78674
rect 128728 78610 128780 78616
rect 128740 75410 128768 78610
rect 128818 78568 128874 78577
rect 128818 78503 128874 78512
rect 128832 76634 128860 78503
rect 128820 76628 128872 76634
rect 128820 76570 128872 76576
rect 128728 75404 128780 75410
rect 128728 75346 128780 75352
rect 128924 75206 128952 79342
rect 129016 78742 129044 79727
rect 129004 78736 129056 78742
rect 129004 78678 129056 78684
rect 129108 77840 129136 79784
rect 129246 79744 129274 80036
rect 129016 77812 129136 77840
rect 129200 79716 129274 79744
rect 129016 77722 129044 77812
rect 129004 77716 129056 77722
rect 129004 77658 129056 77664
rect 129096 77716 129148 77722
rect 129096 77658 129148 77664
rect 129004 77580 129056 77586
rect 129004 77522 129056 77528
rect 128912 75200 128964 75206
rect 128912 75142 128964 75148
rect 128728 75132 128780 75138
rect 128728 75074 128780 75080
rect 128740 9110 128768 75074
rect 128728 9104 128780 9110
rect 128728 9046 128780 9052
rect 128636 7676 128688 7682
rect 128636 7618 128688 7624
rect 128452 5092 128504 5098
rect 128452 5034 128504 5040
rect 129016 3806 129044 77522
rect 129108 9178 129136 77658
rect 129200 77450 129228 79716
rect 129338 79676 129366 80036
rect 129430 79937 129458 80036
rect 129416 79928 129472 79937
rect 129416 79863 129472 79872
rect 129522 79812 129550 80036
rect 129614 79898 129642 80036
rect 129602 79892 129654 79898
rect 129602 79834 129654 79840
rect 129476 79784 129550 79812
rect 129476 79778 129504 79784
rect 129292 79648 129366 79676
rect 129430 79750 129504 79778
rect 129188 77444 129240 77450
rect 129188 77386 129240 77392
rect 129292 75274 129320 79648
rect 129430 79608 129458 79750
rect 129706 79744 129734 80036
rect 129798 79903 129826 80036
rect 129784 79894 129840 79903
rect 129784 79829 129840 79838
rect 129890 79830 129918 80036
rect 129982 79971 130010 80036
rect 129968 79962 130024 79971
rect 130074 79966 130102 80036
rect 129968 79897 130024 79906
rect 130062 79960 130114 79966
rect 130062 79902 130114 79908
rect 130166 79830 130194 80036
rect 130258 79898 130286 80036
rect 130350 79966 130378 80036
rect 130338 79960 130390 79966
rect 130338 79902 130390 79908
rect 130442 79898 130470 80036
rect 130534 79937 130562 80036
rect 130626 79966 130654 80036
rect 130718 79966 130746 80036
rect 130810 79966 130838 80036
rect 130614 79960 130666 79966
rect 130520 79928 130576 79937
rect 130246 79892 130298 79898
rect 130246 79834 130298 79840
rect 130430 79892 130482 79898
rect 130614 79902 130666 79908
rect 130706 79960 130758 79966
rect 130706 79902 130758 79908
rect 130798 79960 130850 79966
rect 130798 79902 130850 79908
rect 130520 79863 130576 79872
rect 130430 79834 130482 79840
rect 129878 79824 129930 79830
rect 129878 79766 129930 79772
rect 130154 79824 130206 79830
rect 130154 79766 130206 79772
rect 130566 79792 130622 79801
rect 129660 79716 129734 79744
rect 130016 79756 130068 79762
rect 129384 79580 129458 79608
rect 129556 79620 129608 79626
rect 129384 78674 129412 79580
rect 129556 79562 129608 79568
rect 129464 79484 129516 79490
rect 129464 79426 129516 79432
rect 129372 78668 129424 78674
rect 129372 78610 129424 78616
rect 129370 78568 129426 78577
rect 129370 78503 129426 78512
rect 129280 75268 129332 75274
rect 129280 75210 129332 75216
rect 129384 64874 129412 78503
rect 129476 77858 129504 79426
rect 129464 77852 129516 77858
rect 129464 77794 129516 77800
rect 129568 75002 129596 79562
rect 129660 75138 129688 79716
rect 130016 79698 130068 79704
rect 130292 79756 130344 79762
rect 130292 79698 130344 79704
rect 130384 79756 130436 79762
rect 130902 79744 130930 80036
rect 130994 79966 131022 80036
rect 130982 79960 131034 79966
rect 130982 79902 131034 79908
rect 131086 79812 131114 80036
rect 131178 79898 131206 80036
rect 131270 79898 131298 80036
rect 131362 79966 131390 80036
rect 131350 79960 131402 79966
rect 131350 79902 131402 79908
rect 131166 79892 131218 79898
rect 131166 79834 131218 79840
rect 131258 79892 131310 79898
rect 131258 79834 131310 79840
rect 131040 79784 131114 79812
rect 131348 79826 131404 79835
rect 131040 79778 131068 79784
rect 130566 79727 130622 79736
rect 130384 79698 130436 79704
rect 129832 79688 129884 79694
rect 129832 79630 129884 79636
rect 129740 79620 129792 79626
rect 129740 79562 129792 79568
rect 129648 75132 129700 75138
rect 129648 75074 129700 75080
rect 129556 74996 129608 75002
rect 129556 74938 129608 74944
rect 129752 73982 129780 79562
rect 129844 78713 129872 79630
rect 130028 78849 130056 79698
rect 130108 79688 130160 79694
rect 130108 79630 130160 79636
rect 130014 78840 130070 78849
rect 130014 78775 130070 78784
rect 129830 78704 129886 78713
rect 129830 78639 129886 78648
rect 130120 78418 130148 79630
rect 129936 78390 130148 78418
rect 129832 77376 129884 77382
rect 129832 77318 129884 77324
rect 129740 73976 129792 73982
rect 129740 73918 129792 73924
rect 129844 70394 129872 77318
rect 129200 64846 129412 64874
rect 129752 70366 129872 70394
rect 129200 22846 129228 64846
rect 129188 22840 129240 22846
rect 129188 22782 129240 22788
rect 129752 16574 129780 70366
rect 129752 16546 129872 16574
rect 129096 9172 129148 9178
rect 129096 9114 129148 9120
rect 129004 3800 129056 3806
rect 129004 3742 129056 3748
rect 129844 3482 129872 16546
rect 129936 5166 129964 78390
rect 130304 77722 130332 79698
rect 130292 77716 130344 77722
rect 130292 77658 130344 77664
rect 130396 77294 130424 79698
rect 130476 79688 130528 79694
rect 130476 79630 130528 79636
rect 130120 77266 130424 77294
rect 130016 75676 130068 75682
rect 130016 75618 130068 75624
rect 130028 6322 130056 75618
rect 130120 9246 130148 77266
rect 130488 75614 130516 79630
rect 130580 78538 130608 79727
rect 130856 79716 130930 79744
rect 130994 79750 131068 79778
rect 131348 79761 131404 79770
rect 130660 79688 130712 79694
rect 130660 79630 130712 79636
rect 130568 78532 130620 78538
rect 130568 78474 130620 78480
rect 130672 75682 130700 79630
rect 130752 79620 130804 79626
rect 130752 79562 130804 79568
rect 130660 75676 130712 75682
rect 130660 75618 130712 75624
rect 130476 75608 130528 75614
rect 130476 75550 130528 75556
rect 130764 75426 130792 79562
rect 130212 75398 130792 75426
rect 130212 9382 130240 75398
rect 130292 75268 130344 75274
rect 130292 75210 130344 75216
rect 130304 44946 130332 75210
rect 130382 74488 130438 74497
rect 130382 74423 130438 74432
rect 130292 44940 130344 44946
rect 130292 44882 130344 44888
rect 130200 9376 130252 9382
rect 130200 9318 130252 9324
rect 130108 9240 130160 9246
rect 130108 9182 130160 9188
rect 130016 6316 130068 6322
rect 130016 6258 130068 6264
rect 129924 5160 129976 5166
rect 129924 5102 129976 5108
rect 130396 3602 130424 74423
rect 130856 70394 130884 79716
rect 130994 79676 131022 79750
rect 131454 79676 131482 80036
rect 131546 79966 131574 80036
rect 131638 79971 131666 80036
rect 131534 79960 131586 79966
rect 131534 79902 131586 79908
rect 131624 79962 131680 79971
rect 131624 79897 131680 79906
rect 131578 79792 131634 79801
rect 131578 79727 131634 79736
rect 130994 79648 131068 79676
rect 130936 79552 130988 79558
rect 130936 79494 130988 79500
rect 130948 76702 130976 79494
rect 130936 76696 130988 76702
rect 130936 76638 130988 76644
rect 131040 75274 131068 79648
rect 131408 79648 131482 79676
rect 131304 79620 131356 79626
rect 131304 79562 131356 79568
rect 131212 79552 131264 79558
rect 131212 79494 131264 79500
rect 131120 79416 131172 79422
rect 131120 79358 131172 79364
rect 131132 79286 131160 79358
rect 131120 79280 131172 79286
rect 131120 79222 131172 79228
rect 131028 75268 131080 75274
rect 131028 75210 131080 75216
rect 131224 73273 131252 79494
rect 131316 77081 131344 79562
rect 131408 77586 131436 79648
rect 131488 79552 131540 79558
rect 131488 79494 131540 79500
rect 131396 77580 131448 77586
rect 131396 77522 131448 77528
rect 131302 77072 131358 77081
rect 131302 77007 131358 77016
rect 131396 76832 131448 76838
rect 131396 76774 131448 76780
rect 131304 75200 131356 75206
rect 131304 75142 131356 75148
rect 131210 73264 131266 73273
rect 131210 73199 131266 73208
rect 130764 70366 130884 70394
rect 130764 64874 130792 70366
rect 130672 64846 130792 64874
rect 130672 3738 130700 64846
rect 131316 6526 131344 75142
rect 131304 6520 131356 6526
rect 131304 6462 131356 6468
rect 131408 6458 131436 76774
rect 131396 6452 131448 6458
rect 131396 6394 131448 6400
rect 131500 6390 131528 79494
rect 131592 10538 131620 79727
rect 131730 79676 131758 80036
rect 131822 79830 131850 80036
rect 131914 79971 131942 80036
rect 131900 79962 131956 79971
rect 131900 79897 131956 79906
rect 132006 79898 132034 80036
rect 131994 79892 132046 79898
rect 131994 79834 132046 79840
rect 131810 79824 131862 79830
rect 131810 79766 131862 79772
rect 131948 79756 132000 79762
rect 132098 79744 132126 80036
rect 132190 79830 132218 80036
rect 132178 79824 132230 79830
rect 132282 79812 132310 80036
rect 132374 79937 132402 80036
rect 132360 79928 132416 79937
rect 132360 79863 132416 79872
rect 132466 79830 132494 80036
rect 132558 79971 132586 80036
rect 132544 79962 132600 79971
rect 132650 79966 132678 80036
rect 132544 79897 132600 79906
rect 132638 79960 132690 79966
rect 132742 79937 132770 80036
rect 132638 79902 132690 79908
rect 132728 79928 132784 79937
rect 132728 79863 132784 79872
rect 132454 79824 132506 79830
rect 132282 79784 132356 79812
rect 132178 79766 132230 79772
rect 132328 79778 132356 79784
rect 132328 79750 132402 79778
rect 132834 79812 132862 80036
rect 132926 79971 132954 80036
rect 132912 79962 132968 79971
rect 133018 79966 133046 80036
rect 132912 79897 132968 79906
rect 133006 79960 133058 79966
rect 133006 79902 133058 79908
rect 132834 79784 132908 79812
rect 132454 79766 132506 79772
rect 131948 79698 132000 79704
rect 132052 79716 132126 79744
rect 131684 79648 131758 79676
rect 131856 79688 131908 79694
rect 131684 76650 131712 79648
rect 131856 79630 131908 79636
rect 131762 78840 131818 78849
rect 131762 78775 131818 78784
rect 131776 78441 131804 78775
rect 131762 78432 131818 78441
rect 131762 78367 131818 78376
rect 131868 78282 131896 79630
rect 131776 78254 131896 78282
rect 131776 76838 131804 78254
rect 131764 76832 131816 76838
rect 131764 76774 131816 76780
rect 131684 76622 131804 76650
rect 131672 76356 131724 76362
rect 131672 76298 131724 76304
rect 131684 20058 131712 76298
rect 131776 71058 131804 76622
rect 131764 71052 131816 71058
rect 131764 70994 131816 71000
rect 131960 70394 131988 79698
rect 132052 75206 132080 79716
rect 132374 79676 132402 79750
rect 132684 79756 132736 79762
rect 132684 79698 132736 79704
rect 132222 79656 132278 79665
rect 132132 79620 132184 79626
rect 132222 79591 132278 79600
rect 132328 79648 132402 79676
rect 132592 79688 132644 79694
rect 132498 79656 132554 79665
rect 132132 79562 132184 79568
rect 132144 76362 132172 79562
rect 132236 76498 132264 79591
rect 132224 76492 132276 76498
rect 132224 76434 132276 76440
rect 132132 76356 132184 76362
rect 132132 76298 132184 76304
rect 132040 75200 132092 75206
rect 132040 75142 132092 75148
rect 131868 70366 131988 70394
rect 132328 70394 132356 79648
rect 132592 79630 132644 79636
rect 132498 79591 132554 79600
rect 132408 79552 132460 79558
rect 132408 79494 132460 79500
rect 132420 78334 132448 79494
rect 132408 78328 132460 78334
rect 132408 78270 132460 78276
rect 132512 78198 132540 79591
rect 132500 78192 132552 78198
rect 132500 78134 132552 78140
rect 132500 77308 132552 77314
rect 132500 77250 132552 77256
rect 132512 75342 132540 77250
rect 132500 75336 132552 75342
rect 132500 75278 132552 75284
rect 132328 70366 132448 70394
rect 131672 20052 131724 20058
rect 131672 19994 131724 20000
rect 131580 10532 131632 10538
rect 131580 10474 131632 10480
rect 131488 6384 131540 6390
rect 131488 6326 131540 6332
rect 131868 3874 131896 70366
rect 132420 5234 132448 70366
rect 132604 5302 132632 79630
rect 132696 75857 132724 79698
rect 132774 79656 132830 79665
rect 132774 79591 132830 79600
rect 132788 77790 132816 79591
rect 132880 79422 132908 79784
rect 132960 79756 133012 79762
rect 133110 79744 133138 80036
rect 133202 79830 133230 80036
rect 133294 79898 133322 80036
rect 133282 79892 133334 79898
rect 133282 79834 133334 79840
rect 133190 79824 133242 79830
rect 133190 79766 133242 79772
rect 133386 79744 133414 80036
rect 133478 79966 133506 80036
rect 133466 79960 133518 79966
rect 133466 79902 133518 79908
rect 133570 79830 133598 80036
rect 133662 79830 133690 80036
rect 133754 79937 133782 80036
rect 133846 79966 133874 80036
rect 133834 79960 133886 79966
rect 133740 79928 133796 79937
rect 133834 79902 133886 79908
rect 133938 79898 133966 80036
rect 134030 79937 134058 80036
rect 134122 79966 134150 80036
rect 134214 79966 134242 80036
rect 134110 79960 134162 79966
rect 134016 79928 134072 79937
rect 133740 79863 133796 79872
rect 133926 79892 133978 79898
rect 134110 79902 134162 79908
rect 134202 79960 134254 79966
rect 134306 79937 134334 80036
rect 134202 79902 134254 79908
rect 134292 79928 134348 79937
rect 134016 79863 134072 79872
rect 134398 79898 134426 80036
rect 134490 79971 134518 80036
rect 134476 79962 134532 79971
rect 134582 79966 134610 80036
rect 134292 79863 134348 79872
rect 134386 79892 134438 79898
rect 134476 79897 134532 79906
rect 134570 79960 134622 79966
rect 134570 79902 134622 79908
rect 134674 79898 134702 80036
rect 134766 79898 134794 80036
rect 134858 79966 134886 80036
rect 134846 79960 134898 79966
rect 134950 79937 134978 80036
rect 135042 79966 135070 80036
rect 135134 79966 135162 80036
rect 135030 79960 135082 79966
rect 134846 79902 134898 79908
rect 134936 79928 134992 79937
rect 133926 79834 133978 79840
rect 134386 79834 134438 79840
rect 134662 79892 134714 79898
rect 134662 79834 134714 79840
rect 134754 79892 134806 79898
rect 135030 79902 135082 79908
rect 135122 79960 135174 79966
rect 135122 79902 135174 79908
rect 134936 79863 134992 79872
rect 134754 79834 134806 79840
rect 133558 79824 133610 79830
rect 133558 79766 133610 79772
rect 133650 79824 133702 79830
rect 133650 79766 133702 79772
rect 134248 79824 134300 79830
rect 135226 79812 135254 80036
rect 134248 79766 134300 79772
rect 135180 79784 135254 79812
rect 133012 79716 133138 79744
rect 133340 79716 133414 79744
rect 133788 79756 133840 79762
rect 132960 79698 133012 79704
rect 132972 79614 133184 79642
rect 132868 79416 132920 79422
rect 132868 79358 132920 79364
rect 132776 77784 132828 77790
rect 132776 77726 132828 77732
rect 132972 76888 133000 79614
rect 133156 79608 133184 79614
rect 133236 79620 133288 79626
rect 133156 79580 133236 79608
rect 133236 79562 133288 79568
rect 133052 79552 133104 79558
rect 133052 79494 133104 79500
rect 132880 76860 133000 76888
rect 132774 76664 132830 76673
rect 132774 76599 132830 76608
rect 132682 75848 132738 75857
rect 132682 75783 132738 75792
rect 132684 75676 132736 75682
rect 132684 75618 132736 75624
rect 132696 6594 132724 75618
rect 132788 7886 132816 76599
rect 132776 7880 132828 7886
rect 132776 7822 132828 7828
rect 132880 7818 132908 76860
rect 133064 76786 133092 79494
rect 133236 79484 133288 79490
rect 133236 79426 133288 79432
rect 133144 79416 133196 79422
rect 133144 79358 133196 79364
rect 132972 76758 133092 76786
rect 132972 10606 133000 76758
rect 133052 76696 133104 76702
rect 133052 76638 133104 76644
rect 133064 10674 133092 76638
rect 133156 74050 133184 79358
rect 133248 76770 133276 79426
rect 133236 76764 133288 76770
rect 133236 76706 133288 76712
rect 133144 74044 133196 74050
rect 133144 73986 133196 73992
rect 133340 70394 133368 79716
rect 133788 79698 133840 79704
rect 133880 79756 133932 79762
rect 133880 79698 133932 79704
rect 133972 79756 134024 79762
rect 133972 79698 134024 79704
rect 133604 79688 133656 79694
rect 133604 79630 133656 79636
rect 133420 79552 133472 79558
rect 133420 79494 133472 79500
rect 133432 77926 133460 79494
rect 133512 78260 133564 78266
rect 133512 78202 133564 78208
rect 133420 77920 133472 77926
rect 133420 77862 133472 77868
rect 133420 76968 133472 76974
rect 133420 76910 133472 76916
rect 133432 75070 133460 76910
rect 133420 75064 133472 75070
rect 133420 75006 133472 75012
rect 133156 70366 133368 70394
rect 133524 70394 133552 78202
rect 133616 75682 133644 79630
rect 133800 76702 133828 79698
rect 133892 77314 133920 79698
rect 133880 77308 133932 77314
rect 133880 77250 133932 77256
rect 133880 76764 133932 76770
rect 133880 76706 133932 76712
rect 133788 76696 133840 76702
rect 133788 76638 133840 76644
rect 133604 75676 133656 75682
rect 133604 75618 133656 75624
rect 133524 70366 133828 70394
rect 133052 10668 133104 10674
rect 133052 10610 133104 10616
rect 132960 10600 133012 10606
rect 132960 10542 133012 10548
rect 132868 7812 132920 7818
rect 132868 7754 132920 7760
rect 132684 6588 132736 6594
rect 132684 6530 132736 6536
rect 133156 5370 133184 70366
rect 133144 5364 133196 5370
rect 133144 5306 133196 5312
rect 132592 5296 132644 5302
rect 132592 5238 132644 5244
rect 132408 5228 132460 5234
rect 132408 5170 132460 5176
rect 131856 3868 131908 3874
rect 131856 3810 131908 3816
rect 130660 3732 130712 3738
rect 130660 3674 130712 3680
rect 133800 3602 133828 70366
rect 130384 3596 130436 3602
rect 130384 3538 130436 3544
rect 133788 3596 133840 3602
rect 133788 3538 133840 3544
rect 131764 3528 131816 3534
rect 129844 3454 130608 3482
rect 131764 3470 131816 3476
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 128372 462 128952 490
rect 130580 480 130608 3454
rect 131776 480 131804 3470
rect 132960 3120 133012 3126
rect 132960 3062 133012 3068
rect 132972 480 133000 3062
rect 128924 354 128952 462
rect 129342 354 129454 480
rect 128924 326 129454 354
rect 129342 -960 129454 326
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 133892 354 133920 76706
rect 133984 76673 134012 79698
rect 134064 79552 134116 79558
rect 134064 79494 134116 79500
rect 133970 76664 134026 76673
rect 133970 76599 134026 76608
rect 134076 73154 134104 79494
rect 134260 77081 134288 79766
rect 134616 79756 134668 79762
rect 134616 79698 134668 79704
rect 134708 79756 134760 79762
rect 134708 79698 134760 79704
rect 134800 79756 134852 79762
rect 134800 79698 134852 79704
rect 134340 79620 134392 79626
rect 134340 79562 134392 79568
rect 134246 77072 134302 77081
rect 134246 77007 134302 77016
rect 134352 76922 134380 79562
rect 134524 77988 134576 77994
rect 134524 77930 134576 77936
rect 133984 73126 134104 73154
rect 134168 76894 134380 76922
rect 133984 70394 134012 73126
rect 133984 70366 134104 70394
rect 134076 7954 134104 70366
rect 134168 14550 134196 76894
rect 134248 76832 134300 76838
rect 134248 76774 134300 76780
rect 134260 18766 134288 76774
rect 134432 76628 134484 76634
rect 134432 76570 134484 76576
rect 134444 70394 134472 76570
rect 134352 70366 134472 70394
rect 134352 21418 134380 70366
rect 134340 21412 134392 21418
rect 134340 21354 134392 21360
rect 134248 18760 134300 18766
rect 134248 18702 134300 18708
rect 134156 14544 134208 14550
rect 134156 14486 134208 14492
rect 134064 7948 134116 7954
rect 134064 7890 134116 7896
rect 134536 4146 134564 77930
rect 134628 76838 134656 79698
rect 134616 76832 134668 76838
rect 134616 76774 134668 76780
rect 134614 76664 134670 76673
rect 134614 76599 134670 76608
rect 134628 70394 134656 76599
rect 134720 74118 134748 79698
rect 134812 77042 134840 79698
rect 134984 79688 135036 79694
rect 134984 79630 135036 79636
rect 135076 79688 135128 79694
rect 135076 79630 135128 79636
rect 134892 79416 134944 79422
rect 134892 79358 134944 79364
rect 134904 77382 134932 79358
rect 134892 77376 134944 77382
rect 134892 77318 134944 77324
rect 134800 77036 134852 77042
rect 134800 76978 134852 76984
rect 134996 75750 135024 79630
rect 135088 76906 135116 79630
rect 135076 76900 135128 76906
rect 135076 76842 135128 76848
rect 135180 76634 135208 79784
rect 135318 79744 135346 80036
rect 135272 79716 135346 79744
rect 135272 77994 135300 79716
rect 135410 79676 135438 80036
rect 135502 79937 135530 80036
rect 135594 79966 135622 80036
rect 135686 79966 135714 80036
rect 135582 79960 135634 79966
rect 135488 79928 135544 79937
rect 135582 79902 135634 79908
rect 135674 79960 135726 79966
rect 135674 79902 135726 79908
rect 135488 79863 135544 79872
rect 135778 79830 135806 80036
rect 135870 79971 135898 80036
rect 135856 79962 135912 79971
rect 135856 79897 135912 79906
rect 135962 79898 135990 80036
rect 136054 79966 136082 80036
rect 136146 79966 136174 80036
rect 136238 79966 136266 80036
rect 136330 79966 136358 80036
rect 136422 79971 136450 80036
rect 136042 79960 136094 79966
rect 136042 79902 136094 79908
rect 136134 79960 136186 79966
rect 136134 79902 136186 79908
rect 136226 79960 136278 79966
rect 136226 79902 136278 79908
rect 136318 79960 136370 79966
rect 136318 79902 136370 79908
rect 136408 79962 136464 79971
rect 136514 79966 136542 80036
rect 136606 79971 136634 80036
rect 135950 79892 136002 79898
rect 136408 79897 136464 79906
rect 136502 79960 136554 79966
rect 136502 79902 136554 79908
rect 136592 79962 136648 79971
rect 136592 79897 136648 79906
rect 135950 79834 136002 79840
rect 135766 79824 135818 79830
rect 135766 79766 135818 79772
rect 136456 79824 136508 79830
rect 136456 79766 136508 79772
rect 136546 79792 136602 79801
rect 135996 79756 136048 79762
rect 135996 79698 136048 79704
rect 136088 79756 136140 79762
rect 136088 79698 136140 79704
rect 135364 79648 135438 79676
rect 135536 79688 135588 79694
rect 135260 77988 135312 77994
rect 135260 77930 135312 77936
rect 135364 77874 135392 79648
rect 135720 79688 135772 79694
rect 135536 79630 135588 79636
rect 135626 79656 135682 79665
rect 135272 77846 135392 77874
rect 135168 76628 135220 76634
rect 135168 76570 135220 76576
rect 134984 75744 135036 75750
rect 134984 75686 135036 75692
rect 135272 74497 135300 77846
rect 135548 76974 135576 79630
rect 135720 79630 135772 79636
rect 135626 79591 135682 79600
rect 135536 76968 135588 76974
rect 135536 76910 135588 76916
rect 135640 76752 135668 79591
rect 135456 76724 135668 76752
rect 135352 76220 135404 76226
rect 135352 76162 135404 76168
rect 135258 74488 135314 74497
rect 135258 74423 135314 74432
rect 134708 74112 134760 74118
rect 134708 74054 134760 74060
rect 134628 70366 134748 70394
rect 134720 6662 134748 70366
rect 135364 6914 135392 76162
rect 135272 6886 135392 6914
rect 134708 6656 134760 6662
rect 134708 6598 134760 6604
rect 134524 4140 134576 4146
rect 134524 4082 134576 4088
rect 135272 480 135300 6886
rect 135456 3126 135484 76724
rect 135534 76664 135590 76673
rect 135732 76650 135760 79630
rect 135904 79620 135956 79626
rect 135904 79562 135956 79568
rect 135812 79552 135864 79558
rect 135812 79494 135864 79500
rect 135534 76599 135590 76608
rect 135640 76622 135760 76650
rect 135548 3194 135576 76599
rect 135640 3534 135668 76622
rect 135720 73908 135772 73914
rect 135720 73850 135772 73856
rect 135628 3528 135680 3534
rect 135628 3470 135680 3476
rect 135732 3330 135760 73850
rect 135720 3324 135772 3330
rect 135720 3266 135772 3272
rect 135536 3188 135588 3194
rect 135536 3130 135588 3136
rect 135824 3126 135852 79494
rect 135916 76770 135944 79562
rect 135904 76764 135956 76770
rect 135904 76706 135956 76712
rect 135904 76628 135956 76634
rect 135904 76570 135956 76576
rect 135444 3120 135496 3126
rect 135444 3062 135496 3068
rect 135812 3120 135864 3126
rect 135812 3062 135864 3068
rect 135916 3058 135944 76570
rect 136008 76226 136036 79698
rect 135996 76220 136048 76226
rect 135996 76162 136048 76168
rect 135996 75744 136048 75750
rect 135996 75686 136048 75692
rect 136008 45014 136036 75686
rect 135996 45008 136048 45014
rect 135996 44950 136048 44956
rect 136100 16574 136128 79698
rect 136364 79620 136416 79626
rect 136364 79562 136416 79568
rect 136376 73914 136404 79562
rect 136468 76634 136496 79766
rect 136546 79727 136602 79736
rect 136698 79744 136726 80036
rect 136790 79966 136818 80036
rect 136778 79960 136830 79966
rect 136778 79902 136830 79908
rect 136882 79898 136910 80036
rect 136870 79892 136922 79898
rect 136870 79834 136922 79840
rect 136974 79830 137002 80036
rect 137066 79971 137094 80036
rect 137052 79962 137108 79971
rect 137158 79966 137186 80036
rect 137250 79966 137278 80036
rect 137052 79897 137108 79906
rect 137146 79960 137198 79966
rect 137146 79902 137198 79908
rect 137238 79960 137290 79966
rect 137238 79902 137290 79908
rect 137342 79898 137370 80036
rect 137330 79892 137382 79898
rect 137330 79834 137382 79840
rect 136962 79824 137014 79830
rect 136962 79766 137014 79772
rect 137100 79824 137152 79830
rect 137100 79766 137152 79772
rect 136456 76628 136508 76634
rect 136456 76570 136508 76576
rect 136560 75750 136588 79727
rect 136698 79716 136864 79744
rect 136640 79620 136692 79626
rect 136640 79562 136692 79568
rect 136652 76634 136680 79562
rect 136732 79484 136784 79490
rect 136732 79426 136784 79432
rect 136640 76628 136692 76634
rect 136640 76570 136692 76576
rect 136548 75744 136600 75750
rect 136548 75686 136600 75692
rect 136364 73908 136416 73914
rect 136364 73850 136416 73856
rect 136100 16546 136496 16574
rect 135904 3052 135956 3058
rect 135904 2994 135956 3000
rect 136468 480 136496 16546
rect 136744 3670 136772 79426
rect 136836 78130 136864 79716
rect 136916 79688 136968 79694
rect 136916 79630 136968 79636
rect 137008 79688 137060 79694
rect 137008 79630 137060 79636
rect 136928 78266 136956 79630
rect 137020 79540 137048 79630
rect 137112 79608 137140 79766
rect 137434 79744 137462 80036
rect 137296 79716 137462 79744
rect 137526 79744 137554 80036
rect 137618 79898 137646 80036
rect 137710 79971 137738 80036
rect 137696 79962 137752 79971
rect 137606 79892 137658 79898
rect 137696 79897 137752 79906
rect 137606 79834 137658 79840
rect 137802 79778 137830 80036
rect 137894 79830 137922 80036
rect 137986 79898 138014 80036
rect 138078 79966 138106 80036
rect 138170 79966 138198 80036
rect 138262 79971 138290 80036
rect 138066 79960 138118 79966
rect 138066 79902 138118 79908
rect 138158 79960 138210 79966
rect 138158 79902 138210 79908
rect 138248 79962 138304 79971
rect 137974 79892 138026 79898
rect 138248 79897 138304 79906
rect 138354 79898 138382 80036
rect 138446 79966 138474 80036
rect 138434 79960 138486 79966
rect 138434 79902 138486 79908
rect 137974 79834 138026 79840
rect 138342 79892 138394 79898
rect 138342 79834 138394 79840
rect 137756 79750 137830 79778
rect 137882 79824 137934 79830
rect 138538 79812 138566 80036
rect 138630 79971 138658 80036
rect 138616 79962 138672 79971
rect 138722 79966 138750 80036
rect 138814 79966 138842 80036
rect 138906 79966 138934 80036
rect 138616 79897 138672 79906
rect 138710 79960 138762 79966
rect 138710 79902 138762 79908
rect 138802 79960 138854 79966
rect 138802 79902 138854 79908
rect 138894 79960 138946 79966
rect 138894 79902 138946 79908
rect 137882 79766 137934 79772
rect 138492 79784 138566 79812
rect 138998 79801 139026 80036
rect 139090 79812 139118 80036
rect 139182 79966 139210 80036
rect 139274 79966 139302 80036
rect 139366 79971 139394 80036
rect 139170 79960 139222 79966
rect 139170 79902 139222 79908
rect 139262 79960 139314 79966
rect 139262 79902 139314 79908
rect 139352 79962 139408 79971
rect 139352 79897 139408 79906
rect 139458 79898 139486 80036
rect 139550 79937 139578 80036
rect 139536 79928 139592 79937
rect 139446 79892 139498 79898
rect 139536 79863 139592 79872
rect 139446 79834 139498 79840
rect 139216 79824 139268 79830
rect 139090 79801 139164 79812
rect 138984 79792 139040 79801
rect 138388 79756 138440 79762
rect 137756 79744 137784 79750
rect 137526 79716 137600 79744
rect 137112 79580 137232 79608
rect 137020 79512 137140 79540
rect 137112 78674 137140 79512
rect 137204 78928 137232 79580
rect 137296 79490 137324 79716
rect 137376 79620 137428 79626
rect 137376 79562 137428 79568
rect 137468 79620 137520 79626
rect 137468 79562 137520 79568
rect 137284 79484 137336 79490
rect 137284 79426 137336 79432
rect 137204 78900 137324 78928
rect 137020 78646 137140 78674
rect 137192 78668 137244 78674
rect 136916 78260 136968 78266
rect 136916 78202 136968 78208
rect 136914 78160 136970 78169
rect 136824 78124 136876 78130
rect 136914 78095 136970 78104
rect 136824 78066 136876 78072
rect 136824 76628 136876 76634
rect 136824 76570 136876 76576
rect 136836 3942 136864 76570
rect 136928 5098 136956 78095
rect 136916 5092 136968 5098
rect 136916 5034 136968 5040
rect 137020 4962 137048 78646
rect 137192 78610 137244 78616
rect 137100 76628 137152 76634
rect 137100 76570 137152 76576
rect 137008 4956 137060 4962
rect 137008 4898 137060 4904
rect 137112 4894 137140 76570
rect 137204 60042 137232 78610
rect 137296 66230 137324 78900
rect 137388 73234 137416 79562
rect 137480 78674 137508 79562
rect 137468 78668 137520 78674
rect 137468 78610 137520 78616
rect 137468 78124 137520 78130
rect 137468 78066 137520 78072
rect 137480 73506 137508 78066
rect 137468 73500 137520 73506
rect 137468 73442 137520 73448
rect 137376 73228 137428 73234
rect 137376 73170 137428 73176
rect 137572 70394 137600 79716
rect 137710 79716 137784 79744
rect 137710 79642 137738 79716
rect 138388 79698 138440 79704
rect 138202 79656 138258 79665
rect 137710 79614 137784 79642
rect 137652 79484 137704 79490
rect 137652 79426 137704 79432
rect 137664 76022 137692 79426
rect 137756 76634 137784 79614
rect 138202 79591 138258 79600
rect 138296 79620 138348 79626
rect 137928 79552 137980 79558
rect 137928 79494 137980 79500
rect 138020 79552 138072 79558
rect 138020 79494 138072 79500
rect 137836 79484 137888 79490
rect 137836 79426 137888 79432
rect 137848 76809 137876 79426
rect 137834 76800 137890 76809
rect 137834 76735 137890 76744
rect 137940 76673 137968 79494
rect 137926 76664 137982 76673
rect 137744 76628 137796 76634
rect 137926 76599 137982 76608
rect 137744 76570 137796 76576
rect 138032 76537 138060 79494
rect 138112 79484 138164 79490
rect 138112 79426 138164 79432
rect 138018 76528 138074 76537
rect 138018 76463 138074 76472
rect 137652 76016 137704 76022
rect 137652 75958 137704 75964
rect 138020 75404 138072 75410
rect 138020 75346 138072 75352
rect 137572 70366 137784 70394
rect 137284 66224 137336 66230
rect 137284 66166 137336 66172
rect 137192 60036 137244 60042
rect 137192 59978 137244 59984
rect 137100 4888 137152 4894
rect 137100 4830 137152 4836
rect 136824 3936 136876 3942
rect 136824 3878 136876 3884
rect 137756 3738 137784 70366
rect 138032 5234 138060 75346
rect 138020 5228 138072 5234
rect 138020 5170 138072 5176
rect 138124 4826 138152 79426
rect 138216 75138 138244 79591
rect 138296 79562 138348 79568
rect 138204 75132 138256 75138
rect 138204 75074 138256 75080
rect 138204 74996 138256 75002
rect 138204 74938 138256 74944
rect 138216 5030 138244 74938
rect 138308 6186 138336 79562
rect 138400 75274 138428 79698
rect 138388 75268 138440 75274
rect 138388 75210 138440 75216
rect 138388 75132 138440 75138
rect 138388 75074 138440 75080
rect 138400 20126 138428 75074
rect 138492 44878 138520 79784
rect 139090 79792 139178 79801
rect 139090 79784 139122 79792
rect 138984 79727 139040 79736
rect 139216 79766 139268 79772
rect 139352 79792 139408 79801
rect 139122 79727 139178 79736
rect 138572 79688 138624 79694
rect 139032 79688 139084 79694
rect 138572 79630 138624 79636
rect 138938 79656 138994 79665
rect 138584 75410 138612 79630
rect 138848 79620 138900 79626
rect 139032 79630 139084 79636
rect 139124 79688 139176 79694
rect 139124 79630 139176 79636
rect 138938 79591 138994 79600
rect 138848 79562 138900 79568
rect 138664 79552 138716 79558
rect 138664 79494 138716 79500
rect 138572 75404 138624 75410
rect 138572 75346 138624 75352
rect 138572 75268 138624 75274
rect 138572 75210 138624 75216
rect 138584 66162 138612 75210
rect 138676 75002 138704 79494
rect 138860 78826 138888 79562
rect 138768 78798 138888 78826
rect 138664 74996 138716 75002
rect 138664 74938 138716 74944
rect 138768 70394 138796 78798
rect 138952 78690 138980 79591
rect 139044 79218 139072 79630
rect 139032 79212 139084 79218
rect 139032 79154 139084 79160
rect 139136 78713 139164 79630
rect 138860 78662 138980 78690
rect 139122 78704 139178 78713
rect 138860 71058 138888 78662
rect 139122 78639 139178 78648
rect 139228 78606 139256 79766
rect 139320 79736 139352 79744
rect 139320 79727 139408 79736
rect 139490 79792 139546 79801
rect 139490 79727 139546 79736
rect 139642 79744 139670 80036
rect 139734 79937 139762 80036
rect 139826 79966 139854 80036
rect 139814 79960 139866 79966
rect 139720 79928 139776 79937
rect 139814 79902 139866 79908
rect 139918 79898 139946 80036
rect 139720 79863 139776 79872
rect 139906 79892 139958 79898
rect 139906 79834 139958 79840
rect 140010 79830 140038 80036
rect 139998 79824 140050 79830
rect 139998 79766 140050 79772
rect 140102 79778 140130 80036
rect 140194 79966 140222 80036
rect 140286 79966 140314 80036
rect 140378 79966 140406 80036
rect 140182 79960 140234 79966
rect 140182 79902 140234 79908
rect 140274 79960 140326 79966
rect 140274 79902 140326 79908
rect 140366 79960 140418 79966
rect 140366 79902 140418 79908
rect 140470 79801 140498 80036
rect 140562 79971 140590 80036
rect 140548 79962 140604 79971
rect 140548 79897 140604 79906
rect 140654 79898 140682 80036
rect 140642 79892 140694 79898
rect 140642 79834 140694 79840
rect 140456 79792 140512 79801
rect 139860 79756 139912 79762
rect 139320 79716 139394 79727
rect 139216 78600 139268 78606
rect 139320 78577 139348 79716
rect 139400 79620 139452 79626
rect 139400 79562 139452 79568
rect 139216 78542 139268 78548
rect 139306 78568 139362 78577
rect 139306 78503 139362 78512
rect 139412 77382 139440 79562
rect 139400 77376 139452 77382
rect 139400 77318 139452 77324
rect 139400 75948 139452 75954
rect 139400 75890 139452 75896
rect 138940 73500 138992 73506
rect 138940 73442 138992 73448
rect 138848 71052 138900 71058
rect 138848 70994 138900 71000
rect 138676 70378 138796 70394
rect 138664 70372 138796 70378
rect 138716 70366 138796 70372
rect 138664 70314 138716 70320
rect 138572 66156 138624 66162
rect 138572 66098 138624 66104
rect 138664 60036 138716 60042
rect 138664 59978 138716 59984
rect 138480 44872 138532 44878
rect 138480 44814 138532 44820
rect 138388 20120 138440 20126
rect 138388 20062 138440 20068
rect 138296 6180 138348 6186
rect 138296 6122 138348 6128
rect 138204 5024 138256 5030
rect 138204 4966 138256 4972
rect 138112 4820 138164 4826
rect 138112 4762 138164 4768
rect 138676 4078 138704 59978
rect 138952 4418 138980 73442
rect 139412 27198 139440 75890
rect 139504 27266 139532 79727
rect 139642 79716 139808 79744
rect 139584 79552 139636 79558
rect 139584 79494 139636 79500
rect 139596 75954 139624 79494
rect 139584 75948 139636 75954
rect 139584 75890 139636 75896
rect 139676 75812 139728 75818
rect 139676 75754 139728 75760
rect 139584 75744 139636 75750
rect 139584 75686 139636 75692
rect 139596 28490 139624 75686
rect 139688 34134 139716 75754
rect 139780 46238 139808 79716
rect 140102 79750 140176 79778
rect 139860 79698 139912 79704
rect 139872 61538 139900 79698
rect 139952 79688 140004 79694
rect 140148 79676 140176 79750
rect 140746 79778 140774 80036
rect 140838 79966 140866 80036
rect 140930 79966 140958 80036
rect 140826 79960 140878 79966
rect 140826 79902 140878 79908
rect 140918 79960 140970 79966
rect 140918 79902 140970 79908
rect 141022 79778 141050 80036
rect 141114 79830 141142 80036
rect 141206 79898 141234 80036
rect 141298 79937 141326 80036
rect 141390 79966 141418 80036
rect 141482 79966 141510 80036
rect 141574 79966 141602 80036
rect 141378 79960 141430 79966
rect 141284 79928 141340 79937
rect 141194 79892 141246 79898
rect 141378 79902 141430 79908
rect 141470 79960 141522 79966
rect 141470 79902 141522 79908
rect 141562 79960 141614 79966
rect 141562 79902 141614 79908
rect 141284 79863 141340 79872
rect 141194 79834 141246 79840
rect 140456 79727 140512 79736
rect 140608 79750 140774 79778
rect 140976 79750 141050 79778
rect 141102 79824 141154 79830
rect 141102 79766 141154 79772
rect 141238 79792 141294 79801
rect 140102 79648 140176 79676
rect 140412 79688 140464 79694
rect 140102 79642 140130 79648
rect 139952 79630 140004 79636
rect 139964 76106 139992 79630
rect 140056 79614 140130 79642
rect 140412 79630 140464 79636
rect 140320 79620 140372 79626
rect 140056 76242 140084 79614
rect 140240 79580 140320 79608
rect 140240 78674 140268 79580
rect 140320 79562 140372 79568
rect 140320 79484 140372 79490
rect 140320 79426 140372 79432
rect 140148 78646 140268 78674
rect 140148 76401 140176 78646
rect 140228 76764 140280 76770
rect 140228 76706 140280 76712
rect 140134 76392 140190 76401
rect 140134 76327 140190 76336
rect 140056 76214 140176 76242
rect 139964 76078 140084 76106
rect 139952 75948 140004 75954
rect 139952 75890 140004 75896
rect 139964 67454 139992 75890
rect 140056 68678 140084 76078
rect 140148 75750 140176 76214
rect 140240 75954 140268 76706
rect 140228 75948 140280 75954
rect 140228 75890 140280 75896
rect 140332 75818 140360 79426
rect 140424 76770 140452 79630
rect 140504 79416 140556 79422
rect 140504 79358 140556 79364
rect 140516 78946 140544 79358
rect 140504 78940 140556 78946
rect 140504 78882 140556 78888
rect 140504 78600 140556 78606
rect 140504 78542 140556 78548
rect 140412 76764 140464 76770
rect 140412 76706 140464 76712
rect 140410 76664 140466 76673
rect 140410 76599 140466 76608
rect 140320 75812 140372 75818
rect 140320 75754 140372 75760
rect 140136 75744 140188 75750
rect 140136 75686 140188 75692
rect 140044 68672 140096 68678
rect 140044 68614 140096 68620
rect 139952 67448 140004 67454
rect 139952 67390 140004 67396
rect 140044 66224 140096 66230
rect 140044 66166 140096 66172
rect 139860 61532 139912 61538
rect 139860 61474 139912 61480
rect 139768 46232 139820 46238
rect 139768 46174 139820 46180
rect 139676 34128 139728 34134
rect 139676 34070 139728 34076
rect 139584 28484 139636 28490
rect 139584 28426 139636 28432
rect 139492 27260 139544 27266
rect 139492 27202 139544 27208
rect 139400 27192 139452 27198
rect 139400 27134 139452 27140
rect 138940 4412 138992 4418
rect 138940 4354 138992 4360
rect 138664 4072 138716 4078
rect 138664 4014 138716 4020
rect 140056 3806 140084 66166
rect 140424 6254 140452 76599
rect 140516 27334 140544 78542
rect 140608 74089 140636 79750
rect 140688 79688 140740 79694
rect 140688 79630 140740 79636
rect 140872 79688 140924 79694
rect 140872 79630 140924 79636
rect 140700 78538 140728 79630
rect 140780 79620 140832 79626
rect 140780 79562 140832 79568
rect 140688 78532 140740 78538
rect 140688 78474 140740 78480
rect 140594 74080 140650 74089
rect 140594 74015 140650 74024
rect 140792 28422 140820 79562
rect 140884 78130 140912 79630
rect 140872 78124 140924 78130
rect 140872 78066 140924 78072
rect 140976 75970 141004 79750
rect 141666 79778 141694 80036
rect 141758 79898 141786 80036
rect 141850 79937 141878 80036
rect 141942 79966 141970 80036
rect 141930 79960 141982 79966
rect 141836 79928 141892 79937
rect 141746 79892 141798 79898
rect 141930 79902 141982 79908
rect 142034 79898 142062 80036
rect 141836 79863 141892 79872
rect 142022 79892 142074 79898
rect 141746 79834 141798 79840
rect 142022 79834 142074 79840
rect 141666 79750 141740 79778
rect 141238 79727 141294 79736
rect 141056 79688 141108 79694
rect 141056 79630 141108 79636
rect 141146 79656 141202 79665
rect 141068 78470 141096 79630
rect 141146 79591 141202 79600
rect 141160 79082 141188 79591
rect 141148 79076 141200 79082
rect 141148 79018 141200 79024
rect 141056 78464 141108 78470
rect 141056 78406 141108 78412
rect 140976 75942 141096 75970
rect 140964 75880 141016 75886
rect 140964 75822 141016 75828
rect 140872 75268 140924 75274
rect 140872 75210 140924 75216
rect 140884 30054 140912 75210
rect 140976 30122 141004 75822
rect 141068 34066 141096 75942
rect 141148 75948 141200 75954
rect 141148 75890 141200 75896
rect 141056 34060 141108 34066
rect 141056 34002 141108 34008
rect 141160 33930 141188 75890
rect 141252 33998 141280 79727
rect 141332 79688 141384 79694
rect 141608 79688 141660 79694
rect 141384 79648 141464 79676
rect 141332 79630 141384 79636
rect 141332 79348 141384 79354
rect 141332 79290 141384 79296
rect 141344 65890 141372 79290
rect 141436 65958 141464 79648
rect 141608 79630 141660 79636
rect 141516 79620 141568 79626
rect 141516 79562 141568 79568
rect 141528 75886 141556 79562
rect 141620 75954 141648 79630
rect 141712 79354 141740 79750
rect 141792 79756 141844 79762
rect 141792 79698 141844 79704
rect 141700 79348 141752 79354
rect 141700 79290 141752 79296
rect 141700 79076 141752 79082
rect 141700 79018 141752 79024
rect 141712 77722 141740 79018
rect 141700 77716 141752 77722
rect 141700 77658 141752 77664
rect 141608 75948 141660 75954
rect 141608 75890 141660 75896
rect 141516 75880 141568 75886
rect 141516 75822 141568 75828
rect 141804 75274 141832 79698
rect 142126 79676 142154 80036
rect 142218 79966 142246 80036
rect 142310 79966 142338 80036
rect 142206 79960 142258 79966
rect 142206 79902 142258 79908
rect 142298 79960 142350 79966
rect 142298 79902 142350 79908
rect 142402 79812 142430 80036
rect 142494 79966 142522 80036
rect 142482 79960 142534 79966
rect 142482 79902 142534 79908
rect 142356 79784 142430 79812
rect 142252 79756 142304 79762
rect 142252 79698 142304 79704
rect 141974 79656 142030 79665
rect 141884 79620 141936 79626
rect 141974 79591 142030 79600
rect 142080 79648 142154 79676
rect 141884 79562 141936 79568
rect 141792 75268 141844 75274
rect 141792 75210 141844 75216
rect 141896 70394 141924 79562
rect 141988 79286 142016 79591
rect 141976 79280 142028 79286
rect 141976 79222 142028 79228
rect 141974 78568 142030 78577
rect 141974 78503 142030 78512
rect 141988 75585 142016 78503
rect 142080 75993 142108 79648
rect 142160 79348 142212 79354
rect 142160 79290 142212 79296
rect 142172 77081 142200 79290
rect 142158 77072 142214 77081
rect 142158 77007 142214 77016
rect 142066 75984 142122 75993
rect 142066 75919 142122 75928
rect 142264 75914 142292 79698
rect 142356 76158 142384 79784
rect 142436 79688 142488 79694
rect 142436 79630 142488 79636
rect 142448 76242 142476 79630
rect 142586 79608 142614 80036
rect 142678 79898 142706 80036
rect 142770 79937 142798 80036
rect 142756 79928 142812 79937
rect 142666 79892 142718 79898
rect 142862 79898 142890 80036
rect 142756 79863 142812 79872
rect 142850 79892 142902 79898
rect 142666 79834 142718 79840
rect 142850 79834 142902 79840
rect 142954 79830 142982 80036
rect 142942 79824 142994 79830
rect 142756 79792 142812 79801
rect 142678 79736 142756 79744
rect 142942 79766 142994 79772
rect 142678 79727 142812 79736
rect 142678 79716 142798 79727
rect 142678 79676 142706 79716
rect 142896 79688 142948 79694
rect 142678 79648 142752 79676
rect 142586 79580 142660 79608
rect 142448 76214 142568 76242
rect 142344 76152 142396 76158
rect 142344 76094 142396 76100
rect 142436 76084 142488 76090
rect 142436 76026 142488 76032
rect 142264 75886 142384 75914
rect 142160 75880 142212 75886
rect 142160 75822 142212 75828
rect 141974 75576 142030 75585
rect 141974 75511 142030 75520
rect 141528 70366 141924 70394
rect 141528 70106 141556 70366
rect 141516 70100 141568 70106
rect 141516 70042 141568 70048
rect 141516 66156 141568 66162
rect 141516 66098 141568 66104
rect 141424 65952 141476 65958
rect 141424 65894 141476 65900
rect 141332 65884 141384 65890
rect 141332 65826 141384 65832
rect 141240 33992 141292 33998
rect 141240 33934 141292 33940
rect 141148 33924 141200 33930
rect 141148 33866 141200 33872
rect 140964 30116 141016 30122
rect 140964 30058 141016 30064
rect 140872 30048 140924 30054
rect 140872 29990 140924 29996
rect 140780 28416 140832 28422
rect 140780 28358 140832 28364
rect 140504 27328 140556 27334
rect 140504 27270 140556 27276
rect 140412 6248 140464 6254
rect 140412 6190 140464 6196
rect 140044 3800 140096 3806
rect 140044 3742 140096 3748
rect 137744 3732 137796 3738
rect 137744 3674 137796 3680
rect 136732 3664 136784 3670
rect 136732 3606 136784 3612
rect 141528 3534 141556 66098
rect 142172 5166 142200 75822
rect 142252 73976 142304 73982
rect 142252 73918 142304 73924
rect 142264 7954 142292 73918
rect 142356 24614 142384 75886
rect 142344 24608 142396 24614
rect 142344 24550 142396 24556
rect 142448 24546 142476 76026
rect 142540 75818 142568 76214
rect 142632 76090 142660 79580
rect 142620 76084 142672 76090
rect 142620 76026 142672 76032
rect 142724 75914 142752 79648
rect 143046 79676 143074 80036
rect 143138 79835 143166 80036
rect 143230 79966 143258 80036
rect 143322 79966 143350 80036
rect 143414 79971 143442 80036
rect 143218 79960 143270 79966
rect 143218 79902 143270 79908
rect 143310 79960 143362 79966
rect 143310 79902 143362 79908
rect 143400 79962 143456 79971
rect 143506 79966 143534 80036
rect 143598 79966 143626 80036
rect 143400 79897 143456 79906
rect 143494 79960 143546 79966
rect 143494 79902 143546 79908
rect 143586 79960 143638 79966
rect 143586 79902 143638 79908
rect 143690 79898 143718 80036
rect 143678 79892 143730 79898
rect 143124 79826 143180 79835
rect 143678 79834 143730 79840
rect 143124 79761 143180 79770
rect 143356 79824 143408 79830
rect 143356 79766 143408 79772
rect 143630 79792 143686 79801
rect 143264 79688 143316 79694
rect 143046 79648 143120 79676
rect 142896 79630 142948 79636
rect 142804 79620 142856 79626
rect 142804 79562 142856 79568
rect 142632 75886 142752 75914
rect 142816 75886 142844 79562
rect 142528 75812 142580 75818
rect 142528 75754 142580 75760
rect 142528 75132 142580 75138
rect 142528 75074 142580 75080
rect 142540 26042 142568 75074
rect 142632 65822 142660 75886
rect 142804 75880 142856 75886
rect 142804 75822 142856 75828
rect 142712 75812 142764 75818
rect 142712 75754 142764 75760
rect 142724 68610 142752 75754
rect 142908 75138 142936 79630
rect 142988 79552 143040 79558
rect 142988 79494 143040 79500
rect 142896 75132 142948 75138
rect 142896 75074 142948 75080
rect 143000 74118 143028 79494
rect 142988 74112 143040 74118
rect 142988 74054 143040 74060
rect 143092 73982 143120 79648
rect 143170 79656 143226 79665
rect 143264 79630 143316 79636
rect 143170 79591 143226 79600
rect 143184 76974 143212 79591
rect 143172 76968 143224 76974
rect 143172 76910 143224 76916
rect 143276 75993 143304 79630
rect 143262 75984 143318 75993
rect 143262 75919 143318 75928
rect 143368 75857 143396 79766
rect 143630 79727 143686 79736
rect 143782 79744 143810 80036
rect 143874 79937 143902 80036
rect 143860 79928 143916 79937
rect 143860 79863 143916 79872
rect 143966 79830 143994 80036
rect 143954 79824 144006 79830
rect 143954 79766 144006 79772
rect 143448 79688 143500 79694
rect 143448 79630 143500 79636
rect 143460 77586 143488 79630
rect 143540 79620 143592 79626
rect 143644 79608 143672 79727
rect 143782 79716 143856 79744
rect 143828 79676 143856 79716
rect 143908 79688 143960 79694
rect 143828 79648 143908 79676
rect 144058 79676 144086 80036
rect 144150 79778 144178 80036
rect 144242 79966 144270 80036
rect 144230 79960 144282 79966
rect 144230 79902 144282 79908
rect 144334 79778 144362 80036
rect 144426 79898 144454 80036
rect 144518 79966 144546 80036
rect 144610 79966 144638 80036
rect 144506 79960 144558 79966
rect 144506 79902 144558 79908
rect 144598 79960 144650 79966
rect 144598 79902 144650 79908
rect 144414 79892 144466 79898
rect 144414 79834 144466 79840
rect 144150 79750 144224 79778
rect 144334 79750 144408 79778
rect 143908 79630 143960 79636
rect 144012 79648 144086 79676
rect 143644 79580 143764 79608
rect 143540 79562 143592 79568
rect 143448 77580 143500 77586
rect 143448 77522 143500 77528
rect 143354 75848 143410 75857
rect 143354 75783 143410 75792
rect 143080 73976 143132 73982
rect 143552 73953 143580 79562
rect 143632 79484 143684 79490
rect 143632 79426 143684 79432
rect 143644 76226 143672 79426
rect 143632 76220 143684 76226
rect 143632 76162 143684 76168
rect 143736 76090 143764 79580
rect 143816 79484 143868 79490
rect 143816 79426 143868 79432
rect 143724 76084 143776 76090
rect 143724 76026 143776 76032
rect 143632 75948 143684 75954
rect 143632 75890 143684 75896
rect 143080 73918 143132 73924
rect 143538 73944 143594 73953
rect 143538 73879 143594 73888
rect 143540 73840 143592 73846
rect 143540 73782 143592 73788
rect 142988 73228 143040 73234
rect 142988 73170 143040 73176
rect 142804 70372 142856 70378
rect 142804 70314 142856 70320
rect 142712 68604 142764 68610
rect 142712 68546 142764 68552
rect 142620 65816 142672 65822
rect 142620 65758 142672 65764
rect 142620 45008 142672 45014
rect 142620 44950 142672 44956
rect 142528 26036 142580 26042
rect 142528 25978 142580 25984
rect 142436 24540 142488 24546
rect 142436 24482 142488 24488
rect 142252 7948 142304 7954
rect 142252 7890 142304 7896
rect 142632 6914 142660 44950
rect 142448 6886 142660 6914
rect 142160 5160 142212 5166
rect 142160 5102 142212 5108
rect 141516 3528 141568 3534
rect 141516 3470 141568 3476
rect 138848 3324 138900 3330
rect 138848 3266 138900 3272
rect 137652 3120 137704 3126
rect 137652 3062 137704 3068
rect 137664 480 137692 3062
rect 138860 480 138888 3266
rect 140044 3188 140096 3194
rect 140044 3130 140096 3136
rect 140056 480 140084 3130
rect 141240 3052 141292 3058
rect 141240 2994 141292 3000
rect 141252 480 141280 2994
rect 142448 480 142476 6886
rect 142816 3466 142844 70314
rect 143000 3874 143028 73170
rect 143552 7886 143580 73782
rect 143644 12034 143672 75890
rect 143724 75880 143776 75886
rect 143724 75822 143776 75828
rect 143736 14822 143764 75822
rect 143828 29918 143856 79426
rect 143908 79348 143960 79354
rect 143908 79290 143960 79296
rect 143920 29986 143948 79290
rect 144012 75954 144040 79648
rect 144092 79552 144144 79558
rect 144092 79494 144144 79500
rect 144000 75948 144052 75954
rect 144000 75890 144052 75896
rect 144000 75812 144052 75818
rect 144000 75754 144052 75760
rect 144012 31482 144040 75754
rect 144104 33862 144132 79494
rect 144196 64462 144224 79750
rect 144276 79620 144328 79626
rect 144276 79562 144328 79568
rect 144288 76906 144316 79562
rect 144380 79472 144408 79750
rect 144460 79688 144512 79694
rect 144458 79656 144460 79665
rect 144552 79688 144604 79694
rect 144512 79656 144514 79665
rect 144702 79676 144730 80036
rect 144552 79630 144604 79636
rect 144656 79648 144730 79676
rect 144458 79591 144514 79600
rect 144380 79444 144500 79472
rect 144368 79348 144420 79354
rect 144368 79290 144420 79296
rect 144380 78946 144408 79290
rect 144368 78940 144420 78946
rect 144368 78882 144420 78888
rect 144366 78840 144422 78849
rect 144366 78775 144422 78784
rect 144276 76900 144328 76906
rect 144276 76842 144328 76848
rect 144276 76084 144328 76090
rect 144276 76026 144328 76032
rect 144288 64530 144316 76026
rect 144380 73846 144408 78775
rect 144472 75886 144500 79444
rect 144460 75880 144512 75886
rect 144460 75822 144512 75828
rect 144564 75818 144592 79630
rect 144656 76129 144684 79648
rect 144794 79642 144822 80036
rect 144886 79971 144914 80036
rect 144872 79962 144928 79971
rect 144872 79897 144928 79906
rect 144978 79898 145006 80036
rect 145070 79971 145098 80036
rect 145056 79962 145112 79971
rect 144966 79892 145018 79898
rect 145056 79897 145112 79906
rect 145162 79898 145190 80036
rect 144966 79834 145018 79840
rect 145150 79892 145202 79898
rect 145150 79834 145202 79840
rect 145254 79812 145282 80036
rect 145346 79966 145374 80036
rect 145334 79960 145386 79966
rect 145334 79902 145386 79908
rect 145010 79792 145066 79801
rect 144920 79756 144972 79762
rect 145254 79784 145328 79812
rect 145010 79727 145066 79736
rect 144920 79698 144972 79704
rect 144794 79614 144868 79642
rect 144736 79552 144788 79558
rect 144736 79494 144788 79500
rect 144748 76294 144776 79494
rect 144840 76945 144868 79614
rect 144932 78606 144960 79698
rect 144920 78600 144972 78606
rect 144920 78542 144972 78548
rect 144826 76936 144882 76945
rect 144826 76871 144882 76880
rect 144736 76288 144788 76294
rect 144736 76230 144788 76236
rect 144642 76120 144698 76129
rect 144642 76055 144698 76064
rect 144644 76016 144696 76022
rect 144644 75958 144696 75964
rect 144920 76016 144972 76022
rect 144920 75958 144972 75964
rect 144552 75812 144604 75818
rect 144552 75754 144604 75760
rect 144368 73840 144420 73846
rect 144368 73782 144420 73788
rect 144656 70394 144684 75958
rect 144472 70366 144684 70394
rect 144276 64524 144328 64530
rect 144276 64466 144328 64472
rect 144184 64456 144236 64462
rect 144184 64398 144236 64404
rect 144092 33856 144144 33862
rect 144092 33798 144144 33804
rect 144000 31476 144052 31482
rect 144000 31418 144052 31424
rect 143908 29980 143960 29986
rect 143908 29922 143960 29928
rect 143816 29912 143868 29918
rect 143816 29854 143868 29860
rect 143724 14816 143776 14822
rect 143724 14758 143776 14764
rect 143632 12028 143684 12034
rect 143632 11970 143684 11976
rect 143540 7880 143592 7886
rect 143540 7822 143592 7828
rect 143540 4412 143592 4418
rect 143540 4354 143592 4360
rect 142988 3868 143040 3874
rect 142988 3810 143040 3816
rect 142804 3460 142856 3466
rect 142804 3402 142856 3408
rect 143552 480 143580 4354
rect 144472 3330 144500 70366
rect 144932 9314 144960 75958
rect 145024 74050 145052 79727
rect 145104 79688 145156 79694
rect 145300 79642 145328 79784
rect 145438 79744 145466 80036
rect 145530 79812 145558 80036
rect 145622 79966 145650 80036
rect 145610 79960 145662 79966
rect 145610 79902 145662 79908
rect 145714 79812 145742 80036
rect 145530 79784 145604 79812
rect 145438 79716 145512 79744
rect 145104 79630 145156 79636
rect 145116 77110 145144 79630
rect 145208 79614 145328 79642
rect 145208 78674 145236 79614
rect 145288 79552 145340 79558
rect 145484 79540 145512 79716
rect 145288 79494 145340 79500
rect 145392 79512 145512 79540
rect 145196 78668 145248 78674
rect 145196 78610 145248 78616
rect 145104 77104 145156 77110
rect 145104 77046 145156 77052
rect 145196 76288 145248 76294
rect 145196 76230 145248 76236
rect 145104 76084 145156 76090
rect 145104 76026 145156 76032
rect 145012 74044 145064 74050
rect 145012 73986 145064 73992
rect 145012 73908 145064 73914
rect 145012 73850 145064 73856
rect 145024 20330 145052 73850
rect 145116 20398 145144 76026
rect 145208 29850 145236 76230
rect 145196 29844 145248 29850
rect 145196 29786 145248 29792
rect 145300 29782 145328 79494
rect 145392 76090 145420 79512
rect 145472 79280 145524 79286
rect 145472 79222 145524 79228
rect 145380 76084 145432 76090
rect 145380 76026 145432 76032
rect 145380 75948 145432 75954
rect 145380 75890 145432 75896
rect 145392 35630 145420 75890
rect 145484 74254 145512 79222
rect 145472 74248 145524 74254
rect 145472 74190 145524 74196
rect 145472 74044 145524 74050
rect 145472 73986 145524 73992
rect 145484 65754 145512 73986
rect 145472 65748 145524 65754
rect 145472 65690 145524 65696
rect 145576 65686 145604 79784
rect 145668 79784 145742 79812
rect 145668 75954 145696 79784
rect 145806 79744 145834 80036
rect 145760 79716 145834 79744
rect 145760 76022 145788 79716
rect 145898 79608 145926 80036
rect 145990 79676 146018 80036
rect 146082 79744 146110 80036
rect 146174 79937 146202 80036
rect 146266 79966 146294 80036
rect 146254 79960 146306 79966
rect 146160 79928 146216 79937
rect 146358 79937 146386 80036
rect 146450 79966 146478 80036
rect 146438 79960 146490 79966
rect 146254 79902 146306 79908
rect 146344 79928 146400 79937
rect 146160 79863 146216 79872
rect 146438 79902 146490 79908
rect 146542 79898 146570 80036
rect 146634 79966 146662 80036
rect 146726 79971 146754 80036
rect 146622 79960 146674 79966
rect 146622 79902 146674 79908
rect 146712 79962 146768 79971
rect 146344 79863 146400 79872
rect 146530 79892 146582 79898
rect 146712 79897 146768 79906
rect 146818 79898 146846 80036
rect 146530 79834 146582 79840
rect 146806 79892 146858 79898
rect 146806 79834 146858 79840
rect 146392 79756 146444 79762
rect 146082 79716 146156 79744
rect 145990 79648 146064 79676
rect 145898 79580 145972 79608
rect 145944 76838 145972 79580
rect 145932 76832 145984 76838
rect 145932 76774 145984 76780
rect 145840 76152 145892 76158
rect 145840 76094 145892 76100
rect 145748 76016 145800 76022
rect 145748 75958 145800 75964
rect 145656 75948 145708 75954
rect 145656 75890 145708 75896
rect 145852 74186 145880 76094
rect 145840 74180 145892 74186
rect 145840 74122 145892 74128
rect 146036 73914 146064 79648
rect 146128 75993 146156 79716
rect 146392 79698 146444 79704
rect 146484 79756 146536 79762
rect 146910 79744 146938 80036
rect 147002 79898 147030 80036
rect 147094 79937 147122 80036
rect 147080 79928 147136 79937
rect 146990 79892 147042 79898
rect 147080 79863 147136 79872
rect 146990 79834 147042 79840
rect 146536 79716 146616 79744
rect 146484 79698 146536 79704
rect 146300 79688 146352 79694
rect 146206 79656 146262 79665
rect 146300 79630 146352 79636
rect 146206 79591 146208 79600
rect 146260 79591 146262 79600
rect 146208 79562 146260 79568
rect 146208 79484 146260 79490
rect 146208 79426 146260 79432
rect 146114 75984 146170 75993
rect 146114 75919 146170 75928
rect 146024 73908 146076 73914
rect 146024 73850 146076 73856
rect 146220 73817 146248 79426
rect 146312 78577 146340 79630
rect 146404 79608 146432 79698
rect 146404 79580 146524 79608
rect 146392 79484 146444 79490
rect 146392 79426 146444 79432
rect 146298 78568 146354 78577
rect 146298 78503 146354 78512
rect 146404 78418 146432 79426
rect 146312 78390 146432 78418
rect 146312 74882 146340 78390
rect 146392 78260 146444 78266
rect 146392 78202 146444 78208
rect 146404 75018 146432 78202
rect 146496 75274 146524 79580
rect 146484 75268 146536 75274
rect 146484 75210 146536 75216
rect 146588 75206 146616 79716
rect 146864 79716 146938 79744
rect 146668 79552 146720 79558
rect 146668 79494 146720 79500
rect 146680 78112 146708 79494
rect 146758 78840 146814 78849
rect 146758 78775 146814 78784
rect 146772 78402 146800 78775
rect 146760 78396 146812 78402
rect 146760 78338 146812 78344
rect 146864 78112 146892 79716
rect 147036 79620 147088 79626
rect 147186 79608 147214 80036
rect 147278 79966 147306 80036
rect 147266 79960 147318 79966
rect 147266 79902 147318 79908
rect 147370 79898 147398 80036
rect 147462 79966 147490 80036
rect 147554 79966 147582 80036
rect 147646 79966 147674 80036
rect 147738 79966 147766 80036
rect 147450 79960 147502 79966
rect 147450 79902 147502 79908
rect 147542 79960 147594 79966
rect 147542 79902 147594 79908
rect 147634 79960 147686 79966
rect 147634 79902 147686 79908
rect 147726 79960 147778 79966
rect 147830 79937 147858 80036
rect 147922 79966 147950 80036
rect 148014 79966 148042 80036
rect 148106 79966 148134 80036
rect 147910 79960 147962 79966
rect 147726 79902 147778 79908
rect 147816 79928 147872 79937
rect 147358 79892 147410 79898
rect 147910 79902 147962 79908
rect 148002 79960 148054 79966
rect 148002 79902 148054 79908
rect 148094 79960 148146 79966
rect 148094 79902 148146 79908
rect 147816 79863 147872 79872
rect 147358 79834 147410 79840
rect 148198 79812 148226 80036
rect 148152 79784 148226 79812
rect 147312 79756 147364 79762
rect 147312 79698 147364 79704
rect 147404 79756 147456 79762
rect 147404 79698 147456 79704
rect 147864 79756 147916 79762
rect 147864 79698 147916 79704
rect 147956 79756 148008 79762
rect 147956 79698 148008 79704
rect 148048 79756 148100 79762
rect 148048 79698 148100 79704
rect 147186 79580 147260 79608
rect 147036 79562 147088 79568
rect 146944 79552 146996 79558
rect 146944 79494 146996 79500
rect 146956 78849 146984 79494
rect 146942 78840 146998 78849
rect 146942 78775 146998 78784
rect 147048 78266 147076 79562
rect 147128 79484 147180 79490
rect 147128 79426 147180 79432
rect 147036 78260 147088 78266
rect 147036 78202 147088 78208
rect 146680 78084 146800 78112
rect 146864 78084 147076 78112
rect 146666 78024 146722 78033
rect 146666 77959 146722 77968
rect 146576 75200 146628 75206
rect 146576 75142 146628 75148
rect 146404 74990 146616 75018
rect 146484 74928 146536 74934
rect 146312 74854 146432 74882
rect 146484 74870 146536 74876
rect 146300 74792 146352 74798
rect 146300 74734 146352 74740
rect 146206 73808 146262 73817
rect 146206 73743 146262 73752
rect 145564 65680 145616 65686
rect 145564 65622 145616 65628
rect 145380 35624 145432 35630
rect 145380 35566 145432 35572
rect 145288 29776 145340 29782
rect 145288 29718 145340 29724
rect 145104 20392 145156 20398
rect 145104 20334 145156 20340
rect 145012 20324 145064 20330
rect 145012 20266 145064 20272
rect 144920 9308 144972 9314
rect 144920 9250 144972 9256
rect 146312 9246 146340 74734
rect 146404 20262 146432 74854
rect 146496 25974 146524 74870
rect 146588 27130 146616 74990
rect 146680 28354 146708 77959
rect 146772 75410 146800 78084
rect 146942 78024 146998 78033
rect 146942 77959 146998 77968
rect 146760 75404 146812 75410
rect 146760 75346 146812 75352
rect 146760 75268 146812 75274
rect 146760 75210 146812 75216
rect 146772 31414 146800 75210
rect 146852 75200 146904 75206
rect 146852 75142 146904 75148
rect 146864 33794 146892 75142
rect 146956 35562 146984 77959
rect 147048 63170 147076 78084
rect 147140 74934 147168 79426
rect 147232 75914 147260 79580
rect 147324 78033 147352 79698
rect 147310 78024 147366 78033
rect 147310 77959 147366 77968
rect 147416 77353 147444 79698
rect 147496 79688 147548 79694
rect 147496 79630 147548 79636
rect 147770 79656 147826 79665
rect 147402 77344 147458 77353
rect 147402 77279 147458 77288
rect 147404 77104 147456 77110
rect 147404 77046 147456 77052
rect 147232 75886 147352 75914
rect 147220 75404 147272 75410
rect 147220 75346 147272 75352
rect 147128 74928 147180 74934
rect 147128 74870 147180 74876
rect 147232 70394 147260 75346
rect 147324 74798 147352 75886
rect 147312 74792 147364 74798
rect 147312 74734 147364 74740
rect 147416 74050 147444 77046
rect 147508 76809 147536 79630
rect 147588 79620 147640 79626
rect 147770 79591 147826 79600
rect 147588 79562 147640 79568
rect 147494 76800 147550 76809
rect 147494 76735 147550 76744
rect 147404 74044 147456 74050
rect 147404 73986 147456 73992
rect 147600 72593 147628 79562
rect 147680 79484 147732 79490
rect 147680 79426 147732 79432
rect 147692 77625 147720 79426
rect 147784 78946 147812 79591
rect 147772 78940 147824 78946
rect 147772 78882 147824 78888
rect 147876 77994 147904 79698
rect 147864 77988 147916 77994
rect 147864 77930 147916 77936
rect 147678 77616 147734 77625
rect 147678 77551 147734 77560
rect 147968 76770 147996 79698
rect 147956 76764 148008 76770
rect 147956 76706 148008 76712
rect 147862 75984 147918 75993
rect 147862 75919 147918 75928
rect 147772 75880 147824 75886
rect 147772 75822 147824 75828
rect 147680 74656 147732 74662
rect 147680 74598 147732 74604
rect 147586 72584 147642 72593
rect 147586 72519 147642 72528
rect 147140 70366 147260 70394
rect 147140 67386 147168 70366
rect 147128 67380 147180 67386
rect 147128 67322 147180 67328
rect 147036 63164 147088 63170
rect 147036 63106 147088 63112
rect 147036 44872 147088 44878
rect 147036 44814 147088 44820
rect 146944 35556 146996 35562
rect 146944 35498 146996 35504
rect 146852 33788 146904 33794
rect 146852 33730 146904 33736
rect 146760 31408 146812 31414
rect 146760 31350 146812 31356
rect 146668 28348 146720 28354
rect 146668 28290 146720 28296
rect 146576 27124 146628 27130
rect 146576 27066 146628 27072
rect 146484 25968 146536 25974
rect 146484 25910 146536 25916
rect 146392 20256 146444 20262
rect 146392 20198 146444 20204
rect 147048 16574 147076 44814
rect 147048 16546 147260 16574
rect 146300 9240 146352 9246
rect 146300 9182 146352 9188
rect 145932 4072 145984 4078
rect 145932 4014 145984 4020
rect 144736 3936 144788 3942
rect 144736 3878 144788 3884
rect 144460 3324 144512 3330
rect 144460 3266 144512 3272
rect 144748 480 144776 3878
rect 145944 480 145972 4014
rect 147232 3602 147260 16546
rect 147692 10606 147720 74598
rect 147784 24478 147812 75822
rect 147876 28286 147904 75919
rect 148060 75914 148088 79698
rect 148152 78198 148180 79784
rect 148290 79744 148318 80036
rect 148382 79966 148410 80036
rect 148474 79966 148502 80036
rect 148370 79960 148422 79966
rect 148370 79902 148422 79908
rect 148462 79960 148514 79966
rect 148462 79902 148514 79908
rect 148566 79744 148594 80036
rect 148658 79937 148686 80036
rect 148750 79966 148778 80036
rect 148738 79960 148790 79966
rect 148644 79928 148700 79937
rect 148738 79902 148790 79908
rect 148644 79863 148700 79872
rect 148244 79716 148318 79744
rect 148520 79716 148594 79744
rect 148842 79744 148870 80036
rect 148934 79971 148962 80036
rect 148920 79962 148976 79971
rect 148920 79897 148976 79906
rect 149026 79812 149054 80036
rect 149118 79966 149146 80036
rect 149106 79960 149158 79966
rect 149210 79937 149238 80036
rect 149106 79902 149158 79908
rect 149196 79928 149252 79937
rect 149302 79898 149330 80036
rect 149196 79863 149252 79872
rect 149290 79892 149342 79898
rect 149290 79834 149342 79840
rect 149026 79784 149100 79812
rect 148842 79716 149008 79744
rect 148140 78192 148192 78198
rect 148140 78134 148192 78140
rect 148140 77988 148192 77994
rect 148140 77930 148192 77936
rect 147968 75886 148088 75914
rect 147968 31346 147996 75886
rect 148048 75812 148100 75818
rect 148048 75754 148100 75760
rect 148060 35426 148088 75754
rect 148152 35494 148180 77930
rect 148244 64394 148272 79716
rect 148324 79620 148376 79626
rect 148324 79562 148376 79568
rect 148336 78282 148364 79562
rect 148416 79348 148468 79354
rect 148416 79290 148468 79296
rect 148428 79150 148456 79290
rect 148416 79144 148468 79150
rect 148416 79086 148468 79092
rect 148336 78254 148456 78282
rect 148324 78192 148376 78198
rect 148324 78134 148376 78140
rect 148336 72690 148364 78134
rect 148428 75886 148456 78254
rect 148416 75880 148468 75886
rect 148416 75822 148468 75828
rect 148520 74662 148548 79716
rect 148874 79656 148930 79665
rect 148600 79620 148652 79626
rect 148600 79562 148652 79568
rect 148784 79620 148836 79626
rect 148874 79591 148930 79600
rect 148784 79562 148836 79568
rect 148612 75818 148640 79562
rect 148796 77897 148824 79562
rect 148782 77888 148838 77897
rect 148782 77823 148838 77832
rect 148888 76702 148916 79591
rect 148876 76696 148928 76702
rect 148876 76638 148928 76644
rect 148692 76220 148744 76226
rect 148692 76162 148744 76168
rect 148600 75812 148652 75818
rect 148600 75754 148652 75760
rect 148508 74656 148560 74662
rect 148508 74598 148560 74604
rect 148324 72684 148376 72690
rect 148324 72626 148376 72632
rect 148704 70394 148732 76162
rect 148980 75993 149008 79716
rect 149072 78441 149100 79784
rect 149150 79792 149206 79801
rect 149394 79778 149422 80036
rect 149486 79966 149514 80036
rect 149474 79960 149526 79966
rect 149474 79902 149526 79908
rect 149578 79778 149606 80036
rect 149670 79966 149698 80036
rect 149762 79966 149790 80036
rect 149658 79960 149710 79966
rect 149658 79902 149710 79908
rect 149750 79960 149802 79966
rect 149750 79902 149802 79908
rect 149150 79727 149206 79736
rect 149256 79750 149422 79778
rect 149532 79750 149606 79778
rect 149704 79824 149756 79830
rect 149704 79766 149756 79772
rect 149058 78432 149114 78441
rect 149058 78367 149114 78376
rect 148966 75984 149022 75993
rect 148966 75919 149022 75928
rect 148704 70366 148824 70394
rect 148796 64874 148824 70366
rect 148704 64846 148824 64874
rect 148232 64388 148284 64394
rect 148232 64330 148284 64336
rect 148140 35488 148192 35494
rect 148140 35430 148192 35436
rect 148048 35420 148100 35426
rect 148048 35362 148100 35368
rect 147956 31340 148008 31346
rect 147956 31282 148008 31288
rect 148704 28558 148732 64846
rect 148692 28552 148744 28558
rect 148692 28494 148744 28500
rect 147864 28280 147916 28286
rect 147864 28222 147916 28228
rect 147772 24472 147824 24478
rect 147772 24414 147824 24420
rect 149164 23390 149192 79727
rect 149256 78062 149284 79750
rect 149336 79688 149388 79694
rect 149336 79630 149388 79636
rect 149244 78056 149296 78062
rect 149244 77998 149296 78004
rect 149348 75914 149376 79630
rect 149428 79620 149480 79626
rect 149428 79562 149480 79568
rect 149256 75886 149376 75914
rect 149256 25906 149284 75886
rect 149336 75268 149388 75274
rect 149336 75210 149388 75216
rect 149348 27062 149376 75210
rect 149440 35358 149468 79562
rect 149428 35352 149480 35358
rect 149428 35294 149480 35300
rect 149532 35290 149560 79750
rect 149612 79688 149664 79694
rect 149612 79630 149664 79636
rect 149624 63102 149652 79630
rect 149716 75274 149744 79766
rect 149854 79744 149882 80036
rect 149946 79898 149974 80036
rect 150038 79966 150066 80036
rect 150026 79960 150078 79966
rect 150026 79902 150078 79908
rect 149934 79892 149986 79898
rect 149934 79834 149986 79840
rect 150130 79801 150158 80036
rect 150116 79792 150172 79801
rect 149854 79716 149928 79744
rect 150116 79727 150172 79736
rect 150222 79744 150250 80036
rect 150314 79971 150342 80036
rect 150300 79962 150356 79971
rect 150300 79897 150356 79906
rect 150406 79898 150434 80036
rect 150394 79892 150446 79898
rect 150394 79834 150446 79840
rect 150498 79744 150526 80036
rect 150222 79716 150296 79744
rect 149796 78056 149848 78062
rect 149796 77998 149848 78004
rect 149704 75268 149756 75274
rect 149704 75210 149756 75216
rect 149808 70394 149836 77998
rect 149900 72622 149928 79716
rect 149980 79620 150032 79626
rect 149980 79562 150032 79568
rect 149992 78713 150020 79562
rect 150072 79552 150124 79558
rect 150072 79494 150124 79500
rect 149978 78704 150034 78713
rect 149978 78639 150034 78648
rect 150084 77994 150112 79494
rect 150268 78577 150296 79716
rect 150452 79716 150526 79744
rect 150590 79744 150618 80036
rect 150682 79812 150710 80036
rect 150774 79937 150802 80036
rect 150866 79966 150894 80036
rect 150854 79960 150906 79966
rect 150760 79928 150816 79937
rect 150854 79902 150906 79908
rect 150760 79863 150816 79872
rect 150682 79784 150848 79812
rect 150590 79716 150664 79744
rect 150348 79688 150400 79694
rect 150348 79630 150400 79636
rect 150254 78568 150310 78577
rect 150254 78503 150310 78512
rect 150164 78124 150216 78130
rect 150164 78066 150216 78072
rect 150072 77988 150124 77994
rect 150072 77930 150124 77936
rect 150176 77110 150204 78066
rect 150164 77104 150216 77110
rect 150164 77046 150216 77052
rect 149888 72616 149940 72622
rect 149888 72558 149940 72564
rect 149716 70366 149836 70394
rect 149716 67318 149744 70366
rect 149704 67312 149756 67318
rect 149704 67254 149756 67260
rect 149612 63096 149664 63102
rect 149612 63038 149664 63044
rect 149520 35284 149572 35290
rect 149520 35226 149572 35232
rect 149336 27056 149388 27062
rect 149336 26998 149388 27004
rect 149244 25900 149296 25906
rect 149244 25842 149296 25848
rect 149152 23384 149204 23390
rect 149152 23326 149204 23332
rect 150360 11966 150388 79630
rect 150452 74390 150480 79716
rect 150532 79620 150584 79626
rect 150532 79562 150584 79568
rect 150544 76158 150572 79562
rect 150532 76152 150584 76158
rect 150532 76094 150584 76100
rect 150440 74384 150492 74390
rect 150440 74326 150492 74332
rect 150532 73772 150584 73778
rect 150532 73714 150584 73720
rect 150348 11960 150400 11966
rect 150348 11902 150400 11908
rect 147680 10600 147732 10606
rect 147680 10542 147732 10548
rect 148324 5092 148376 5098
rect 148324 5034 148376 5040
rect 147128 3596 147180 3602
rect 147128 3538 147180 3544
rect 147220 3596 147272 3602
rect 147220 3538 147272 3544
rect 147140 480 147168 3538
rect 148336 480 148364 5034
rect 150544 4010 150572 73714
rect 150636 5114 150664 79716
rect 150716 79688 150768 79694
rect 150716 79630 150768 79636
rect 150728 5522 150756 79630
rect 150820 6798 150848 79784
rect 150958 79744 150986 80036
rect 151050 79966 151078 80036
rect 151038 79960 151090 79966
rect 151038 79902 151090 79908
rect 151142 79812 151170 80036
rect 151234 79898 151262 80036
rect 151222 79892 151274 79898
rect 151222 79834 151274 79840
rect 151096 79784 151170 79812
rect 150958 79716 151032 79744
rect 150900 76628 150952 76634
rect 150900 76570 150952 76576
rect 150808 6792 150860 6798
rect 150808 6734 150860 6740
rect 150912 6662 150940 76570
rect 151004 6730 151032 79716
rect 151096 76634 151124 79784
rect 151326 79744 151354 80036
rect 151418 79937 151446 80036
rect 151404 79928 151460 79937
rect 151510 79898 151538 80036
rect 151602 79966 151630 80036
rect 151590 79960 151642 79966
rect 151590 79902 151642 79908
rect 151694 79898 151722 80036
rect 151404 79863 151460 79872
rect 151498 79892 151550 79898
rect 151498 79834 151550 79840
rect 151682 79892 151734 79898
rect 151682 79834 151734 79840
rect 151786 79801 151814 80036
rect 151280 79716 151354 79744
rect 151772 79792 151828 79801
rect 151772 79727 151828 79736
rect 151878 79744 151906 80036
rect 151970 79937 151998 80036
rect 151956 79928 152012 79937
rect 152062 79898 152090 80036
rect 151956 79863 152012 79872
rect 152050 79892 152102 79898
rect 152050 79834 152102 79840
rect 152002 79792 152058 79801
rect 151878 79716 151952 79744
rect 152002 79727 152058 79736
rect 152154 79744 152182 80036
rect 152246 79966 152274 80036
rect 152234 79960 152286 79966
rect 152234 79902 152286 79908
rect 152338 79812 152366 80036
rect 152292 79784 152366 79812
rect 151176 79688 151228 79694
rect 151176 79630 151228 79636
rect 151084 76628 151136 76634
rect 151084 76570 151136 76576
rect 151188 70394 151216 79630
rect 151280 73778 151308 79716
rect 151360 79620 151412 79626
rect 151360 79562 151412 79568
rect 151728 79620 151780 79626
rect 151728 79562 151780 79568
rect 151820 79620 151872 79626
rect 151820 79562 151872 79568
rect 151268 73772 151320 73778
rect 151268 73714 151320 73720
rect 151096 70366 151216 70394
rect 151372 70394 151400 79562
rect 151636 79552 151688 79558
rect 151636 79494 151688 79500
rect 151648 76673 151676 79494
rect 151634 76664 151690 76673
rect 151634 76599 151690 76608
rect 151740 76537 151768 79562
rect 151726 76528 151782 76537
rect 151726 76463 151782 76472
rect 151372 70366 151584 70394
rect 150992 6724 151044 6730
rect 150992 6666 151044 6672
rect 150900 6656 150952 6662
rect 150900 6598 150952 6604
rect 151096 6594 151124 70366
rect 151084 6588 151136 6594
rect 151084 6530 151136 6536
rect 150728 5494 150940 5522
rect 150636 5086 150848 5114
rect 150624 4956 150676 4962
rect 150624 4898 150676 4904
rect 150532 4004 150584 4010
rect 150532 3946 150584 3952
rect 149520 3800 149572 3806
rect 149520 3742 149572 3748
rect 149532 480 149560 3742
rect 150636 480 150664 4898
rect 150820 3398 150848 5086
rect 150912 4078 150940 5494
rect 151556 4146 151584 70366
rect 151832 9178 151860 79562
rect 151924 76566 151952 79716
rect 151912 76560 151964 76566
rect 151912 76502 151964 76508
rect 151912 76356 151964 76362
rect 151912 76298 151964 76304
rect 151924 13462 151952 76298
rect 152016 76226 152044 79727
rect 152154 79716 152228 79744
rect 152200 77042 152228 79716
rect 152188 77036 152240 77042
rect 152188 76978 152240 76984
rect 152292 76786 152320 79784
rect 152430 79744 152458 80036
rect 152108 76758 152320 76786
rect 152384 79716 152458 79744
rect 152522 79744 152550 80036
rect 152614 79937 152642 80036
rect 152706 79966 152734 80036
rect 152694 79960 152746 79966
rect 152600 79928 152656 79937
rect 152798 79937 152826 80036
rect 152890 79966 152918 80036
rect 152982 79966 153010 80036
rect 153074 79966 153102 80036
rect 153166 79971 153194 80036
rect 152878 79960 152930 79966
rect 152694 79902 152746 79908
rect 152784 79928 152840 79937
rect 152600 79863 152656 79872
rect 152878 79902 152930 79908
rect 152970 79960 153022 79966
rect 152970 79902 153022 79908
rect 153062 79960 153114 79966
rect 153062 79902 153114 79908
rect 153152 79962 153208 79971
rect 153258 79966 153286 80036
rect 153152 79897 153208 79906
rect 153246 79960 153298 79966
rect 153246 79902 153298 79908
rect 152784 79863 152840 79872
rect 152648 79824 152700 79830
rect 152648 79766 152700 79772
rect 153016 79824 153068 79830
rect 153016 79766 153068 79772
rect 153106 79792 153162 79801
rect 152522 79716 152596 79744
rect 152004 76220 152056 76226
rect 152004 76162 152056 76168
rect 152004 73908 152056 73914
rect 152004 73850 152056 73856
rect 151912 13456 151964 13462
rect 151912 13398 151964 13404
rect 152016 13394 152044 73850
rect 152108 21690 152136 76758
rect 152384 76650 152412 79716
rect 152462 79656 152518 79665
rect 152462 79591 152518 79600
rect 152476 77926 152504 79591
rect 152464 77920 152516 77926
rect 152464 77862 152516 77868
rect 152464 77036 152516 77042
rect 152464 76978 152516 76984
rect 152188 76628 152240 76634
rect 152188 76570 152240 76576
rect 152292 76622 152412 76650
rect 152200 25838 152228 76570
rect 152292 76362 152320 76622
rect 152372 76560 152424 76566
rect 152372 76502 152424 76508
rect 152280 76356 152332 76362
rect 152280 76298 152332 76304
rect 152280 76220 152332 76226
rect 152280 76162 152332 76168
rect 152292 26994 152320 76162
rect 152384 64326 152412 76502
rect 152476 67182 152504 76978
rect 152568 76634 152596 79716
rect 152556 76628 152608 76634
rect 152556 76570 152608 76576
rect 152660 73914 152688 79766
rect 152740 79756 152792 79762
rect 152740 79698 152792 79704
rect 152752 78577 152780 79698
rect 152832 79688 152884 79694
rect 152832 79630 152884 79636
rect 152738 78568 152794 78577
rect 152738 78503 152794 78512
rect 152844 76537 152872 79630
rect 152924 79620 152976 79626
rect 152924 79562 152976 79568
rect 152830 76528 152886 76537
rect 152830 76463 152886 76472
rect 152648 73908 152700 73914
rect 152648 73850 152700 73856
rect 152936 73154 152964 79562
rect 153028 76673 153056 79766
rect 153106 79727 153162 79736
rect 153120 78198 153148 79727
rect 153350 79676 153378 80036
rect 153198 79656 153254 79665
rect 153198 79591 153254 79600
rect 153304 79648 153378 79676
rect 153442 79676 153470 80036
rect 153534 79744 153562 80036
rect 153626 79898 153654 80036
rect 153718 79937 153746 80036
rect 153704 79928 153760 79937
rect 153614 79892 153666 79898
rect 153704 79863 153760 79872
rect 153614 79834 153666 79840
rect 153810 79744 153838 80036
rect 153534 79716 153700 79744
rect 153442 79648 153516 79676
rect 153108 78192 153160 78198
rect 153108 78134 153160 78140
rect 153212 77330 153240 79591
rect 153120 77302 153240 77330
rect 153014 76664 153070 76673
rect 153014 76599 153070 76608
rect 153120 73914 153148 77302
rect 153200 77240 153252 77246
rect 153200 77182 153252 77188
rect 153108 73908 153160 73914
rect 153108 73850 153160 73856
rect 152752 73126 152964 73154
rect 152752 72554 152780 73126
rect 152740 72548 152792 72554
rect 152740 72490 152792 72496
rect 153212 72486 153240 77182
rect 153304 76634 153332 79648
rect 153384 79484 153436 79490
rect 153384 79426 153436 79432
rect 153396 77081 153424 79426
rect 153488 77246 153516 79648
rect 153568 79620 153620 79626
rect 153568 79562 153620 79568
rect 153580 77314 153608 79562
rect 153568 77308 153620 77314
rect 153568 77250 153620 77256
rect 153476 77240 153528 77246
rect 153476 77182 153528 77188
rect 153382 77072 153438 77081
rect 153382 77007 153438 77016
rect 153476 77036 153528 77042
rect 153476 76978 153528 76984
rect 153382 76664 153438 76673
rect 153292 76628 153344 76634
rect 153382 76599 153438 76608
rect 153292 76570 153344 76576
rect 153292 74452 153344 74458
rect 153292 74394 153344 74400
rect 153200 72480 153252 72486
rect 153200 72422 153252 72428
rect 152556 71052 152608 71058
rect 152556 70994 152608 71000
rect 152464 67176 152516 67182
rect 152464 67118 152516 67124
rect 152372 64320 152424 64326
rect 152372 64262 152424 64268
rect 152280 26988 152332 26994
rect 152280 26930 152332 26936
rect 152188 25832 152240 25838
rect 152188 25774 152240 25780
rect 152096 21684 152148 21690
rect 152096 21626 152148 21632
rect 152004 13388 152056 13394
rect 152004 13330 152056 13336
rect 151820 9172 151872 9178
rect 151820 9114 151872 9120
rect 151544 4140 151596 4146
rect 151544 4082 151596 4088
rect 150900 4072 150952 4078
rect 150900 4014 150952 4020
rect 151820 3868 151872 3874
rect 151820 3810 151872 3816
rect 150808 3392 150860 3398
rect 150808 3334 150860 3340
rect 151832 480 151860 3810
rect 152568 3806 152596 70994
rect 153304 10538 153332 74394
rect 153396 13326 153424 76599
rect 153488 23254 153516 76978
rect 153568 76628 153620 76634
rect 153568 76570 153620 76576
rect 153580 31210 153608 76570
rect 153672 65618 153700 79716
rect 153764 79716 153838 79744
rect 153764 68474 153792 79716
rect 153902 79676 153930 80036
rect 153994 79744 154022 80036
rect 154086 79937 154114 80036
rect 154072 79928 154128 79937
rect 154072 79863 154128 79872
rect 154178 79801 154206 80036
rect 154164 79792 154220 79801
rect 153994 79716 154068 79744
rect 154164 79727 154220 79736
rect 153856 79648 153930 79676
rect 153856 74458 153884 79648
rect 154040 76650 154068 79716
rect 154270 79676 154298 80036
rect 154362 79744 154390 80036
rect 154454 79937 154482 80036
rect 154440 79928 154496 79937
rect 154440 79863 154496 79872
rect 154546 79812 154574 80036
rect 154500 79784 154574 79812
rect 154362 79716 154436 79744
rect 154270 79648 154344 79676
rect 154120 79552 154172 79558
rect 154120 79494 154172 79500
rect 154132 77042 154160 79494
rect 154316 78334 154344 79648
rect 154304 78328 154356 78334
rect 154304 78270 154356 78276
rect 154120 77036 154172 77042
rect 154120 76978 154172 76984
rect 154408 76673 154436 79716
rect 154394 76664 154450 76673
rect 154040 76622 154344 76650
rect 154210 76392 154266 76401
rect 154210 76327 154266 76336
rect 153844 74452 153896 74458
rect 153844 74394 153896 74400
rect 153752 68468 153804 68474
rect 153752 68410 153804 68416
rect 153660 65612 153712 65618
rect 153660 65554 153712 65560
rect 154224 64874 154252 76327
rect 154316 70394 154344 76622
rect 154394 76599 154450 76608
rect 154500 76537 154528 79784
rect 154638 79744 154666 80036
rect 154730 79937 154758 80036
rect 154822 79966 154850 80036
rect 154810 79960 154862 79966
rect 154716 79928 154772 79937
rect 154810 79902 154862 79908
rect 154716 79863 154772 79872
rect 154914 79812 154942 80036
rect 154776 79784 154942 79812
rect 154638 79716 154712 79744
rect 154578 79656 154634 79665
rect 154578 79591 154634 79600
rect 154486 76528 154542 76537
rect 154486 76463 154542 76472
rect 154592 76294 154620 79591
rect 154580 76288 154632 76294
rect 154580 76230 154632 76236
rect 154684 76226 154712 79716
rect 154776 76634 154804 79784
rect 155006 79744 155034 80036
rect 154868 79716 155034 79744
rect 154764 76628 154816 76634
rect 154764 76570 154816 76576
rect 154764 76356 154816 76362
rect 154764 76298 154816 76304
rect 154672 76220 154724 76226
rect 154672 76162 154724 76168
rect 154580 74588 154632 74594
rect 154580 74530 154632 74536
rect 154316 70366 154528 70394
rect 154132 64846 154252 64874
rect 154132 31278 154160 64846
rect 154120 31272 154172 31278
rect 154120 31214 154172 31220
rect 153568 31204 153620 31210
rect 153568 31146 153620 31152
rect 153476 23248 153528 23254
rect 153476 23190 153528 23196
rect 153384 13320 153436 13326
rect 153384 13262 153436 13268
rect 153292 10532 153344 10538
rect 153292 10474 153344 10480
rect 154500 5098 154528 70366
rect 154592 14618 154620 74530
rect 154776 73386 154804 76298
rect 154684 73358 154804 73386
rect 154684 14754 154712 73358
rect 154764 73296 154816 73302
rect 154764 73238 154816 73244
rect 154672 14748 154724 14754
rect 154672 14690 154724 14696
rect 154776 14686 154804 73238
rect 154868 16182 154896 79716
rect 155098 79676 155126 80036
rect 154960 79648 155126 79676
rect 154960 23186 154988 79648
rect 155190 79608 155218 80036
rect 155282 79744 155310 80036
rect 155374 79898 155402 80036
rect 155466 79937 155494 80036
rect 155452 79928 155508 79937
rect 155362 79892 155414 79898
rect 155452 79863 155508 79872
rect 155362 79834 155414 79840
rect 155406 79792 155462 79801
rect 155282 79716 155356 79744
rect 155558 79744 155586 80036
rect 155650 79778 155678 80036
rect 155742 79937 155770 80036
rect 155728 79928 155784 79937
rect 155834 79898 155862 80036
rect 155728 79863 155784 79872
rect 155822 79892 155874 79898
rect 155822 79834 155874 79840
rect 155926 79778 155954 80036
rect 156018 79898 156046 80036
rect 156110 79937 156138 80036
rect 156202 79966 156230 80036
rect 156190 79960 156242 79966
rect 156096 79928 156152 79937
rect 156006 79892 156058 79898
rect 156190 79902 156242 79908
rect 156294 79898 156322 80036
rect 156386 79966 156414 80036
rect 156478 79966 156506 80036
rect 156374 79960 156426 79966
rect 156374 79902 156426 79908
rect 156466 79960 156518 79966
rect 156570 79937 156598 80036
rect 156466 79902 156518 79908
rect 156556 79928 156612 79937
rect 156096 79863 156152 79872
rect 156282 79892 156334 79898
rect 156006 79834 156058 79840
rect 156556 79863 156612 79872
rect 156282 79834 156334 79840
rect 156662 79830 156690 80036
rect 156754 79898 156782 80036
rect 156846 79966 156874 80036
rect 156834 79960 156886 79966
rect 156834 79902 156886 79908
rect 156742 79892 156794 79898
rect 156742 79834 156794 79840
rect 156938 79830 156966 80036
rect 155650 79750 155724 79778
rect 155406 79727 155462 79736
rect 155144 79580 155218 79608
rect 155040 79348 155092 79354
rect 155040 79290 155092 79296
rect 155052 78305 155080 79290
rect 155038 78296 155094 78305
rect 155038 78231 155094 78240
rect 155038 78160 155094 78169
rect 155038 78095 155094 78104
rect 155052 24410 155080 78095
rect 155144 76362 155172 79580
rect 155224 79484 155276 79490
rect 155224 79426 155276 79432
rect 155236 79218 155264 79426
rect 155224 79212 155276 79218
rect 155224 79154 155276 79160
rect 155224 78872 155276 78878
rect 155224 78814 155276 78820
rect 155236 78470 155264 78814
rect 155224 78464 155276 78470
rect 155224 78406 155276 78412
rect 155224 77512 155276 77518
rect 155224 77454 155276 77460
rect 155236 77382 155264 77454
rect 155224 77376 155276 77382
rect 155224 77318 155276 77324
rect 155224 76628 155276 76634
rect 155224 76570 155276 76576
rect 155132 76356 155184 76362
rect 155132 76298 155184 76304
rect 155132 76220 155184 76226
rect 155132 76162 155184 76168
rect 155144 63034 155172 76162
rect 155236 65550 155264 76570
rect 155328 70038 155356 79716
rect 155420 73302 155448 79727
rect 155512 79716 155586 79744
rect 155512 74594 155540 79716
rect 155696 79642 155724 79750
rect 155776 79756 155828 79762
rect 155776 79698 155828 79704
rect 155880 79750 155954 79778
rect 156374 79824 156426 79830
rect 156650 79824 156702 79830
rect 156510 79792 156566 79801
rect 156426 79772 156510 79778
rect 156374 79766 156510 79772
rect 156386 79750 156510 79766
rect 155604 79614 155724 79642
rect 155604 76673 155632 79614
rect 155590 76664 155646 76673
rect 155590 76599 155646 76608
rect 155788 75886 155816 79698
rect 155880 79608 155908 79750
rect 156650 79766 156702 79772
rect 156926 79824 156978 79830
rect 157030 79812 157058 80036
rect 157122 79937 157150 80036
rect 157108 79928 157164 79937
rect 157108 79863 157164 79872
rect 157030 79784 157104 79812
rect 157214 79801 157242 80036
rect 157306 79830 157334 80036
rect 157398 79898 157426 80036
rect 157386 79892 157438 79898
rect 157386 79834 157438 79840
rect 157490 79830 157518 80036
rect 157294 79824 157346 79830
rect 156926 79766 156978 79772
rect 156510 79727 156566 79736
rect 156052 79688 156104 79694
rect 156052 79630 156104 79636
rect 156144 79688 156196 79694
rect 156144 79630 156196 79636
rect 156236 79688 156288 79694
rect 156604 79688 156656 79694
rect 156236 79630 156288 79636
rect 156418 79656 156474 79665
rect 155880 79580 156000 79608
rect 155868 79484 155920 79490
rect 155868 79426 155920 79432
rect 155776 75880 155828 75886
rect 155776 75822 155828 75828
rect 155880 74866 155908 79426
rect 155972 77625 156000 79580
rect 155958 77616 156014 77625
rect 155958 77551 156014 77560
rect 155868 74860 155920 74866
rect 155868 74802 155920 74808
rect 155500 74588 155552 74594
rect 155500 74530 155552 74536
rect 155960 73500 156012 73506
rect 155960 73442 156012 73448
rect 155408 73296 155460 73302
rect 155408 73238 155460 73244
rect 155316 70032 155368 70038
rect 155316 69974 155368 69980
rect 155224 65544 155276 65550
rect 155224 65486 155276 65492
rect 155132 63028 155184 63034
rect 155132 62970 155184 62976
rect 155040 24404 155092 24410
rect 155040 24346 155092 24352
rect 154948 23180 155000 23186
rect 154948 23122 155000 23128
rect 154856 16176 154908 16182
rect 154856 16118 154908 16124
rect 154764 14680 154816 14686
rect 154764 14622 154816 14628
rect 154580 14612 154632 14618
rect 154580 14554 154632 14560
rect 155972 7818 156000 73442
rect 156064 10470 156092 79630
rect 156156 77246 156184 79630
rect 156144 77240 156196 77246
rect 156144 77182 156196 77188
rect 156144 76628 156196 76634
rect 156144 76570 156196 76576
rect 156052 10464 156104 10470
rect 156052 10406 156104 10412
rect 156156 10402 156184 76570
rect 156248 16114 156276 79630
rect 156604 79630 156656 79636
rect 156418 79591 156474 79600
rect 156512 79620 156564 79626
rect 156328 79552 156380 79558
rect 156328 79494 156380 79500
rect 156340 77314 156368 79494
rect 156328 77308 156380 77314
rect 156328 77250 156380 77256
rect 156432 76786 156460 79591
rect 156512 79562 156564 79568
rect 156340 76758 156460 76786
rect 156236 16108 156288 16114
rect 156236 16050 156288 16056
rect 156340 16046 156368 76758
rect 156418 76664 156474 76673
rect 156418 76599 156474 76608
rect 156432 32774 156460 76599
rect 156524 73506 156552 79562
rect 156616 76634 156644 79630
rect 156972 79552 157024 79558
rect 156972 79494 157024 79500
rect 156696 79416 156748 79422
rect 156696 79358 156748 79364
rect 156708 79218 156736 79358
rect 156696 79212 156748 79218
rect 156696 79154 156748 79160
rect 156984 77897 157012 79494
rect 157076 78169 157104 79784
rect 157200 79792 157256 79801
rect 157294 79766 157346 79772
rect 157478 79824 157530 79830
rect 157478 79766 157530 79772
rect 157200 79727 157256 79736
rect 157156 79688 157208 79694
rect 157156 79630 157208 79636
rect 157248 79688 157300 79694
rect 157248 79630 157300 79636
rect 157340 79688 157392 79694
rect 157582 79676 157610 80036
rect 157674 79744 157702 80036
rect 157766 79937 157794 80036
rect 157752 79928 157808 79937
rect 157858 79898 157886 80036
rect 157752 79863 157808 79872
rect 157846 79892 157898 79898
rect 157846 79834 157898 79840
rect 157950 79744 157978 80036
rect 157674 79716 157748 79744
rect 157340 79630 157392 79636
rect 157536 79648 157610 79676
rect 157062 78160 157118 78169
rect 157062 78095 157118 78104
rect 157064 77988 157116 77994
rect 157064 77930 157116 77936
rect 156970 77888 157026 77897
rect 156970 77823 157026 77832
rect 156972 77240 157024 77246
rect 156972 77182 157024 77188
rect 156604 76628 156656 76634
rect 156604 76570 156656 76576
rect 156696 76628 156748 76634
rect 156696 76570 156748 76576
rect 156512 73500 156564 73506
rect 156512 73442 156564 73448
rect 156708 70394 156736 76570
rect 156984 76378 157012 77182
rect 156524 70366 156736 70394
rect 156800 76350 157012 76378
rect 156524 58682 156552 70366
rect 156800 69970 156828 76350
rect 156972 75880 157024 75886
rect 156972 75822 157024 75828
rect 156880 74384 156932 74390
rect 156880 74326 156932 74332
rect 156788 69964 156840 69970
rect 156788 69906 156840 69912
rect 156892 68542 156920 74326
rect 156880 68536 156932 68542
rect 156880 68478 156932 68484
rect 156512 58676 156564 58682
rect 156512 58618 156564 58624
rect 156420 32768 156472 32774
rect 156420 32710 156472 32716
rect 156984 31142 157012 75822
rect 157076 73154 157104 77930
rect 157168 76634 157196 79630
rect 157260 76673 157288 79630
rect 157246 76664 157302 76673
rect 157156 76628 157208 76634
rect 157246 76599 157302 76608
rect 157156 76570 157208 76576
rect 157352 75342 157380 79630
rect 157432 79620 157484 79626
rect 157432 79562 157484 79568
rect 157444 77042 157472 79562
rect 157536 77654 157564 79648
rect 157616 79552 157668 79558
rect 157616 79494 157668 79500
rect 157524 77648 157576 77654
rect 157524 77590 157576 77596
rect 157432 77036 157484 77042
rect 157432 76978 157484 76984
rect 157628 76786 157656 79494
rect 157444 76758 157656 76786
rect 157340 75336 157392 75342
rect 157340 75278 157392 75284
rect 157076 73126 157380 73154
rect 157352 71058 157380 73126
rect 157340 71052 157392 71058
rect 157340 70994 157392 71000
rect 156972 31136 157024 31142
rect 156972 31078 157024 31084
rect 156328 16040 156380 16046
rect 156328 15982 156380 15988
rect 157444 11830 157472 76758
rect 157522 76664 157578 76673
rect 157720 76634 157748 79716
rect 157812 79716 157978 79744
rect 158042 79744 158070 80036
rect 158134 79898 158162 80036
rect 158122 79892 158174 79898
rect 158122 79834 158174 79840
rect 158226 79744 158254 80036
rect 158318 79801 158346 80036
rect 158042 79716 158116 79744
rect 157522 76599 157578 76608
rect 157708 76628 157760 76634
rect 157536 11898 157564 76599
rect 157708 76570 157760 76576
rect 157616 75948 157668 75954
rect 157616 75890 157668 75896
rect 157628 13258 157656 75890
rect 157708 73976 157760 73982
rect 157708 73918 157760 73924
rect 157720 17542 157748 73918
rect 157812 17610 157840 79716
rect 157984 79620 158036 79626
rect 157984 79562 158036 79568
rect 157892 79484 157944 79490
rect 157892 79426 157944 79432
rect 157904 76786 157932 79426
rect 157996 79218 158024 79562
rect 157984 79212 158036 79218
rect 157984 79154 158036 79160
rect 157904 76758 158024 76786
rect 157892 76628 157944 76634
rect 157892 76570 157944 76576
rect 157904 61470 157932 76570
rect 157996 75449 158024 76758
rect 158088 75954 158116 79716
rect 158180 79716 158254 79744
rect 158304 79792 158360 79801
rect 158304 79727 158360 79736
rect 158410 79744 158438 80036
rect 158502 79937 158530 80036
rect 158488 79928 158544 79937
rect 158488 79863 158544 79872
rect 158594 79744 158622 80036
rect 158686 79966 158714 80036
rect 158778 79966 158806 80036
rect 158674 79960 158726 79966
rect 158674 79902 158726 79908
rect 158766 79960 158818 79966
rect 158766 79902 158818 79908
rect 158870 79812 158898 80036
rect 158410 79716 158484 79744
rect 158076 75948 158128 75954
rect 158076 75890 158128 75896
rect 157982 75440 158038 75449
rect 157982 75375 158038 75384
rect 157984 75336 158036 75342
rect 157984 75278 158036 75284
rect 157996 62966 158024 75278
rect 158180 73982 158208 79716
rect 158258 79656 158314 79665
rect 158258 79591 158314 79600
rect 158352 79620 158404 79626
rect 158272 75682 158300 79591
rect 158352 79562 158404 79568
rect 158364 77722 158392 79562
rect 158352 77716 158404 77722
rect 158352 77658 158404 77664
rect 158456 76537 158484 79716
rect 158548 79716 158622 79744
rect 158732 79784 158898 79812
rect 158548 76673 158576 79716
rect 158628 79620 158680 79626
rect 158628 79562 158680 79568
rect 158640 77790 158668 79562
rect 158628 77784 158680 77790
rect 158628 77726 158680 77732
rect 158628 77036 158680 77042
rect 158628 76978 158680 76984
rect 158534 76664 158590 76673
rect 158534 76599 158590 76608
rect 158442 76528 158498 76537
rect 158442 76463 158498 76472
rect 158444 76152 158496 76158
rect 158444 76094 158496 76100
rect 158260 75676 158312 75682
rect 158260 75618 158312 75624
rect 158456 73982 158484 76094
rect 158168 73976 158220 73982
rect 158168 73918 158220 73924
rect 158444 73976 158496 73982
rect 158444 73918 158496 73924
rect 158640 64874 158668 76978
rect 158732 76566 158760 79784
rect 158962 79744 158990 80036
rect 159054 79971 159082 80036
rect 159040 79962 159096 79971
rect 159040 79897 159096 79906
rect 159146 79778 159174 80036
rect 159238 79898 159266 80036
rect 159226 79892 159278 79898
rect 159226 79834 159278 79840
rect 158824 79716 158990 79744
rect 159100 79750 159174 79778
rect 158720 76560 158772 76566
rect 158720 76502 158772 76508
rect 158720 72956 158772 72962
rect 158720 72898 158772 72904
rect 158548 64846 158668 64874
rect 157984 62960 158036 62966
rect 157984 62902 158036 62908
rect 157892 61464 157944 61470
rect 157892 61406 157944 61412
rect 157800 17604 157852 17610
rect 157800 17546 157852 17552
rect 157708 17536 157760 17542
rect 157708 17478 157760 17484
rect 157616 13252 157668 13258
rect 157616 13194 157668 13200
rect 157524 11892 157576 11898
rect 157524 11834 157576 11840
rect 157432 11824 157484 11830
rect 157432 11766 157484 11772
rect 156144 10396 156196 10402
rect 156144 10338 156196 10344
rect 155960 7812 156012 7818
rect 155960 7754 156012 7760
rect 158548 6526 158576 64846
rect 158536 6520 158588 6526
rect 158536 6462 158588 6468
rect 158732 6390 158760 72898
rect 158824 13190 158852 79716
rect 158994 79656 159050 79665
rect 158904 79620 158956 79626
rect 158994 79591 159050 79600
rect 158904 79562 158956 79568
rect 158916 78674 158944 79562
rect 159008 79218 159036 79591
rect 158996 79212 159048 79218
rect 158996 79154 159048 79160
rect 159100 78962 159128 79750
rect 159330 79744 159358 80036
rect 159422 79898 159450 80036
rect 159410 79892 159462 79898
rect 159410 79834 159462 79840
rect 159514 79778 159542 80036
rect 159606 79966 159634 80036
rect 159594 79960 159646 79966
rect 159594 79902 159646 79908
rect 159468 79750 159542 79778
rect 159330 79716 159404 79744
rect 159180 79688 159232 79694
rect 159180 79630 159232 79636
rect 159008 78934 159128 78962
rect 158904 78668 158956 78674
rect 158904 78610 158956 78616
rect 158904 78124 158956 78130
rect 158904 78066 158956 78072
rect 158916 14550 158944 78066
rect 159008 75750 159036 78934
rect 159192 77858 159220 79630
rect 159180 77852 159232 77858
rect 159180 77794 159232 77800
rect 159376 76786 159404 79716
rect 159468 79506 159496 79750
rect 159698 79744 159726 80036
rect 159790 79966 159818 80036
rect 159778 79960 159830 79966
rect 159778 79902 159830 79908
rect 159882 79744 159910 80036
rect 159974 79937 160002 80036
rect 159960 79928 160016 79937
rect 159960 79863 160016 79872
rect 160066 79812 160094 80036
rect 159652 79716 159726 79744
rect 159836 79716 159910 79744
rect 160020 79784 160094 79812
rect 159468 79478 159588 79506
rect 159456 79416 159508 79422
rect 159456 79358 159508 79364
rect 159100 76758 159404 76786
rect 158996 75744 159048 75750
rect 158996 75686 159048 75692
rect 158996 73772 159048 73778
rect 158996 73714 159048 73720
rect 159008 72962 159036 73714
rect 158996 72956 159048 72962
rect 158996 72898 159048 72904
rect 159100 60042 159128 76758
rect 159468 76650 159496 79358
rect 159560 78130 159588 79478
rect 159548 78124 159600 78130
rect 159548 78066 159600 78072
rect 159652 78010 159680 79716
rect 159732 79620 159784 79626
rect 159732 79562 159784 79568
rect 159744 78033 159772 79562
rect 159192 76622 159496 76650
rect 159560 77982 159680 78010
rect 159730 78024 159786 78033
rect 159192 67114 159220 76622
rect 159272 76560 159324 76566
rect 159272 76502 159324 76508
rect 159284 68406 159312 76502
rect 159560 75614 159588 77982
rect 159730 77959 159786 77968
rect 159640 77920 159692 77926
rect 159640 77862 159692 77868
rect 159652 76634 159680 77862
rect 159640 76628 159692 76634
rect 159640 76570 159692 76576
rect 159548 75608 159600 75614
rect 159548 75550 159600 75556
rect 159640 74860 159692 74866
rect 159640 74802 159692 74808
rect 159652 70394 159680 74802
rect 159836 73778 159864 79716
rect 159914 79656 159970 79665
rect 160020 79626 160048 79784
rect 160158 79744 160186 80036
rect 160112 79716 160186 79744
rect 159914 79591 159916 79600
rect 159968 79591 159970 79600
rect 160008 79620 160060 79626
rect 159916 79562 159968 79568
rect 160008 79562 160060 79568
rect 159916 79484 159968 79490
rect 159916 79426 159968 79432
rect 159824 73772 159876 73778
rect 159824 73714 159876 73720
rect 159928 73154 159956 79426
rect 160008 79416 160060 79422
rect 160008 79358 160060 79364
rect 160020 76265 160048 79358
rect 160112 78849 160140 79716
rect 160250 79676 160278 80036
rect 160342 79898 160370 80036
rect 160330 79892 160382 79898
rect 160330 79834 160382 79840
rect 160434 79744 160462 80036
rect 160526 79812 160554 80036
rect 160618 79966 160646 80036
rect 160710 79971 160738 80036
rect 160606 79960 160658 79966
rect 160606 79902 160658 79908
rect 160696 79962 160752 79971
rect 160696 79897 160752 79906
rect 160802 79830 160830 80036
rect 160894 79937 160922 80036
rect 160880 79928 160936 79937
rect 160880 79863 160936 79872
rect 160652 79824 160704 79830
rect 160526 79784 160600 79812
rect 160434 79716 160508 79744
rect 160204 79648 160278 79676
rect 160374 79656 160430 79665
rect 160098 78840 160154 78849
rect 160098 78775 160154 78784
rect 160204 76616 160232 79648
rect 160374 79591 160376 79600
rect 160428 79591 160430 79600
rect 160376 79562 160428 79568
rect 160284 79552 160336 79558
rect 160284 79494 160336 79500
rect 160296 77353 160324 79494
rect 160374 79112 160430 79121
rect 160374 79047 160430 79056
rect 160282 77344 160338 77353
rect 160282 77279 160338 77288
rect 160112 76588 160232 76616
rect 160006 76256 160062 76265
rect 160006 76191 160062 76200
rect 159928 73126 160048 73154
rect 159652 70366 159772 70394
rect 159272 68400 159324 68406
rect 159272 68342 159324 68348
rect 159180 67108 159232 67114
rect 159180 67050 159232 67056
rect 159088 60036 159140 60042
rect 159088 59978 159140 59984
rect 159744 35222 159772 70366
rect 159732 35216 159784 35222
rect 159732 35158 159784 35164
rect 160020 32706 160048 73126
rect 160008 32700 160060 32706
rect 160008 32642 160060 32648
rect 158904 14544 158956 14550
rect 158904 14486 158956 14492
rect 158812 13184 158864 13190
rect 158812 13126 158864 13132
rect 160112 7750 160140 76588
rect 160284 76560 160336 76566
rect 160284 76502 160336 76508
rect 160192 75200 160244 75206
rect 160192 75142 160244 75148
rect 160204 13122 160232 75142
rect 160296 17406 160324 76502
rect 160388 76401 160416 79047
rect 160374 76392 160430 76401
rect 160374 76327 160430 76336
rect 160376 76152 160428 76158
rect 160376 76094 160428 76100
rect 160388 18834 160416 76094
rect 160480 18902 160508 79716
rect 160572 76566 160600 79784
rect 160652 79766 160704 79772
rect 160790 79824 160842 79830
rect 160986 79778 161014 80036
rect 161078 79830 161106 80036
rect 160790 79766 160842 79772
rect 160560 76560 160612 76566
rect 160560 76502 160612 76508
rect 160560 76220 160612 76226
rect 160560 76162 160612 76168
rect 160572 20058 160600 76162
rect 160664 21622 160692 79766
rect 160940 79750 161014 79778
rect 161066 79824 161118 79830
rect 161066 79766 161118 79772
rect 160836 79688 160888 79694
rect 160742 79656 160798 79665
rect 160836 79630 160888 79636
rect 160742 79591 160798 79600
rect 160756 76158 160784 79591
rect 160744 76152 160796 76158
rect 160744 76094 160796 76100
rect 160848 75206 160876 79630
rect 160940 76226 160968 79750
rect 161170 79744 161198 80036
rect 161262 79937 161290 80036
rect 161354 79966 161382 80036
rect 161342 79960 161394 79966
rect 161248 79928 161304 79937
rect 161342 79902 161394 79908
rect 161248 79863 161304 79872
rect 161446 79744 161474 80036
rect 161170 79716 161244 79744
rect 161112 79620 161164 79626
rect 161112 79562 161164 79568
rect 161020 79552 161072 79558
rect 161020 79494 161072 79500
rect 161032 78878 161060 79494
rect 161020 78872 161072 78878
rect 161020 78814 161072 78820
rect 161020 78192 161072 78198
rect 161020 78134 161072 78140
rect 160928 76220 160980 76226
rect 160928 76162 160980 76168
rect 160836 75200 160888 75206
rect 160836 75142 160888 75148
rect 161032 67250 161060 78134
rect 161124 76537 161152 79562
rect 161216 78470 161244 79716
rect 161400 79716 161474 79744
rect 161538 79744 161566 80036
rect 161630 79937 161658 80036
rect 161616 79928 161672 79937
rect 161616 79863 161672 79872
rect 161722 79812 161750 80036
rect 161676 79784 161750 79812
rect 161538 79716 161612 79744
rect 161296 79688 161348 79694
rect 161296 79630 161348 79636
rect 161204 78464 161256 78470
rect 161204 78406 161256 78412
rect 161308 77926 161336 79630
rect 161296 77920 161348 77926
rect 161296 77862 161348 77868
rect 161400 76673 161428 79716
rect 161480 79620 161532 79626
rect 161480 79562 161532 79568
rect 161386 76664 161442 76673
rect 161386 76599 161442 76608
rect 161110 76528 161166 76537
rect 161110 76463 161166 76472
rect 161020 67244 161072 67250
rect 161020 67186 161072 67192
rect 160652 21616 160704 21622
rect 160652 21558 160704 21564
rect 160560 20052 160612 20058
rect 160560 19994 160612 20000
rect 160558 19952 160614 19961
rect 160558 19887 160614 19896
rect 160468 18896 160520 18902
rect 160468 18838 160520 18844
rect 160376 18828 160428 18834
rect 160376 18770 160428 18776
rect 160284 17400 160336 17406
rect 160284 17342 160336 17348
rect 160192 13116 160244 13122
rect 160192 13058 160244 13064
rect 160100 7744 160152 7750
rect 160100 7686 160152 7692
rect 160572 6914 160600 19887
rect 160112 6886 160600 6914
rect 158720 6384 158772 6390
rect 158720 6326 158772 6332
rect 156604 6248 156656 6254
rect 156604 6190 156656 6196
rect 154488 5092 154540 5098
rect 154488 5034 154540 5040
rect 152556 3800 152608 3806
rect 152556 3742 152608 3748
rect 154212 3732 154264 3738
rect 154212 3674 154264 3680
rect 153016 3324 153068 3330
rect 153016 3266 153068 3272
rect 153028 480 153056 3266
rect 154224 480 154252 3674
rect 155408 3664 155460 3670
rect 155408 3606 155460 3612
rect 155420 480 155448 3606
rect 156616 480 156644 6190
rect 157800 4888 157852 4894
rect 157800 4830 157852 4836
rect 158902 4856 158958 4865
rect 157812 480 157840 4830
rect 158902 4791 158958 4800
rect 158916 480 158944 4791
rect 160112 480 160140 6886
rect 161492 6322 161520 79562
rect 161584 76566 161612 79716
rect 161676 78266 161704 79784
rect 161814 79744 161842 80036
rect 161906 79966 161934 80036
rect 161998 79966 162026 80036
rect 161894 79960 161946 79966
rect 161894 79902 161946 79908
rect 161986 79960 162038 79966
rect 161986 79902 162038 79908
rect 162090 79812 162118 80036
rect 161768 79716 161842 79744
rect 161938 79792 161994 79801
rect 161938 79727 161994 79736
rect 162044 79784 162118 79812
rect 161664 78260 161716 78266
rect 161664 78202 161716 78208
rect 161572 76560 161624 76566
rect 161572 76502 161624 76508
rect 161572 75948 161624 75954
rect 161572 75890 161624 75896
rect 161584 7682 161612 75890
rect 161664 73636 161716 73642
rect 161664 73578 161716 73584
rect 161676 9110 161704 73578
rect 161768 19990 161796 79716
rect 161848 79620 161900 79626
rect 161848 79562 161900 79568
rect 161860 75410 161888 79562
rect 161848 75404 161900 75410
rect 161848 75346 161900 75352
rect 161848 74792 161900 74798
rect 161848 74734 161900 74740
rect 161860 21554 161888 74734
rect 161952 32638 161980 79727
rect 162044 75954 162072 79784
rect 162182 79744 162210 80036
rect 162274 79898 162302 80036
rect 162262 79892 162314 79898
rect 162262 79834 162314 79840
rect 162366 79744 162394 80036
rect 162458 79937 162486 80036
rect 162444 79928 162500 79937
rect 162550 79898 162578 80036
rect 162444 79863 162500 79872
rect 162538 79892 162590 79898
rect 162538 79834 162590 79840
rect 162642 79801 162670 80036
rect 162734 79966 162762 80036
rect 162722 79960 162774 79966
rect 162722 79902 162774 79908
rect 162628 79792 162684 79801
rect 162136 79716 162210 79744
rect 162320 79716 162394 79744
rect 162492 79756 162544 79762
rect 162032 75948 162084 75954
rect 162032 75890 162084 75896
rect 162136 73642 162164 79716
rect 162214 79656 162270 79665
rect 162214 79591 162270 79600
rect 162228 77246 162256 79591
rect 162216 77240 162268 77246
rect 162216 77182 162268 77188
rect 162216 76560 162268 76566
rect 162216 76502 162268 76508
rect 162124 73636 162176 73642
rect 162124 73578 162176 73584
rect 162228 70394 162256 76502
rect 162320 74798 162348 79716
rect 162826 79744 162854 80036
rect 162918 79801 162946 80036
rect 163010 79966 163038 80036
rect 162998 79960 163050 79966
rect 162998 79902 163050 79908
rect 162628 79727 162684 79736
rect 162492 79698 162544 79704
rect 162780 79716 162854 79744
rect 162904 79792 162960 79801
rect 163102 79744 163130 80036
rect 162904 79727 162960 79736
rect 163056 79716 163130 79744
rect 163194 79744 163222 80036
rect 163286 79937 163314 80036
rect 163272 79928 163328 79937
rect 163378 79898 163406 80036
rect 163272 79863 163328 79872
rect 163366 79892 163418 79898
rect 163366 79834 163418 79840
rect 163318 79792 163374 79801
rect 163194 79716 163268 79744
rect 163470 79744 163498 80036
rect 163318 79727 163374 79736
rect 162400 78328 162452 78334
rect 162400 78270 162452 78276
rect 162308 74792 162360 74798
rect 162308 74734 162360 74740
rect 162044 70366 162256 70394
rect 162044 67046 162072 70366
rect 162032 67040 162084 67046
rect 162032 66982 162084 66988
rect 162412 64874 162440 78270
rect 162504 78130 162532 79698
rect 162676 79688 162728 79694
rect 162674 79656 162676 79665
rect 162728 79656 162730 79665
rect 162674 79591 162730 79600
rect 162780 78577 162808 79716
rect 162860 79620 162912 79626
rect 162860 79562 162912 79568
rect 162766 78568 162822 78577
rect 162766 78503 162822 78512
rect 162492 78124 162544 78130
rect 162492 78066 162544 78072
rect 162674 77616 162730 77625
rect 162674 77551 162730 77560
rect 162688 73154 162716 77551
rect 162768 77036 162820 77042
rect 162768 76978 162820 76984
rect 162780 76294 162808 76978
rect 162768 76288 162820 76294
rect 162768 76230 162820 76236
rect 162688 73126 162808 73154
rect 162780 70394 162808 73126
rect 162872 72729 162900 79562
rect 162952 79552 163004 79558
rect 162952 79494 163004 79500
rect 162858 72720 162914 72729
rect 162858 72655 162914 72664
rect 162228 64846 162440 64874
rect 162504 70366 162808 70394
rect 162228 64258 162256 64846
rect 162216 64252 162268 64258
rect 162216 64194 162268 64200
rect 162504 42090 162532 70366
rect 162492 42084 162544 42090
rect 162492 42026 162544 42032
rect 161940 32632 161992 32638
rect 161940 32574 161992 32580
rect 161848 21548 161900 21554
rect 161848 21490 161900 21496
rect 162860 20120 162912 20126
rect 162860 20062 162912 20068
rect 161756 19984 161808 19990
rect 161756 19926 161808 19932
rect 161664 9104 161716 9110
rect 161664 9046 161716 9052
rect 161572 7676 161624 7682
rect 161572 7618 161624 7624
rect 161480 6316 161532 6322
rect 161480 6258 161532 6264
rect 162492 6180 162544 6186
rect 162492 6122 162544 6128
rect 161294 3360 161350 3369
rect 161294 3295 161350 3304
rect 161308 480 161336 3295
rect 162504 480 162532 6122
rect 162872 3482 162900 20062
rect 162964 4962 162992 79494
rect 163056 76566 163084 79716
rect 163136 79620 163188 79626
rect 163136 79562 163188 79568
rect 163044 76560 163096 76566
rect 163044 76502 163096 76508
rect 163044 76288 163096 76294
rect 163044 76230 163096 76236
rect 163056 9042 163084 76230
rect 163148 10334 163176 79562
rect 163240 79490 163268 79716
rect 163228 79484 163280 79490
rect 163228 79426 163280 79432
rect 163228 79348 163280 79354
rect 163228 79290 163280 79296
rect 163240 78674 163268 79290
rect 163228 78668 163280 78674
rect 163228 78610 163280 78616
rect 163228 76356 163280 76362
rect 163228 76298 163280 76304
rect 163240 17338 163268 76298
rect 163332 21486 163360 79727
rect 163424 79716 163498 79744
rect 163562 79744 163590 80036
rect 163654 79966 163682 80036
rect 163642 79960 163694 79966
rect 163642 79902 163694 79908
rect 163746 79744 163774 80036
rect 163838 79898 163866 80036
rect 163826 79892 163878 79898
rect 163826 79834 163878 79840
rect 163930 79744 163958 80036
rect 164022 79937 164050 80036
rect 164008 79928 164064 79937
rect 164008 79863 164064 79872
rect 164114 79812 164142 80036
rect 163562 79716 163636 79744
rect 163746 79716 163820 79744
rect 163424 79558 163452 79716
rect 163504 79620 163556 79626
rect 163504 79562 163556 79568
rect 163412 79552 163464 79558
rect 163412 79494 163464 79500
rect 163412 79348 163464 79354
rect 163412 79290 163464 79296
rect 163424 78713 163452 79290
rect 163410 78704 163466 78713
rect 163410 78639 163466 78648
rect 163412 76560 163464 76566
rect 163412 76502 163464 76508
rect 163424 32570 163452 76502
rect 163516 57322 163544 79562
rect 163608 62898 163636 79716
rect 163688 79620 163740 79626
rect 163688 79562 163740 79568
rect 163700 76294 163728 79562
rect 163688 76288 163740 76294
rect 163688 76230 163740 76236
rect 163792 70394 163820 79716
rect 163884 79716 163958 79744
rect 164068 79784 164142 79812
rect 163884 76362 163912 79716
rect 163962 79656 164018 79665
rect 163962 79591 164018 79600
rect 163976 78062 164004 79591
rect 164068 79121 164096 79784
rect 164206 79744 164234 80036
rect 164160 79716 164234 79744
rect 164298 79744 164326 80036
rect 164390 79898 164418 80036
rect 164378 79892 164430 79898
rect 164378 79834 164430 79840
rect 164482 79744 164510 80036
rect 164574 79937 164602 80036
rect 164560 79928 164616 79937
rect 164560 79863 164616 79872
rect 164666 79812 164694 80036
rect 164758 79966 164786 80036
rect 164746 79960 164798 79966
rect 164746 79902 164798 79908
rect 164666 79784 164740 79812
rect 164298 79716 164372 79744
rect 164482 79716 164556 79744
rect 164160 79665 164188 79716
rect 164146 79656 164202 79665
rect 164146 79591 164202 79600
rect 164240 79620 164292 79626
rect 164240 79562 164292 79568
rect 164148 79280 164200 79286
rect 164148 79222 164200 79228
rect 164054 79112 164110 79121
rect 164054 79047 164110 79056
rect 164056 79008 164108 79014
rect 164056 78950 164108 78956
rect 164068 78402 164096 78950
rect 164056 78396 164108 78402
rect 164056 78338 164108 78344
rect 163964 78056 164016 78062
rect 163964 77998 164016 78004
rect 164160 77518 164188 79222
rect 164148 77512 164200 77518
rect 164148 77454 164200 77460
rect 163872 76356 163924 76362
rect 163872 76298 163924 76304
rect 163792 70366 164004 70394
rect 163596 62892 163648 62898
rect 163596 62834 163648 62840
rect 163504 57316 163556 57322
rect 163504 57258 163556 57264
rect 163412 32564 163464 32570
rect 163412 32506 163464 32512
rect 163320 21480 163372 21486
rect 163320 21422 163372 21428
rect 163228 17332 163280 17338
rect 163228 17274 163280 17280
rect 163136 10328 163188 10334
rect 163136 10270 163188 10276
rect 163044 9036 163096 9042
rect 163044 8978 163096 8984
rect 162952 4956 163004 4962
rect 162952 4898 163004 4904
rect 163976 3738 164004 70366
rect 164252 7614 164280 79562
rect 164344 79422 164372 79716
rect 164332 79416 164384 79422
rect 164332 79358 164384 79364
rect 164422 79384 164478 79393
rect 164422 79319 164478 79328
rect 164332 79144 164384 79150
rect 164436 79121 164464 79319
rect 164332 79086 164384 79092
rect 164422 79112 164478 79121
rect 164344 78538 164372 79086
rect 164422 79047 164478 79056
rect 164332 78532 164384 78538
rect 164332 78474 164384 78480
rect 164528 77518 164556 79716
rect 164608 79688 164660 79694
rect 164608 79630 164660 79636
rect 164516 77512 164568 77518
rect 164516 77454 164568 77460
rect 164422 76664 164478 76673
rect 164422 76599 164478 76608
rect 164332 76560 164384 76566
rect 164332 76502 164384 76508
rect 164344 14482 164372 76502
rect 164436 21418 164464 76599
rect 164516 76356 164568 76362
rect 164516 76298 164568 76304
rect 164528 23050 164556 76298
rect 164620 23118 164648 79630
rect 164712 76566 164740 79784
rect 164850 79744 164878 80036
rect 164942 79937 164970 80036
rect 164928 79928 164984 79937
rect 164928 79863 164984 79872
rect 165034 79812 165062 80036
rect 164988 79784 165062 79812
rect 164850 79716 164924 79744
rect 164790 79248 164846 79257
rect 164790 79183 164846 79192
rect 164804 79082 164832 79183
rect 164792 79076 164844 79082
rect 164792 79018 164844 79024
rect 164792 78464 164844 78470
rect 164792 78406 164844 78412
rect 164804 78305 164832 78406
rect 164790 78296 164846 78305
rect 164790 78231 164846 78240
rect 164792 77376 164844 77382
rect 164792 77318 164844 77324
rect 164700 76560 164752 76566
rect 164700 76502 164752 76508
rect 164804 76294 164832 77318
rect 164792 76288 164844 76294
rect 164792 76230 164844 76236
rect 164792 75744 164844 75750
rect 164792 75686 164844 75692
rect 164804 75546 164832 75686
rect 164792 75540 164844 75546
rect 164792 75482 164844 75488
rect 164700 74996 164752 75002
rect 164700 74938 164752 74944
rect 164712 26926 164740 74938
rect 164792 73840 164844 73846
rect 164792 73782 164844 73788
rect 164804 57254 164832 73782
rect 164896 69834 164924 79716
rect 164988 75002 165016 79784
rect 165126 79744 165154 80036
rect 165218 79830 165246 80036
rect 165206 79824 165258 79830
rect 165310 79801 165338 80036
rect 165206 79766 165258 79772
rect 165296 79792 165352 79801
rect 165080 79716 165154 79744
rect 165296 79727 165352 79736
rect 165402 79744 165430 80036
rect 165494 79812 165522 80036
rect 165586 79937 165614 80036
rect 165572 79928 165628 79937
rect 165572 79863 165628 79872
rect 165494 79784 165568 79812
rect 165402 79716 165476 79744
rect 164976 74996 165028 75002
rect 164976 74938 165028 74944
rect 165080 73846 165108 79716
rect 165250 79656 165306 79665
rect 165250 79591 165306 79600
rect 165344 79620 165396 79626
rect 165160 79076 165212 79082
rect 165160 79018 165212 79024
rect 165172 78606 165200 79018
rect 165160 78600 165212 78606
rect 165160 78542 165212 78548
rect 165158 78296 165214 78305
rect 165158 78231 165214 78240
rect 165172 77897 165200 78231
rect 165158 77888 165214 77897
rect 165158 77823 165214 77832
rect 165160 77308 165212 77314
rect 165160 77250 165212 77256
rect 165172 73846 165200 77250
rect 165068 73840 165120 73846
rect 165068 73782 165120 73788
rect 165160 73840 165212 73846
rect 165160 73782 165212 73788
rect 165264 72418 165292 79591
rect 165344 79562 165396 79568
rect 165356 76362 165384 79562
rect 165448 76673 165476 79716
rect 165434 76664 165490 76673
rect 165434 76599 165490 76608
rect 165540 76537 165568 79784
rect 165678 79744 165706 80036
rect 165770 79898 165798 80036
rect 165758 79892 165810 79898
rect 165758 79834 165810 79840
rect 165862 79812 165890 80036
rect 165954 79937 165982 80036
rect 166046 79966 166074 80036
rect 166138 79966 166166 80036
rect 166230 79966 166258 80036
rect 166034 79960 166086 79966
rect 165940 79928 165996 79937
rect 166034 79902 166086 79908
rect 166126 79960 166178 79966
rect 166126 79902 166178 79908
rect 166218 79960 166270 79966
rect 166218 79902 166270 79908
rect 166322 79898 166350 80036
rect 165940 79863 165996 79872
rect 166310 79892 166362 79898
rect 166310 79834 166362 79840
rect 165988 79824 166040 79830
rect 165862 79801 165936 79812
rect 165862 79792 165950 79801
rect 165862 79784 165894 79792
rect 165678 79716 165752 79744
rect 165988 79766 166040 79772
rect 165894 79727 165950 79736
rect 165620 79620 165672 79626
rect 165620 79562 165672 79568
rect 165526 76528 165582 76537
rect 165526 76463 165582 76472
rect 165344 76356 165396 76362
rect 165344 76298 165396 76304
rect 165252 72412 165304 72418
rect 165252 72354 165304 72360
rect 164884 69828 164936 69834
rect 164884 69770 164936 69776
rect 164792 57248 164844 57254
rect 164792 57190 164844 57196
rect 164700 26920 164752 26926
rect 164700 26862 164752 26868
rect 164608 23112 164660 23118
rect 164608 23054 164660 23060
rect 164516 23044 164568 23050
rect 164516 22986 164568 22992
rect 164424 21412 164476 21418
rect 164424 21354 164476 21360
rect 164332 14476 164384 14482
rect 164332 14418 164384 14424
rect 164240 7608 164292 7614
rect 164240 7550 164292 7556
rect 165632 4894 165660 79562
rect 165724 78402 165752 79716
rect 165896 79688 165948 79694
rect 165896 79630 165948 79636
rect 165804 79552 165856 79558
rect 165804 79494 165856 79500
rect 165712 78396 165764 78402
rect 165712 78338 165764 78344
rect 165712 76560 165764 76566
rect 165712 76502 165764 76508
rect 165620 4888 165672 4894
rect 165620 4830 165672 4836
rect 165724 4826 165752 76502
rect 165816 11762 165844 79494
rect 165908 22982 165936 79630
rect 165896 22976 165948 22982
rect 165896 22918 165948 22924
rect 166000 22914 166028 79766
rect 166080 79756 166132 79762
rect 166414 79744 166442 80036
rect 166132 79716 166212 79744
rect 166080 79698 166132 79704
rect 166078 79656 166134 79665
rect 166078 79591 166134 79600
rect 166092 25770 166120 79591
rect 166184 29714 166212 79716
rect 166276 79716 166442 79744
rect 166506 79744 166534 80036
rect 166598 79812 166626 80036
rect 166690 79966 166718 80036
rect 166678 79960 166730 79966
rect 166782 79937 166810 80036
rect 166678 79902 166730 79908
rect 166768 79928 166824 79937
rect 166768 79863 166824 79872
rect 166598 79784 166764 79812
rect 166506 79716 166580 79744
rect 166276 31074 166304 79716
rect 166448 79484 166500 79490
rect 166448 79426 166500 79432
rect 166354 78840 166410 78849
rect 166354 78775 166356 78784
rect 166408 78775 166410 78784
rect 166356 78746 166408 78752
rect 166460 78606 166488 79426
rect 166448 78600 166500 78606
rect 166448 78542 166500 78548
rect 166448 77512 166500 77518
rect 166448 77454 166500 77460
rect 166460 75274 166488 77454
rect 166448 75268 166500 75274
rect 166448 75210 166500 75216
rect 166552 71774 166580 79716
rect 166630 79656 166686 79665
rect 166630 79591 166686 79600
rect 166460 71746 166580 71774
rect 166460 70394 166488 71746
rect 166368 70366 166488 70394
rect 166368 61402 166396 70366
rect 166644 69766 166672 79591
rect 166736 76566 166764 79784
rect 166874 79744 166902 80036
rect 166966 79801 166994 80036
rect 166828 79716 166902 79744
rect 166952 79792 167008 79801
rect 166952 79727 167008 79736
rect 167058 79744 167086 80036
rect 167150 79937 167178 80036
rect 167136 79928 167192 79937
rect 167136 79863 167192 79872
rect 167242 79812 167270 80036
rect 167334 79937 167362 80036
rect 167320 79928 167376 79937
rect 167320 79863 167376 79872
rect 167242 79784 167316 79812
rect 167058 79716 167132 79744
rect 166828 76673 166856 79716
rect 166908 79620 166960 79626
rect 166908 79562 166960 79568
rect 167000 79620 167052 79626
rect 167000 79562 167052 79568
rect 166814 76664 166870 76673
rect 166814 76599 166870 76608
rect 166724 76560 166776 76566
rect 166724 76502 166776 76508
rect 166920 75177 166948 79562
rect 166906 75168 166962 75177
rect 166906 75103 166962 75112
rect 166632 69760 166684 69766
rect 166632 69702 166684 69708
rect 166356 61396 166408 61402
rect 166356 61338 166408 61344
rect 166264 31068 166316 31074
rect 166264 31010 166316 31016
rect 166172 29708 166224 29714
rect 166172 29650 166224 29656
rect 166080 25764 166132 25770
rect 166080 25706 166132 25712
rect 165988 22908 166040 22914
rect 165988 22850 166040 22856
rect 167012 15910 167040 79562
rect 167104 77314 167132 79716
rect 167182 79656 167238 79665
rect 167182 79591 167238 79600
rect 167092 77308 167144 77314
rect 167092 77250 167144 77256
rect 167092 72140 167144 72146
rect 167092 72082 167144 72088
rect 167104 17270 167132 72082
rect 167196 24342 167224 79591
rect 167184 24336 167236 24342
rect 167184 24278 167236 24284
rect 167288 24274 167316 79784
rect 167426 79778 167454 80036
rect 167518 79971 167546 80036
rect 167504 79962 167560 79971
rect 167610 79966 167638 80036
rect 167702 79966 167730 80036
rect 167794 79966 167822 80036
rect 167886 79966 167914 80036
rect 167504 79897 167560 79906
rect 167598 79960 167650 79966
rect 167598 79902 167650 79908
rect 167690 79960 167742 79966
rect 167690 79902 167742 79908
rect 167782 79960 167834 79966
rect 167782 79902 167834 79908
rect 167874 79960 167926 79966
rect 167874 79902 167926 79908
rect 167380 79750 167454 79778
rect 167276 24268 167328 24274
rect 167276 24210 167328 24216
rect 167380 24206 167408 79750
rect 167552 79688 167604 79694
rect 167552 79630 167604 79636
rect 167736 79688 167788 79694
rect 167736 79630 167788 79636
rect 167460 79620 167512 79626
rect 167460 79562 167512 79568
rect 167472 29646 167500 79562
rect 167564 76566 167592 79630
rect 167644 79416 167696 79422
rect 167644 79358 167696 79364
rect 167656 77994 167684 79358
rect 167644 77988 167696 77994
rect 167644 77930 167696 77936
rect 167748 76650 167776 79630
rect 167978 79608 168006 80036
rect 168070 79676 168098 80036
rect 168162 79966 168190 80036
rect 168150 79960 168202 79966
rect 168150 79902 168202 79908
rect 168254 79778 168282 80036
rect 168346 79966 168374 80036
rect 168438 79971 168466 80036
rect 168334 79960 168386 79966
rect 168334 79902 168386 79908
rect 168424 79962 168480 79971
rect 168424 79897 168480 79906
rect 168530 79898 168558 80036
rect 168622 79898 168650 80036
rect 168518 79892 168570 79898
rect 168518 79834 168570 79840
rect 168610 79892 168662 79898
rect 168610 79834 168662 79840
rect 168562 79792 168618 79801
rect 168254 79750 168328 79778
rect 168196 79688 168248 79694
rect 168070 79648 168144 79676
rect 167978 79580 168052 79608
rect 167828 79552 167880 79558
rect 167828 79494 167880 79500
rect 167656 76622 167776 76650
rect 167552 76560 167604 76566
rect 167552 76502 167604 76508
rect 167550 76392 167606 76401
rect 167550 76327 167606 76336
rect 167564 32502 167592 76327
rect 167656 66910 167684 76622
rect 167736 76560 167788 76566
rect 167736 76502 167788 76508
rect 167748 66978 167776 76502
rect 167840 75342 167868 79494
rect 167920 77240 167972 77246
rect 167920 77182 167972 77188
rect 167932 76566 167960 77182
rect 167920 76560 167972 76566
rect 167920 76502 167972 76508
rect 167828 75336 167880 75342
rect 167828 75278 167880 75284
rect 168024 72146 168052 79580
rect 168116 78713 168144 79648
rect 168300 79665 168328 79750
rect 168380 79756 168432 79762
rect 168714 79778 168742 80036
rect 168806 79966 168834 80036
rect 168794 79960 168846 79966
rect 168794 79902 168846 79908
rect 168898 79898 168926 80036
rect 168990 79966 169018 80036
rect 168978 79960 169030 79966
rect 168978 79902 169030 79908
rect 169082 79898 169110 80036
rect 169174 79898 169202 80036
rect 168886 79892 168938 79898
rect 168886 79834 168938 79840
rect 169070 79892 169122 79898
rect 169070 79834 169122 79840
rect 169162 79892 169214 79898
rect 169162 79834 169214 79840
rect 168562 79727 168618 79736
rect 168668 79750 168742 79778
rect 168932 79756 168984 79762
rect 168380 79698 168432 79704
rect 168196 79630 168248 79636
rect 168286 79656 168342 79665
rect 168102 78704 168158 78713
rect 168102 78639 168158 78648
rect 168208 76673 168236 79630
rect 168286 79591 168342 79600
rect 168288 79552 168340 79558
rect 168288 79494 168340 79500
rect 168300 77382 168328 79494
rect 168288 77376 168340 77382
rect 168288 77318 168340 77324
rect 168288 77240 168340 77246
rect 168288 77182 168340 77188
rect 168194 76664 168250 76673
rect 168194 76599 168250 76608
rect 168300 73154 168328 77182
rect 168392 76362 168420 79698
rect 168472 79688 168524 79694
rect 168472 79630 168524 79636
rect 168380 76356 168432 76362
rect 168380 76298 168432 76304
rect 168300 73126 168420 73154
rect 168012 72140 168064 72146
rect 168012 72082 168064 72088
rect 167736 66972 167788 66978
rect 167736 66914 167788 66920
rect 167644 66904 167696 66910
rect 167644 66846 167696 66852
rect 167552 32496 167604 32502
rect 167552 32438 167604 32444
rect 167460 29640 167512 29646
rect 167460 29582 167512 29588
rect 167368 24200 167420 24206
rect 167368 24142 167420 24148
rect 168392 18698 168420 73126
rect 168484 18766 168512 79630
rect 168576 74526 168604 79727
rect 168668 78742 168696 79750
rect 168932 79698 168984 79704
rect 169024 79756 169076 79762
rect 169266 79744 169294 80036
rect 169358 79937 169386 80036
rect 169344 79928 169400 79937
rect 169344 79863 169400 79872
rect 169450 79778 169478 80036
rect 169542 79898 169570 80036
rect 169530 79892 169582 79898
rect 169530 79834 169582 79840
rect 169024 79698 169076 79704
rect 169220 79716 169294 79744
rect 169404 79750 169478 79778
rect 168748 79688 168800 79694
rect 168748 79630 168800 79636
rect 168656 78736 168708 78742
rect 168656 78678 168708 78684
rect 168760 76616 168788 79630
rect 168840 79620 168892 79626
rect 168840 79562 168892 79568
rect 168852 77246 168880 79562
rect 168840 77240 168892 77246
rect 168840 77182 168892 77188
rect 168668 76588 168788 76616
rect 168564 74520 168616 74526
rect 168564 74462 168616 74468
rect 168564 72344 168616 72350
rect 168564 72286 168616 72292
rect 168472 18760 168524 18766
rect 168472 18702 168524 18708
rect 168380 18692 168432 18698
rect 168380 18634 168432 18640
rect 168576 18630 168604 72286
rect 168668 22846 168696 76588
rect 168838 76528 168894 76537
rect 168838 76463 168894 76472
rect 168748 76356 168800 76362
rect 168748 76298 168800 76304
rect 168760 24138 168788 76298
rect 168852 25634 168880 76463
rect 168944 62830 168972 79698
rect 169036 75954 169064 79698
rect 169116 79688 169168 79694
rect 169116 79630 169168 79636
rect 169024 75948 169076 75954
rect 169024 75890 169076 75896
rect 169128 72350 169156 79630
rect 169116 72344 169168 72350
rect 169116 72286 169168 72292
rect 169220 70394 169248 79716
rect 169404 79608 169432 79750
rect 169634 79744 169662 80036
rect 169726 79812 169754 80036
rect 169818 79966 169846 80036
rect 169806 79960 169858 79966
rect 169806 79902 169858 79908
rect 169910 79812 169938 80036
rect 170002 79937 170030 80036
rect 169988 79928 170044 79937
rect 169988 79863 170044 79872
rect 169726 79784 169800 79812
rect 169588 79716 169662 79744
rect 169484 79688 169536 79694
rect 169484 79630 169536 79636
rect 169312 79580 169432 79608
rect 169312 75206 169340 79580
rect 169392 79484 169444 79490
rect 169392 79426 169444 79432
rect 169404 78849 169432 79426
rect 169390 78840 169446 78849
rect 169390 78775 169446 78784
rect 169392 77376 169444 77382
rect 169392 77318 169444 77324
rect 169404 76673 169432 77318
rect 169390 76664 169446 76673
rect 169390 76599 169446 76608
rect 169300 75200 169352 75206
rect 169300 75142 169352 75148
rect 169036 70366 169248 70394
rect 169036 64190 169064 70366
rect 169496 68338 169524 79630
rect 169588 76537 169616 79716
rect 169668 79620 169720 79626
rect 169668 79562 169720 79568
rect 169574 76528 169630 76537
rect 169574 76463 169630 76472
rect 169680 76362 169708 79562
rect 169668 76356 169720 76362
rect 169668 76298 169720 76304
rect 169772 76129 169800 79784
rect 169864 79784 169938 79812
rect 169758 76120 169814 76129
rect 169758 76055 169814 76064
rect 169864 75993 169892 79784
rect 170094 79778 170122 80036
rect 170186 79966 170214 80036
rect 170174 79960 170226 79966
rect 170174 79902 170226 79908
rect 170278 79801 170306 80036
rect 170370 79966 170398 80036
rect 170462 79966 170490 80036
rect 170358 79960 170410 79966
rect 170358 79902 170410 79908
rect 170450 79960 170502 79966
rect 170450 79902 170502 79908
rect 170554 79898 170582 80036
rect 170646 79966 170674 80036
rect 170738 79966 170766 80036
rect 170634 79960 170686 79966
rect 170634 79902 170686 79908
rect 170726 79960 170778 79966
rect 170830 79937 170858 80036
rect 170726 79902 170778 79908
rect 170816 79928 170872 79937
rect 170542 79892 170594 79898
rect 170922 79898 170950 80036
rect 171014 79898 171042 80036
rect 170816 79863 170872 79872
rect 170910 79892 170962 79898
rect 170542 79834 170594 79840
rect 170910 79834 170962 79840
rect 171002 79892 171054 79898
rect 171002 79834 171054 79840
rect 170772 79824 170824 79830
rect 170264 79792 170320 79801
rect 170094 79750 170168 79778
rect 170036 79688 170088 79694
rect 169942 79656 169998 79665
rect 170036 79630 170088 79636
rect 169942 79591 169998 79600
rect 169850 75984 169906 75993
rect 169850 75919 169906 75928
rect 169852 75880 169904 75886
rect 169758 75848 169814 75857
rect 169852 75822 169904 75828
rect 169758 75783 169814 75792
rect 169484 68332 169536 68338
rect 169484 68274 169536 68280
rect 169024 64184 169076 64190
rect 169024 64126 169076 64132
rect 168932 62824 168984 62830
rect 168932 62766 168984 62772
rect 168840 25628 168892 25634
rect 168840 25570 168892 25576
rect 168748 24132 168800 24138
rect 168748 24074 168800 24080
rect 168656 22840 168708 22846
rect 168656 22782 168708 22788
rect 168564 18624 168616 18630
rect 168564 18566 168616 18572
rect 167092 17264 167144 17270
rect 167092 17206 167144 17212
rect 167000 15904 167052 15910
rect 167000 15846 167052 15852
rect 165804 11756 165856 11762
rect 165804 11698 165856 11704
rect 169772 6254 169800 75783
rect 169760 6248 169812 6254
rect 169760 6190 169812 6196
rect 169864 6186 169892 75822
rect 169956 8974 169984 79591
rect 170048 25566 170076 79630
rect 170140 78713 170168 79750
rect 170586 79792 170642 79801
rect 170264 79727 170320 79736
rect 170404 79756 170456 79762
rect 171106 79778 171134 80036
rect 171198 79898 171226 80036
rect 171186 79892 171238 79898
rect 171186 79834 171238 79840
rect 171290 79778 171318 80036
rect 170772 79766 170824 79772
rect 170586 79727 170642 79736
rect 170404 79698 170456 79704
rect 170312 79688 170364 79694
rect 170416 79665 170444 79698
rect 170312 79630 170364 79636
rect 170402 79656 170458 79665
rect 170126 78704 170182 78713
rect 170126 78639 170182 78648
rect 170128 78532 170180 78538
rect 170128 78474 170180 78480
rect 170140 32434 170168 78474
rect 170220 77852 170272 77858
rect 170220 77794 170272 77800
rect 170232 77518 170260 77794
rect 170220 77512 170272 77518
rect 170220 77454 170272 77460
rect 170324 76265 170352 79630
rect 170402 79591 170458 79600
rect 170496 79620 170548 79626
rect 170496 79562 170548 79568
rect 170404 79552 170456 79558
rect 170404 79494 170456 79500
rect 170310 76256 170366 76265
rect 170310 76191 170366 76200
rect 170220 75132 170272 75138
rect 170220 75074 170272 75080
rect 170232 69018 170260 75074
rect 170416 71774 170444 79494
rect 170508 75886 170536 79562
rect 170600 78538 170628 79727
rect 170680 79484 170732 79490
rect 170680 79426 170732 79432
rect 170692 78849 170720 79426
rect 170678 78840 170734 78849
rect 170678 78775 170734 78784
rect 170588 78532 170640 78538
rect 170588 78474 170640 78480
rect 170680 75948 170732 75954
rect 170680 75890 170732 75896
rect 170496 75880 170548 75886
rect 170496 75822 170548 75828
rect 170324 71746 170444 71774
rect 170324 69698 170352 71746
rect 170312 69692 170364 69698
rect 170312 69634 170364 69640
rect 170220 69012 170272 69018
rect 170220 68954 170272 68960
rect 170128 32428 170180 32434
rect 170128 32370 170180 32376
rect 170692 25702 170720 75890
rect 170784 75138 170812 79766
rect 170864 79756 170916 79762
rect 170864 79698 170916 79704
rect 171060 79750 171134 79778
rect 171244 79750 171318 79778
rect 170876 75857 170904 79698
rect 171060 79665 171088 79750
rect 171140 79688 171192 79694
rect 171046 79656 171102 79665
rect 170956 79620 171008 79626
rect 171140 79630 171192 79636
rect 171046 79591 171102 79600
rect 170956 79562 171008 79568
rect 170968 78713 170996 79562
rect 171152 78849 171180 79630
rect 171244 79422 171272 79750
rect 171382 79694 171410 80036
rect 171474 79744 171502 80036
rect 171566 79937 171594 80036
rect 171552 79928 171608 79937
rect 171552 79863 171608 79872
rect 171658 79778 171686 80036
rect 171750 79937 171778 80036
rect 171736 79928 171792 79937
rect 171842 79898 171870 80036
rect 171934 79937 171962 80036
rect 172026 79966 172054 80036
rect 172014 79960 172066 79966
rect 171920 79928 171976 79937
rect 171736 79863 171792 79872
rect 171830 79892 171882 79898
rect 172014 79902 172066 79908
rect 171920 79863 171976 79872
rect 171830 79834 171882 79840
rect 171968 79824 172020 79830
rect 171658 79750 171824 79778
rect 171968 79766 172020 79772
rect 171474 79716 171548 79744
rect 171370 79688 171422 79694
rect 171370 79630 171422 79636
rect 171232 79416 171284 79422
rect 171232 79358 171284 79364
rect 171520 79354 171548 79716
rect 171600 79688 171652 79694
rect 171600 79630 171652 79636
rect 171508 79348 171560 79354
rect 171508 79290 171560 79296
rect 171138 78840 171194 78849
rect 171138 78775 171194 78784
rect 170954 78704 171010 78713
rect 170954 78639 171010 78648
rect 171508 78600 171560 78606
rect 171508 78542 171560 78548
rect 171322 78296 171378 78305
rect 171322 78231 171378 78240
rect 171138 78160 171194 78169
rect 171138 78095 171194 78104
rect 171152 77489 171180 78095
rect 171336 77625 171364 78231
rect 171520 77897 171548 78542
rect 171612 78198 171640 79630
rect 171796 78674 171824 79750
rect 171876 79756 171928 79762
rect 171876 79698 171928 79704
rect 171888 79490 171916 79698
rect 171876 79484 171928 79490
rect 171876 79426 171928 79432
rect 171692 78668 171744 78674
rect 171692 78610 171744 78616
rect 171784 78668 171836 78674
rect 171784 78610 171836 78616
rect 171600 78192 171652 78198
rect 171600 78134 171652 78140
rect 171506 77888 171562 77897
rect 171506 77823 171562 77832
rect 171416 77648 171468 77654
rect 171322 77616 171378 77625
rect 171416 77590 171468 77596
rect 171322 77551 171378 77560
rect 171138 77480 171194 77489
rect 171138 77415 171194 77424
rect 170862 75848 170918 75857
rect 170862 75783 170918 75792
rect 170772 75132 170824 75138
rect 170772 75074 170824 75080
rect 171428 70394 171456 77590
rect 171428 70366 171640 70394
rect 171612 43450 171640 70366
rect 171704 69902 171732 78610
rect 171876 78396 171928 78402
rect 171876 78338 171928 78344
rect 171888 75914 171916 78338
rect 171980 77840 172008 79766
rect 172118 79744 172146 80036
rect 172072 79716 172146 79744
rect 172210 79744 172238 80036
rect 172302 79966 172330 80036
rect 172290 79960 172342 79966
rect 172394 79937 172422 80036
rect 172290 79902 172342 79908
rect 172380 79928 172436 79937
rect 172380 79863 172436 79872
rect 172486 79744 172514 80036
rect 172578 79937 172606 80036
rect 172564 79928 172620 79937
rect 172564 79863 172620 79872
rect 172210 79716 172284 79744
rect 172072 78441 172100 79716
rect 172058 78432 172114 78441
rect 172058 78367 172114 78376
rect 172256 78169 172284 79716
rect 172348 79716 172514 79744
rect 172348 78606 172376 79716
rect 172670 79676 172698 80036
rect 172624 79648 172698 79676
rect 172762 79676 172790 80036
rect 172854 79778 172882 80036
rect 172946 79966 172974 80036
rect 172934 79960 172986 79966
rect 172934 79902 172986 79908
rect 172854 79750 172928 79778
rect 172762 79648 172836 79676
rect 172336 78600 172388 78606
rect 172336 78542 172388 78548
rect 172242 78160 172298 78169
rect 172242 78095 172298 78104
rect 171980 77812 172100 77840
rect 171966 77752 172022 77761
rect 171966 77687 172022 77696
rect 171796 75886 171916 75914
rect 171692 69896 171744 69902
rect 171692 69838 171744 69844
rect 171692 69012 171744 69018
rect 171692 68954 171744 68960
rect 171600 43444 171652 43450
rect 171600 43386 171652 43392
rect 171704 33114 171732 68954
rect 171692 33108 171744 33114
rect 171692 33050 171744 33056
rect 170680 25696 170732 25702
rect 170680 25638 170732 25644
rect 170036 25560 170088 25566
rect 170036 25502 170088 25508
rect 169944 8968 169996 8974
rect 169944 8910 169996 8916
rect 169852 6180 169904 6186
rect 169852 6122 169904 6128
rect 169576 5228 169628 5234
rect 169576 5170 169628 5176
rect 164884 4820 164936 4826
rect 164884 4762 164936 4768
rect 165712 4820 165764 4826
rect 165712 4762 165764 4768
rect 163964 3732 164016 3738
rect 163964 3674 164016 3680
rect 162872 3454 163728 3482
rect 163700 480 163728 3454
rect 164896 480 164924 4762
rect 168380 3800 168432 3806
rect 168380 3742 168432 3748
rect 167184 3596 167236 3602
rect 167184 3538 167236 3544
rect 166080 3528 166132 3534
rect 166080 3470 166132 3476
rect 166092 480 166120 3470
rect 167196 480 167224 3538
rect 168392 480 168420 3742
rect 169588 480 169616 5170
rect 171796 3602 171824 75886
rect 171876 72412 171928 72418
rect 171876 72354 171928 72360
rect 171888 3670 171916 72354
rect 171980 17474 172008 77687
rect 172072 77586 172100 77812
rect 172428 77716 172480 77722
rect 172428 77658 172480 77664
rect 172150 77616 172206 77625
rect 172060 77580 172112 77586
rect 172150 77551 172206 77560
rect 172060 77522 172112 77528
rect 172060 76288 172112 76294
rect 172060 76230 172112 76236
rect 171968 17468 172020 17474
rect 171968 17410 172020 17416
rect 171968 5024 172020 5030
rect 171968 4966 172020 4972
rect 171876 3664 171928 3670
rect 171876 3606 171928 3612
rect 171784 3596 171836 3602
rect 171784 3538 171836 3544
rect 170772 3460 170824 3466
rect 170772 3402 170824 3408
rect 170784 480 170812 3402
rect 171980 480 172008 4966
rect 172072 3942 172100 76230
rect 172164 37942 172192 77551
rect 172334 77480 172390 77489
rect 172334 77415 172390 77424
rect 172244 76356 172296 76362
rect 172244 76298 172296 76304
rect 172152 37936 172204 37942
rect 172152 37878 172204 37884
rect 172060 3936 172112 3942
rect 172060 3878 172112 3884
rect 172256 3874 172284 76298
rect 172348 39370 172376 77415
rect 172440 40730 172468 77658
rect 172624 77178 172652 79648
rect 172612 77172 172664 77178
rect 172612 77114 172664 77120
rect 172808 76430 172836 79648
rect 172900 76498 172928 79750
rect 173038 79744 173066 80036
rect 172992 79716 173066 79744
rect 172992 79529 173020 79716
rect 173130 79676 173158 80036
rect 173222 79801 173250 80036
rect 173208 79792 173264 79801
rect 173314 79778 173342 80036
rect 173406 79898 173434 80036
rect 173498 79966 173526 80036
rect 173486 79960 173538 79966
rect 173486 79902 173538 79908
rect 173394 79892 173446 79898
rect 173394 79834 173446 79840
rect 173590 79812 173618 80036
rect 173498 79784 173618 79812
rect 173314 79750 173388 79778
rect 173208 79727 173264 79736
rect 173256 79688 173308 79694
rect 173130 79648 173204 79676
rect 172978 79520 173034 79529
rect 172978 79455 173034 79464
rect 173072 79484 173124 79490
rect 173072 79426 173124 79432
rect 173084 78985 173112 79426
rect 173070 78976 173126 78985
rect 173070 78911 173126 78920
rect 173176 78849 173204 79648
rect 173256 79630 173308 79636
rect 173268 79393 173296 79630
rect 173360 79529 173388 79750
rect 173498 79540 173526 79784
rect 173682 79778 173710 80036
rect 173774 79898 173802 80036
rect 173866 79966 173894 80036
rect 173958 79966 173986 80036
rect 174050 79966 174078 80036
rect 174142 79966 174170 80036
rect 173854 79960 173906 79966
rect 173854 79902 173906 79908
rect 173946 79960 173998 79966
rect 173946 79902 173998 79908
rect 174038 79960 174090 79966
rect 174038 79902 174090 79908
rect 174130 79960 174182 79966
rect 174130 79902 174182 79908
rect 174234 79914 174262 80036
rect 173762 79892 173814 79898
rect 174234 79886 174400 79914
rect 173762 79834 173814 79840
rect 173900 79824 173952 79830
rect 173682 79750 173756 79778
rect 173900 79766 173952 79772
rect 173992 79824 174044 79830
rect 173992 79766 174044 79772
rect 174176 79824 174228 79830
rect 174176 79766 174228 79772
rect 173624 79688 173676 79694
rect 173622 79656 173624 79665
rect 173676 79656 173678 79665
rect 173622 79591 173678 79600
rect 173346 79520 173402 79529
rect 173346 79455 173402 79464
rect 173452 79512 173526 79540
rect 173254 79384 173310 79393
rect 173254 79319 173310 79328
rect 173452 79121 173480 79512
rect 173438 79112 173494 79121
rect 173438 79047 173494 79056
rect 173728 78878 173756 79750
rect 173808 79756 173860 79762
rect 173808 79698 173860 79704
rect 173716 78872 173768 78878
rect 173162 78840 173218 78849
rect 173716 78814 173768 78820
rect 173162 78775 173218 78784
rect 173820 78470 173848 79698
rect 173912 79218 173940 79766
rect 174004 79257 174032 79766
rect 174188 79558 174216 79766
rect 174176 79552 174228 79558
rect 174176 79494 174228 79500
rect 173990 79248 174046 79257
rect 173900 79212 173952 79218
rect 173990 79183 174046 79192
rect 173900 79154 173952 79160
rect 173808 78464 173860 78470
rect 173808 78406 173860 78412
rect 173992 78396 174044 78402
rect 173992 78338 174044 78344
rect 173164 77308 173216 77314
rect 173164 77250 173216 77256
rect 172888 76492 172940 76498
rect 172888 76434 172940 76440
rect 172796 76424 172848 76430
rect 172796 76366 172848 76372
rect 172518 60072 172574 60081
rect 172518 60007 172574 60016
rect 172428 40724 172480 40730
rect 172428 40666 172480 40672
rect 172336 39364 172388 39370
rect 172336 39306 172388 39312
rect 172532 16574 172560 60007
rect 172532 16546 172744 16574
rect 172244 3868 172296 3874
rect 172244 3810 172296 3816
rect 134126 354 134238 480
rect 133892 326 134238 354
rect 134126 -960 134238 326
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 172716 354 172744 16546
rect 173176 3534 173204 77250
rect 173254 77208 173310 77217
rect 173254 77143 173310 77152
rect 173164 3528 173216 3534
rect 173164 3470 173216 3476
rect 173268 3330 173296 77143
rect 173898 75712 173954 75721
rect 173898 75647 173954 75656
rect 173348 74520 173400 74526
rect 173348 74462 173400 74468
rect 173360 3466 173388 74462
rect 173348 3460 173400 3466
rect 173348 3402 173400 3408
rect 173256 3324 173308 3330
rect 173256 3266 173308 3272
rect 173134 354 173246 480
rect 172716 326 173246 354
rect 173912 354 173940 75647
rect 174004 23322 174032 78338
rect 174372 71774 174400 79886
rect 174464 77654 174492 80242
rect 174556 78402 174584 80430
rect 174740 79626 174768 80446
rect 174832 80034 174860 80650
rect 174820 80028 174872 80034
rect 174820 79970 174872 79976
rect 174728 79620 174780 79626
rect 174728 79562 174780 79568
rect 174924 79354 174952 80650
rect 175924 80640 175976 80646
rect 175924 80582 175976 80588
rect 175096 80436 175148 80442
rect 175096 80378 175148 80384
rect 175108 79801 175136 80378
rect 175740 80164 175792 80170
rect 175740 80106 175792 80112
rect 175094 79792 175150 79801
rect 175094 79727 175150 79736
rect 174912 79348 174964 79354
rect 174912 79290 174964 79296
rect 174544 78396 174596 78402
rect 174544 78338 174596 78344
rect 174544 77784 174596 77790
rect 174544 77726 174596 77732
rect 174452 77648 174504 77654
rect 174452 77590 174504 77596
rect 174188 71746 174400 71774
rect 174188 70394 174216 71746
rect 174096 70366 174216 70394
rect 174096 45558 174124 70366
rect 174084 45552 174136 45558
rect 174084 45494 174136 45500
rect 173992 23316 174044 23322
rect 173992 23258 174044 23264
rect 174556 15978 174584 77726
rect 175752 77246 175780 80106
rect 175936 80102 175964 80582
rect 177028 80164 177080 80170
rect 177028 80106 177080 80112
rect 175924 80096 175976 80102
rect 175924 80038 175976 80044
rect 176658 79928 176714 79937
rect 176658 79863 176714 79872
rect 176672 78878 176700 79863
rect 176660 78872 176712 78878
rect 176566 78840 176622 78849
rect 176660 78814 176712 78820
rect 176566 78775 176622 78784
rect 176580 78606 176608 78775
rect 176568 78600 176620 78606
rect 176568 78542 176620 78548
rect 175924 77512 175976 77518
rect 175924 77454 175976 77460
rect 175740 77240 175792 77246
rect 175740 77182 175792 77188
rect 175278 69592 175334 69601
rect 175278 69527 175334 69536
rect 175292 16574 175320 69527
rect 175292 16546 175504 16574
rect 174544 15972 174596 15978
rect 174544 15914 174596 15920
rect 175476 480 175504 16546
rect 175936 6458 175964 77454
rect 177040 77450 177068 80106
rect 178512 80073 178540 80951
rect 178590 80880 178646 80889
rect 178590 80815 178646 80824
rect 178498 80064 178554 80073
rect 178498 79999 178554 80008
rect 178132 79280 178184 79286
rect 178132 79222 178184 79228
rect 177028 77444 177080 77450
rect 177028 77386 177080 77392
rect 177302 76120 177358 76129
rect 177302 76055 177358 76064
rect 176658 75576 176714 75585
rect 176658 75511 176714 75520
rect 176672 11694 176700 75511
rect 177316 73166 177344 76055
rect 177304 73160 177356 73166
rect 177304 73102 177356 73108
rect 178144 64874 178172 79222
rect 178604 78674 178632 80815
rect 178592 78668 178644 78674
rect 178592 78610 178644 78616
rect 178682 72720 178738 72729
rect 178682 72655 178738 72664
rect 178052 64846 178172 64874
rect 176752 27328 176804 27334
rect 176752 27270 176804 27276
rect 176660 11688 176712 11694
rect 176660 11630 176712 11636
rect 176764 6914 176792 27270
rect 178052 16574 178080 64846
rect 178052 16546 178632 16574
rect 177856 11688 177908 11694
rect 177856 11630 177908 11636
rect 176672 6886 176792 6914
rect 175924 6452 175976 6458
rect 175924 6394 175976 6400
rect 176672 480 176700 6886
rect 177868 480 177896 11630
rect 174238 354 174350 480
rect 173912 326 174350 354
rect 173134 -960 173246 326
rect 174238 -960 174350 326
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 178604 354 178632 16546
rect 178696 3806 178724 72655
rect 179616 71738 179644 135487
rect 180076 79354 180104 191830
rect 180156 151836 180208 151842
rect 180156 151778 180208 151784
rect 180168 81161 180196 151778
rect 180248 144900 180300 144906
rect 180248 144842 180300 144848
rect 180260 120086 180288 144842
rect 180340 140208 180392 140214
rect 180340 140150 180392 140156
rect 180352 128314 180380 140150
rect 180340 128308 180392 128314
rect 180340 128250 180392 128256
rect 180812 124137 180840 231066
rect 188344 205692 188396 205698
rect 188344 205634 188396 205640
rect 180892 162920 180944 162926
rect 180892 162862 180944 162868
rect 180904 133113 180932 162862
rect 182180 162172 182232 162178
rect 182180 162114 182232 162120
rect 181168 141772 181220 141778
rect 181168 141714 181220 141720
rect 181076 141364 181128 141370
rect 181076 141306 181128 141312
rect 180982 138680 181038 138689
rect 180982 138615 181038 138624
rect 180890 133104 180946 133113
rect 180890 133039 180946 133048
rect 180798 124128 180854 124137
rect 180798 124063 180854 124072
rect 180248 120080 180300 120086
rect 180248 120022 180300 120028
rect 180248 111852 180300 111858
rect 180248 111794 180300 111800
rect 180154 81152 180210 81161
rect 180154 81087 180210 81096
rect 180260 80442 180288 111794
rect 180340 99408 180392 99414
rect 180340 99350 180392 99356
rect 180352 81433 180380 99350
rect 180996 88330 181024 138615
rect 181088 115161 181116 141306
rect 181180 116657 181208 141714
rect 181258 137592 181314 137601
rect 181258 137527 181314 137536
rect 181166 116648 181222 116657
rect 181166 116583 181222 116592
rect 181074 115152 181130 115161
rect 181074 115087 181130 115096
rect 180984 88324 181036 88330
rect 180984 88266 181036 88272
rect 180996 88233 181024 88266
rect 180982 88224 181038 88233
rect 180982 88159 181038 88168
rect 180338 81424 180394 81433
rect 180338 81359 180394 81368
rect 180248 80436 180300 80442
rect 180248 80378 180300 80384
rect 180064 79348 180116 79354
rect 180064 79290 180116 79296
rect 180064 77920 180116 77926
rect 180064 77862 180116 77868
rect 179604 71732 179656 71738
rect 179604 71674 179656 71680
rect 179420 27260 179472 27266
rect 179420 27202 179472 27208
rect 179432 16574 179460 27202
rect 179432 16546 180012 16574
rect 178684 3800 178736 3806
rect 178684 3742 178736 3748
rect 179984 3482 180012 16546
rect 180076 5030 180104 77862
rect 180800 46232 180852 46238
rect 180800 46174 180852 46180
rect 180812 16574 180840 46174
rect 181272 33046 181300 137527
rect 182192 130121 182220 162114
rect 182272 144492 182324 144498
rect 182272 144434 182324 144440
rect 182178 130112 182234 130121
rect 182178 130047 182234 130056
rect 182284 128625 182312 144434
rect 182548 144424 182600 144430
rect 182548 144366 182600 144372
rect 182456 144356 182508 144362
rect 182456 144298 182508 144304
rect 182364 139528 182416 139534
rect 182364 139470 182416 139476
rect 182376 134609 182404 139470
rect 182362 134600 182418 134609
rect 182362 134535 182418 134544
rect 182364 134496 182416 134502
rect 182364 134438 182416 134444
rect 182270 128616 182326 128625
rect 182270 128551 182326 128560
rect 182180 128308 182232 128314
rect 182180 128250 182232 128256
rect 182192 112169 182220 128250
rect 182272 120080 182324 120086
rect 182272 120022 182324 120028
rect 182284 113665 182312 120022
rect 182376 118153 182404 134438
rect 182468 125633 182496 144298
rect 182560 127129 182588 144366
rect 182824 141704 182876 141710
rect 182824 141646 182876 141652
rect 182732 140140 182784 140146
rect 182732 140082 182784 140088
rect 182640 140072 182692 140078
rect 182640 140014 182692 140020
rect 182652 134502 182680 140014
rect 182640 134496 182692 134502
rect 182640 134438 182692 134444
rect 182744 134314 182772 140082
rect 182652 134286 182772 134314
rect 182546 127120 182602 127129
rect 182546 127055 182602 127064
rect 182454 125624 182510 125633
rect 182454 125559 182510 125568
rect 182652 121145 182680 134286
rect 182836 122834 182864 141646
rect 184204 125656 184256 125662
rect 184204 125598 184256 125604
rect 182744 122806 182864 122834
rect 182638 121136 182694 121145
rect 182638 121071 182694 121080
rect 182744 119649 182772 122806
rect 182730 119640 182786 119649
rect 182730 119575 182786 119584
rect 182362 118144 182418 118153
rect 182362 118079 182418 118088
rect 182270 113656 182326 113665
rect 182270 113591 182326 113600
rect 182178 112160 182234 112169
rect 182178 112095 182234 112104
rect 183284 111784 183336 111790
rect 183284 111726 183336 111732
rect 183296 110673 183324 111726
rect 183282 110664 183338 110673
rect 183282 110599 183338 110608
rect 183468 110424 183520 110430
rect 183468 110366 183520 110372
rect 183480 109177 183508 110366
rect 183466 109168 183522 109177
rect 183466 109103 183522 109112
rect 182272 108996 182324 109002
rect 182272 108938 182324 108944
rect 182284 107681 182312 108938
rect 182270 107672 182326 107681
rect 182270 107607 182326 107616
rect 183468 106276 183520 106282
rect 183468 106218 183520 106224
rect 183480 106185 183508 106218
rect 183466 106176 183522 106185
rect 183466 106111 183522 106120
rect 183468 104848 183520 104854
rect 183468 104790 183520 104796
rect 183480 104689 183508 104790
rect 183466 104680 183522 104689
rect 183466 104615 183522 104624
rect 183468 103488 183520 103494
rect 183468 103430 183520 103436
rect 183480 103193 183508 103430
rect 183466 103184 183522 103193
rect 183466 103119 183522 103128
rect 182916 102128 182968 102134
rect 182916 102070 182968 102076
rect 182928 101697 182956 102070
rect 182914 101688 182970 101697
rect 182914 101623 182970 101632
rect 182916 100700 182968 100706
rect 182916 100642 182968 100648
rect 182928 100201 182956 100642
rect 182914 100192 182970 100201
rect 182914 100127 182970 100136
rect 183100 99340 183152 99346
rect 183100 99282 183152 99288
rect 183112 98705 183140 99282
rect 183098 98696 183154 98705
rect 183098 98631 183154 98640
rect 183468 97980 183520 97986
rect 183468 97922 183520 97928
rect 183480 97209 183508 97922
rect 183466 97200 183522 97209
rect 183466 97135 183522 97144
rect 183192 96620 183244 96626
rect 183192 96562 183244 96568
rect 183204 95713 183232 96562
rect 183190 95704 183246 95713
rect 183190 95639 183246 95648
rect 183284 95192 183336 95198
rect 183284 95134 183336 95140
rect 183296 94217 183324 95134
rect 183282 94208 183338 94217
rect 183282 94143 183338 94152
rect 183284 93832 183336 93838
rect 183284 93774 183336 93780
rect 183296 92721 183324 93774
rect 183282 92712 183338 92721
rect 183282 92647 183338 92656
rect 183468 92472 183520 92478
rect 183468 92414 183520 92420
rect 183480 91225 183508 92414
rect 183466 91216 183522 91225
rect 183466 91151 183522 91160
rect 182178 89720 182234 89729
rect 182178 89655 182180 89664
rect 182232 89655 182234 89664
rect 182180 89626 182232 89632
rect 184216 86766 184244 125598
rect 188356 89690 188384 205634
rect 207032 198014 207060 230588
rect 236012 230574 236578 230602
rect 207020 198008 207072 198014
rect 207020 197950 207072 197956
rect 236012 196722 236040 230574
rect 266556 228410 266584 230588
rect 266544 228404 266596 228410
rect 266544 228346 266596 228352
rect 267004 228404 267056 228410
rect 267004 228346 267056 228352
rect 236000 196716 236052 196722
rect 236000 196658 236052 196664
rect 267016 195906 267044 228346
rect 296732 199442 296760 230588
rect 296720 199436 296772 199442
rect 296720 199378 296772 199384
rect 327092 196654 327120 230588
rect 356532 228410 356560 230588
rect 356520 228404 356572 228410
rect 356520 228346 356572 228352
rect 385040 220788 385092 220794
rect 385040 220730 385092 220736
rect 385052 217938 385080 220730
rect 386524 219434 386552 230588
rect 391216 227798 391244 232222
rect 393964 231872 394016 231878
rect 393964 231814 394016 231820
rect 388444 227792 388496 227798
rect 388444 227734 388496 227740
rect 391204 227792 391256 227798
rect 391204 227734 391256 227740
rect 391296 227792 391348 227798
rect 391296 227734 391348 227740
rect 386432 219406 386552 219434
rect 380900 217932 380952 217938
rect 380900 217874 380952 217880
rect 385040 217932 385092 217938
rect 385040 217874 385092 217880
rect 380912 215490 380940 217874
rect 375472 215484 375524 215490
rect 375472 215426 375524 215432
rect 380900 215484 380952 215490
rect 380900 215426 380952 215432
rect 375484 213994 375512 215426
rect 375472 213988 375524 213994
rect 375472 213930 375524 213936
rect 371884 213920 371936 213926
rect 371884 213862 371936 213868
rect 371896 205766 371924 213862
rect 370504 205760 370556 205766
rect 370504 205702 370556 205708
rect 371884 205760 371936 205766
rect 371884 205702 371936 205708
rect 327080 196648 327132 196654
rect 327080 196590 327132 196596
rect 267004 195900 267056 195906
rect 267004 195842 267056 195848
rect 366364 174548 366416 174554
rect 366364 174490 366416 174496
rect 226984 165640 227036 165646
rect 226984 165582 227036 165588
rect 188344 89684 188396 89690
rect 188344 89626 188396 89632
rect 226996 88330 227024 165582
rect 365536 136264 365588 136270
rect 365536 136206 365588 136212
rect 365548 133958 365576 136206
rect 362224 133952 362276 133958
rect 362224 133894 362276 133900
rect 365536 133952 365588 133958
rect 365536 133894 365588 133900
rect 355968 119400 356020 119406
rect 355968 119342 356020 119348
rect 355980 116890 356008 119342
rect 352564 116884 352616 116890
rect 352564 116826 352616 116832
rect 355968 116884 356020 116890
rect 355968 116826 356020 116832
rect 352576 110498 352604 116826
rect 362236 111790 362264 133894
rect 366376 119406 366404 174490
rect 370516 140826 370544 205702
rect 384396 205488 384448 205494
rect 384396 205430 384448 205436
rect 384408 203386 384436 205430
rect 385684 204264 385736 204270
rect 385684 204206 385736 204212
rect 382924 203380 382976 203386
rect 382924 203322 382976 203328
rect 384396 203380 384448 203386
rect 384396 203322 384448 203328
rect 382936 196926 382964 203322
rect 380900 196920 380952 196926
rect 380900 196862 380952 196868
rect 382924 196920 382976 196926
rect 382924 196862 382976 196868
rect 380164 193996 380216 194002
rect 380164 193938 380216 193944
rect 380176 174554 380204 193938
rect 380912 193866 380940 196862
rect 385696 194002 385724 204206
rect 386432 195974 386460 219406
rect 388456 205494 388484 227734
rect 391308 225010 391336 227734
rect 389088 225004 389140 225010
rect 389088 224946 389140 224952
rect 391296 225004 391348 225010
rect 391296 224946 391348 224952
rect 389100 220794 389128 224946
rect 389088 220788 389140 220794
rect 389088 220730 389140 220736
rect 391204 213172 391256 213178
rect 391204 213114 391256 213120
rect 388444 205488 388496 205494
rect 388444 205430 388496 205436
rect 391216 204270 391244 213114
rect 391204 204264 391256 204270
rect 391204 204206 391256 204212
rect 386420 195968 386472 195974
rect 386420 195910 386472 195916
rect 385684 193996 385736 194002
rect 385684 193938 385736 193944
rect 380900 193860 380952 193866
rect 380900 193802 380952 193808
rect 387064 189100 387116 189106
rect 387064 189042 387116 189048
rect 387076 174554 387104 189042
rect 380164 174548 380216 174554
rect 380164 174490 380216 174496
rect 385684 174548 385736 174554
rect 385684 174490 385736 174496
rect 387064 174548 387116 174554
rect 387064 174490 387116 174496
rect 385696 167142 385724 174490
rect 384304 167136 384356 167142
rect 384304 167078 384356 167084
rect 385684 167136 385736 167142
rect 385684 167078 385736 167084
rect 384316 165306 384344 167078
rect 380900 165300 380952 165306
rect 380900 165242 380952 165248
rect 384304 165300 384356 165306
rect 384304 165242 384356 165248
rect 380912 163130 380940 165242
rect 380256 163124 380308 163130
rect 380256 163066 380308 163072
rect 380900 163124 380952 163130
rect 380900 163066 380952 163072
rect 380268 157418 380296 163066
rect 378876 157412 378928 157418
rect 378876 157354 378928 157360
rect 380256 157412 380308 157418
rect 380256 157354 380308 157360
rect 378888 154154 378916 157354
rect 377404 154148 377456 154154
rect 377404 154090 377456 154096
rect 378876 154148 378928 154154
rect 378876 154090 378928 154096
rect 367376 140820 367428 140826
rect 367376 140762 367428 140768
rect 370504 140820 370556 140826
rect 370504 140762 370556 140768
rect 367388 136270 367416 140762
rect 377416 139874 377444 154090
rect 375012 139868 375064 139874
rect 375012 139810 375064 139816
rect 377404 139868 377456 139874
rect 377404 139810 377456 139816
rect 375024 137426 375052 139810
rect 373264 137420 373316 137426
rect 373264 137362 373316 137368
rect 375012 137420 375064 137426
rect 375012 137362 375064 137368
rect 367376 136264 367428 136270
rect 367376 136206 367428 136212
rect 373276 129810 373304 137362
rect 373264 129804 373316 129810
rect 373264 129746 373316 129752
rect 369860 129736 369912 129742
rect 369860 129678 369912 129684
rect 369872 127106 369900 129678
rect 369780 127078 369900 127106
rect 369780 125186 369808 127078
rect 367744 125180 367796 125186
rect 367744 125122 367796 125128
rect 369768 125180 369820 125186
rect 369768 125122 369820 125128
rect 366364 119400 366416 119406
rect 366364 119342 366416 119348
rect 362224 111784 362276 111790
rect 362224 111726 362276 111732
rect 349528 110492 349580 110498
rect 349528 110434 349580 110440
rect 352564 110492 352616 110498
rect 352564 110434 352616 110440
rect 349540 105602 349568 110434
rect 367756 110430 367784 125122
rect 367744 110424 367796 110430
rect 367744 110366 367796 110372
rect 346400 105596 346452 105602
rect 346400 105538 346452 105544
rect 349528 105596 349580 105602
rect 349528 105538 349580 105544
rect 346412 102202 346440 105538
rect 343640 102196 343692 102202
rect 343640 102138 343692 102144
rect 346400 102196 346452 102202
rect 346400 102138 346452 102144
rect 343652 94994 343680 102138
rect 339224 94988 339276 94994
rect 339224 94930 339276 94936
rect 343640 94988 343692 94994
rect 343640 94930 343692 94936
rect 339236 91798 339264 94930
rect 329104 91792 329156 91798
rect 329104 91734 329156 91740
rect 339224 91792 339276 91798
rect 339224 91734 339276 91740
rect 226984 88324 227036 88330
rect 226984 88266 227036 88272
rect 182180 86760 182232 86766
rect 182178 86728 182180 86737
rect 184204 86760 184256 86766
rect 182232 86728 182234 86737
rect 184204 86702 184256 86708
rect 182178 86663 182234 86672
rect 182640 85604 182692 85610
rect 182640 85546 182692 85552
rect 182652 85241 182680 85546
rect 182638 85232 182694 85241
rect 182638 85167 182694 85176
rect 182822 83736 182878 83745
rect 182822 83671 182878 83680
rect 182454 82240 182510 82249
rect 182454 82175 182510 82184
rect 182468 81462 182496 82175
rect 182456 81456 182508 81462
rect 182456 81398 182508 81404
rect 182180 80300 182232 80306
rect 182180 80242 182232 80248
rect 181260 33040 181312 33046
rect 181260 32982 181312 32988
rect 180812 16546 181024 16574
rect 180064 5024 180116 5030
rect 180064 4966 180116 4972
rect 179984 3454 180288 3482
rect 180260 480 180288 3454
rect 179022 354 179134 480
rect 178604 326 179134 354
rect 179022 -960 179134 326
rect 180218 -960 180330 480
rect 180996 354 181024 16546
rect 181414 354 181526 480
rect 180996 326 181526 354
rect 182192 354 182220 80242
rect 182836 46918 182864 83671
rect 200120 80232 200172 80238
rect 200120 80174 200172 80180
rect 195980 79144 196032 79150
rect 195980 79086 196032 79092
rect 194598 74080 194654 74089
rect 194598 74015 194654 74024
rect 184940 68672 184992 68678
rect 184940 68614 184992 68620
rect 182824 46912 182876 46918
rect 182824 46854 182876 46860
rect 183560 27192 183612 27198
rect 183560 27134 183612 27140
rect 183572 16574 183600 27134
rect 183572 16546 183784 16574
rect 183756 480 183784 16546
rect 184952 11694 184980 68614
rect 189080 67448 189132 67454
rect 189080 67390 189132 67396
rect 185032 61532 185084 61538
rect 185032 61474 185084 61480
rect 184940 11688 184992 11694
rect 184940 11630 184992 11636
rect 185044 6914 185072 61474
rect 187700 34128 187752 34134
rect 187700 34070 187752 34076
rect 186320 28484 186372 28490
rect 186320 28426 186372 28432
rect 186332 16574 186360 28426
rect 187712 16574 187740 34070
rect 189092 16574 189120 67390
rect 193218 65512 193274 65521
rect 193218 65447 193274 65456
rect 190460 28552 190512 28558
rect 190460 28494 190512 28500
rect 186332 16546 186912 16574
rect 187712 16546 188568 16574
rect 189092 16546 189304 16574
rect 186136 11688 186188 11694
rect 186136 11630 186188 11636
rect 184952 6886 185072 6914
rect 184952 480 184980 6886
rect 186148 480 186176 11630
rect 182518 354 182630 480
rect 182192 326 182630 354
rect 181414 -960 181526 326
rect 182518 -960 182630 326
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 186884 354 186912 16546
rect 188540 480 188568 16546
rect 187302 354 187414 480
rect 186884 326 187414 354
rect 187302 -960 187414 326
rect 188498 -960 188610 480
rect 189276 354 189304 16546
rect 189694 354 189806 480
rect 189276 326 189806 354
rect 190472 354 190500 28494
rect 191838 19000 191894 19009
rect 191838 18935 191894 18944
rect 191852 16574 191880 18935
rect 191852 16546 192064 16574
rect 192036 480 192064 16546
rect 193232 480 193260 65447
rect 193310 28520 193366 28529
rect 193310 28455 193366 28464
rect 193324 16574 193352 28455
rect 194612 16574 194640 74015
rect 195992 16574 196020 79086
rect 197360 77104 197412 77110
rect 197360 77046 197412 77052
rect 197372 16574 197400 77046
rect 198740 34060 198792 34066
rect 198740 34002 198792 34008
rect 193324 16546 194456 16574
rect 194612 16546 195192 16574
rect 195992 16546 196848 16574
rect 197372 16546 197952 16574
rect 194428 480 194456 16546
rect 190798 354 190910 480
rect 190472 326 190910 354
rect 189694 -960 189806 326
rect 190798 -960 190910 326
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195164 354 195192 16546
rect 196820 480 196848 16546
rect 197924 480 197952 16546
rect 195582 354 195694 480
rect 195164 326 195694 354
rect 195582 -960 195694 326
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198752 354 198780 34002
rect 200132 16574 200160 80174
rect 231860 80164 231912 80170
rect 231860 80106 231912 80112
rect 213920 79008 213972 79014
rect 213920 78950 213972 78956
rect 211804 77036 211856 77042
rect 211804 76978 211856 76984
rect 209780 74248 209832 74254
rect 209780 74190 209832 74196
rect 202880 65952 202932 65958
rect 202880 65894 202932 65900
rect 201500 33992 201552 33998
rect 201500 33934 201552 33940
rect 200132 16546 200344 16574
rect 200316 480 200344 16546
rect 201512 11694 201540 33934
rect 201592 28416 201644 28422
rect 201592 28358 201644 28364
rect 201500 11688 201552 11694
rect 201500 11630 201552 11636
rect 201604 6914 201632 28358
rect 202892 16574 202920 65894
rect 207020 65884 207072 65890
rect 207020 65826 207072 65832
rect 205640 33924 205692 33930
rect 205640 33866 205692 33872
rect 204260 30116 204312 30122
rect 204260 30058 204312 30064
rect 204272 16574 204300 30058
rect 205652 16574 205680 33866
rect 202892 16546 203472 16574
rect 204272 16546 205128 16574
rect 205652 16546 206232 16574
rect 202696 11688 202748 11694
rect 202696 11630 202748 11636
rect 201512 6886 201632 6914
rect 201512 480 201540 6886
rect 202708 480 202736 11630
rect 199078 354 199190 480
rect 198752 326 199190 354
rect 199078 -960 199190 326
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203444 354 203472 16546
rect 205100 480 205128 16546
rect 206204 480 206232 16546
rect 203862 354 203974 480
rect 203444 326 203974 354
rect 203862 -960 203974 326
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207032 354 207060 65826
rect 208400 30048 208452 30054
rect 208400 29990 208452 29996
rect 208412 16574 208440 29990
rect 208412 16546 208624 16574
rect 208596 480 208624 16546
rect 209792 480 209820 74190
rect 209872 70100 209924 70106
rect 209872 70042 209924 70048
rect 209884 16574 209912 70042
rect 209884 16546 211016 16574
rect 210988 480 211016 16546
rect 211816 3262 211844 76978
rect 213932 16574 213960 78950
rect 226340 76968 226392 76974
rect 226340 76910 226392 76916
rect 216680 74180 216732 74186
rect 216680 74122 216732 74128
rect 215300 24608 215352 24614
rect 215300 24550 215352 24556
rect 213932 16546 214512 16574
rect 213366 10704 213422 10713
rect 213366 10639 213422 10648
rect 212172 3324 212224 3330
rect 212172 3266 212224 3272
rect 211804 3256 211856 3262
rect 211804 3198 211856 3204
rect 212184 480 212212 3266
rect 213380 480 213408 10639
rect 214484 480 214512 16546
rect 207358 354 207470 480
rect 207032 326 207470 354
rect 207358 -960 207470 326
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215312 354 215340 24550
rect 216692 16574 216720 74122
rect 223580 74112 223632 74118
rect 223580 74054 223632 74060
rect 218060 68604 218112 68610
rect 218060 68546 218112 68552
rect 216692 16546 216904 16574
rect 216876 480 216904 16546
rect 218072 480 218100 68546
rect 220820 65816 220872 65822
rect 220820 65758 220872 65764
rect 218152 24540 218204 24546
rect 218152 24482 218204 24488
rect 218164 16574 218192 24482
rect 220832 16574 220860 65758
rect 222200 26036 222252 26042
rect 222200 25978 222252 25984
rect 222212 16574 222240 25978
rect 218164 16546 219296 16574
rect 220832 16546 221136 16574
rect 222212 16546 222792 16574
rect 219268 480 219296 16546
rect 220452 5160 220504 5166
rect 220452 5102 220504 5108
rect 220464 480 220492 5102
rect 215638 354 215750 480
rect 215312 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221108 354 221136 16546
rect 222764 480 222792 16546
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223592 354 223620 74054
rect 225144 7948 225196 7954
rect 225144 7890 225196 7896
rect 225156 480 225184 7890
rect 226352 480 226380 76910
rect 230478 73944 230534 73953
rect 230478 73879 230534 73888
rect 227718 59936 227774 59945
rect 227718 59871 227774 59880
rect 226430 34096 226486 34105
rect 226430 34031 226486 34040
rect 226444 16574 226472 34031
rect 227732 16574 227760 59871
rect 229098 28384 229154 28393
rect 229098 28319 229154 28328
rect 229112 16574 229140 28319
rect 230492 16574 230520 73879
rect 226444 16546 227576 16574
rect 227732 16546 228312 16574
rect 229112 16546 229416 16574
rect 230492 16546 231072 16574
rect 227548 480 227576 16546
rect 223918 354 224030 480
rect 223592 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228284 354 228312 16546
rect 228702 354 228814 480
rect 228284 326 228814 354
rect 229388 354 229416 16546
rect 231044 480 231072 16546
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 228702 -960 228814 326
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 231872 354 231900 80106
rect 252560 80096 252612 80102
rect 252560 80038 252612 80044
rect 249800 79076 249852 79082
rect 249800 79018 249852 79024
rect 247684 78328 247736 78334
rect 247684 78270 247736 78276
rect 247038 76936 247094 76945
rect 240140 76900 240192 76906
rect 247038 76871 247094 76880
rect 240140 76842 240192 76848
rect 234620 64524 234672 64530
rect 234620 64466 234672 64472
rect 233240 29980 233292 29986
rect 233240 29922 233292 29928
rect 233252 16574 233280 29922
rect 233252 16546 233464 16574
rect 233436 480 233464 16546
rect 234632 11694 234660 64466
rect 238760 64456 238812 64462
rect 238760 64398 238812 64404
rect 234712 33856 234764 33862
rect 234712 33798 234764 33804
rect 234620 11688 234672 11694
rect 234620 11630 234672 11636
rect 234724 6914 234752 33798
rect 236000 29912 236052 29918
rect 236000 29854 236052 29860
rect 236012 16574 236040 29854
rect 238772 16574 238800 64398
rect 236012 16546 236592 16574
rect 238772 16546 239352 16574
rect 235816 11688 235868 11694
rect 235816 11630 235868 11636
rect 234632 6886 234752 6914
rect 234632 480 234660 6886
rect 235828 480 235856 11630
rect 232198 354 232310 480
rect 231872 326 232310 354
rect 232198 -960 232310 326
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 16546
rect 237656 12028 237708 12034
rect 237656 11970 237708 11976
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 237668 354 237696 11970
rect 239324 480 239352 16546
rect 238086 354 238198 480
rect 237668 326 238198 354
rect 236982 -960 237094 326
rect 238086 -960 238198 326
rect 239282 -960 239394 480
rect 240152 354 240180 76842
rect 244278 73808 244334 73817
rect 244278 73743 244334 73752
rect 242900 31476 242952 31482
rect 242900 31418 242952 31424
rect 241704 14816 241756 14822
rect 241704 14758 241756 14764
rect 241716 480 241744 14758
rect 242912 4214 242940 31418
rect 244292 16574 244320 73743
rect 247052 16574 247080 76871
rect 247696 20194 247724 78270
rect 248418 20224 248474 20233
rect 247684 20188 247736 20194
rect 248418 20159 248474 20168
rect 247684 20130 247736 20136
rect 244292 16546 245240 16574
rect 247052 16546 247632 16574
rect 242992 7880 243044 7886
rect 242992 7822 243044 7828
rect 242900 4208 242952 4214
rect 242900 4150 242952 4156
rect 243004 3482 243032 7822
rect 244096 4208 244148 4214
rect 244096 4150 244148 4156
rect 242912 3454 243032 3482
rect 242912 480 242940 3454
rect 244108 480 244136 4150
rect 245212 480 245240 16546
rect 246394 7712 246450 7721
rect 246394 7647 246450 7656
rect 246408 480 246436 7647
rect 247604 480 247632 16546
rect 240478 354 240590 480
rect 240152 326 240590 354
rect 240478 -960 240590 326
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248432 354 248460 20159
rect 249812 16574 249840 79018
rect 251180 74044 251232 74050
rect 251180 73986 251232 73992
rect 249812 16546 250024 16574
rect 249996 480 250024 16546
rect 251192 4214 251220 73986
rect 251272 65748 251324 65754
rect 251272 65690 251324 65696
rect 251180 4208 251232 4214
rect 251180 4150 251232 4156
rect 251284 3482 251312 65690
rect 252572 16574 252600 80038
rect 267740 78940 267792 78946
rect 267740 78882 267792 78888
rect 253204 78260 253256 78266
rect 253204 78202 253256 78208
rect 253216 20126 253244 78202
rect 260840 76832 260892 76838
rect 260840 76774 260892 76780
rect 256700 65680 256752 65686
rect 256700 65622 256752 65628
rect 253940 29844 253992 29850
rect 253940 29786 253992 29792
rect 253204 20120 253256 20126
rect 253204 20062 253256 20068
rect 253952 16574 253980 29786
rect 255320 20392 255372 20398
rect 255320 20334 255372 20340
rect 255332 16574 255360 20334
rect 252572 16546 253520 16574
rect 253952 16546 254256 16574
rect 255332 16546 255912 16574
rect 252376 4208 252428 4214
rect 252376 4150 252428 4156
rect 251192 3454 251312 3482
rect 251192 480 251220 3454
rect 252388 480 252416 4150
rect 253492 480 253520 16546
rect 248758 354 248870 480
rect 248432 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254228 354 254256 16546
rect 255884 480 255912 16546
rect 254646 354 254758 480
rect 254228 326 254758 354
rect 254646 -960 254758 326
rect 255842 -960 255954 480
rect 256712 354 256740 65622
rect 259460 35624 259512 35630
rect 259460 35566 259512 35572
rect 258080 29776 258132 29782
rect 258080 29718 258132 29724
rect 258092 16574 258120 29718
rect 258092 16546 258304 16574
rect 258276 480 258304 16546
rect 259472 480 259500 35566
rect 260852 16574 260880 76774
rect 266358 33960 266414 33969
rect 266358 33895 266414 33904
rect 262220 20324 262272 20330
rect 262220 20266 262272 20272
rect 262232 16574 262260 20266
rect 266372 16574 266400 33895
rect 260852 16546 261800 16574
rect 262232 16546 262536 16574
rect 266372 16546 266584 16574
rect 260656 9308 260708 9314
rect 260656 9250 260708 9256
rect 260668 480 260696 9250
rect 261772 480 261800 16546
rect 257038 354 257150 480
rect 256712 326 257150 354
rect 257038 -960 257150 326
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 354 262536 16546
rect 264150 9208 264206 9217
rect 264150 9143 264206 9152
rect 264164 480 264192 9143
rect 265346 7576 265402 7585
rect 265346 7511 265402 7520
rect 265360 480 265388 7511
rect 266556 480 266584 16546
rect 267752 480 267780 78882
rect 329116 78878 329144 91734
rect 393976 80646 394004 231814
rect 395356 223582 395384 232290
rect 395448 227798 395476 232358
rect 396460 232354 396488 673202
rect 396724 430636 396776 430642
rect 396724 430578 396776 430584
rect 396540 240100 396592 240106
rect 396540 240042 396592 240048
rect 396552 238814 396580 240042
rect 396540 238808 396592 238814
rect 396540 238750 396592 238756
rect 396632 238740 396684 238746
rect 396632 238682 396684 238688
rect 396540 238672 396592 238678
rect 396540 238614 396592 238620
rect 396448 232348 396500 232354
rect 396448 232290 396500 232296
rect 396552 232286 396580 238614
rect 396644 232422 396672 238682
rect 396632 232416 396684 232422
rect 396632 232358 396684 232364
rect 396540 232280 396592 232286
rect 396540 232222 396592 232228
rect 395436 227792 395488 227798
rect 395436 227734 395488 227740
rect 394056 223576 394108 223582
rect 394056 223518 394108 223524
rect 395344 223576 395396 223582
rect 395344 223518 395396 223524
rect 394068 189106 394096 223518
rect 394424 218136 394476 218142
rect 394424 218078 394476 218084
rect 394436 213178 394464 218078
rect 394424 213172 394476 213178
rect 394424 213114 394476 213120
rect 394056 189100 394108 189106
rect 394056 189042 394108 189048
rect 396736 81025 396764 430578
rect 396908 378208 396960 378214
rect 396908 378150 396960 378156
rect 396816 271924 396868 271930
rect 396816 271866 396868 271872
rect 396722 81016 396778 81025
rect 396722 80951 396778 80960
rect 396828 80782 396856 271866
rect 396920 80889 396948 378150
rect 397092 324352 397144 324358
rect 397092 324294 397144 324300
rect 396906 80880 396962 80889
rect 396906 80815 396962 80824
rect 396816 80776 396868 80782
rect 397104 80753 397132 324294
rect 396816 80718 396868 80724
rect 397090 80744 397146 80753
rect 397090 80679 397146 80688
rect 393964 80640 394016 80646
rect 393964 80582 394016 80588
rect 329104 78872 329156 78878
rect 397472 78849 397500 703520
rect 410524 700460 410576 700466
rect 410524 700402 410576 700408
rect 409144 700392 409196 700398
rect 409144 700334 409196 700340
rect 407764 700324 407816 700330
rect 407764 700266 407816 700272
rect 406384 670744 406436 670750
rect 406384 670686 406436 670692
rect 405004 616888 405056 616894
rect 405004 616830 405056 616836
rect 403624 563100 403676 563106
rect 403624 563042 403676 563048
rect 400864 510672 400916 510678
rect 400864 510614 400916 510620
rect 399484 456816 399536 456822
rect 399484 456758 399536 456764
rect 398104 418192 398156 418198
rect 398104 418134 398156 418140
rect 397552 343664 397604 343670
rect 397552 343606 397604 343612
rect 397564 218142 397592 343606
rect 397552 218136 397604 218142
rect 397552 218078 397604 218084
rect 398116 144294 398144 418134
rect 398196 311908 398248 311914
rect 398196 311850 398248 311856
rect 398104 144288 398156 144294
rect 398104 144230 398156 144236
rect 398208 142934 398236 311850
rect 398196 142928 398248 142934
rect 398196 142870 398248 142876
rect 399496 97986 399524 456758
rect 400876 99346 400904 510614
rect 403636 100706 403664 563042
rect 405016 102134 405044 616830
rect 406396 103494 406424 670686
rect 407776 104854 407804 700266
rect 409156 106282 409184 700334
rect 410536 109002 410564 700402
rect 412652 141642 412680 703582
rect 413480 703474 413508 703582
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 413664 703474 413692 703520
rect 413480 703446 413692 703474
rect 429856 700466 429884 703520
rect 429844 700460 429896 700466
rect 429844 700402 429896 700408
rect 421564 404388 421616 404394
rect 421564 404330 421616 404336
rect 418804 351960 418856 351966
rect 418804 351902 418856 351908
rect 417424 298172 417476 298178
rect 417424 298114 417476 298120
rect 414664 244316 414716 244322
rect 414664 244258 414716 244264
rect 412640 141636 412692 141642
rect 412640 141578 412692 141584
rect 410524 108996 410576 109002
rect 410524 108938 410576 108944
rect 409144 106276 409196 106282
rect 409144 106218 409196 106224
rect 407764 104848 407816 104854
rect 407764 104790 407816 104796
rect 406384 103488 406436 103494
rect 406384 103430 406436 103436
rect 405004 102128 405056 102134
rect 405004 102070 405056 102076
rect 403624 100700 403676 100706
rect 403624 100642 403676 100648
rect 400864 99340 400916 99346
rect 400864 99282 400916 99288
rect 399484 97980 399536 97986
rect 399484 97922 399536 97928
rect 414676 92478 414704 244258
rect 417436 93838 417464 298114
rect 418816 95198 418844 351902
rect 418896 258120 418948 258126
rect 418896 258062 418948 258068
rect 418908 142866 418936 258062
rect 418896 142860 418948 142866
rect 418896 142802 418948 142808
rect 421576 96626 421604 404330
rect 421564 96620 421616 96626
rect 421564 96562 421616 96568
rect 418804 95192 418856 95198
rect 418804 95134 418856 95140
rect 417424 93832 417476 93838
rect 417424 93774 417476 93780
rect 414664 92472 414716 92478
rect 414664 92414 414716 92420
rect 430578 80200 430634 80209
rect 430578 80135 430634 80144
rect 329104 78814 329156 78820
rect 397458 78840 397514 78849
rect 397458 78775 397514 78784
rect 322204 78192 322256 78198
rect 322204 78134 322256 78140
rect 282918 76800 282974 76809
rect 282918 76735 282974 76744
rect 288440 76764 288492 76770
rect 270500 67380 270552 67386
rect 270500 67322 270552 67328
rect 269120 33788 269172 33794
rect 269120 33730 269172 33736
rect 267832 31408 267884 31414
rect 267832 31350 267884 31356
rect 267844 16574 267872 31350
rect 269132 16574 269160 33730
rect 270512 16574 270540 67322
rect 274640 63164 274692 63170
rect 274640 63106 274692 63112
rect 271880 28348 271932 28354
rect 271880 28290 271932 28296
rect 271892 16574 271920 28290
rect 273260 20256 273312 20262
rect 273260 20198 273312 20204
rect 267844 16546 268424 16574
rect 269132 16546 270080 16574
rect 270512 16546 270816 16574
rect 271892 16546 272472 16574
rect 262926 354 263038 480
rect 262508 326 263038 354
rect 262926 -960 263038 326
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268396 354 268424 16546
rect 270052 480 270080 16546
rect 268814 354 268926 480
rect 268396 326 268926 354
rect 268814 -960 268926 326
rect 270010 -960 270122 480
rect 270788 354 270816 16546
rect 272444 480 272472 16546
rect 271206 354 271318 480
rect 270788 326 271318 354
rect 271206 -960 271318 326
rect 272402 -960 272514 480
rect 273272 354 273300 20198
rect 274652 16574 274680 63106
rect 280158 44840 280214 44849
rect 280158 44775 280214 44784
rect 276020 35556 276072 35562
rect 276020 35498 276072 35504
rect 274652 16546 274864 16574
rect 274836 480 274864 16546
rect 276032 4214 276060 35498
rect 276112 27124 276164 27130
rect 276112 27066 276164 27072
rect 276020 4208 276072 4214
rect 276020 4150 276072 4156
rect 276124 3482 276152 27066
rect 278780 25968 278832 25974
rect 278780 25910 278832 25916
rect 278792 16574 278820 25910
rect 280172 16574 280200 44775
rect 282932 16574 282960 76735
rect 288440 76706 288492 76712
rect 284298 72584 284354 72593
rect 284298 72519 284354 72528
rect 278792 16546 279096 16574
rect 280172 16546 280752 16574
rect 282932 16546 283144 16574
rect 278320 9240 278372 9246
rect 278320 9182 278372 9188
rect 276756 4208 276808 4214
rect 276756 4150 276808 4156
rect 276032 3454 276152 3482
rect 276032 480 276060 3454
rect 273598 354 273710 480
rect 273272 326 273710 354
rect 273598 -960 273710 326
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 276768 354 276796 4150
rect 278332 480 278360 9182
rect 277094 354 277206 480
rect 276768 326 277206 354
rect 277094 -960 277206 326
rect 278290 -960 278402 480
rect 279068 354 279096 16546
rect 280724 480 280752 16546
rect 281538 10568 281594 10577
rect 281538 10503 281594 10512
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281552 354 281580 10503
rect 283116 480 283144 16546
rect 284312 480 284340 72519
rect 284392 71052 284444 71058
rect 284392 70994 284444 71000
rect 284404 16574 284432 70994
rect 287060 35488 287112 35494
rect 287060 35430 287112 35436
rect 285680 28280 285732 28286
rect 285680 28222 285732 28228
rect 285692 16574 285720 28222
rect 287072 16574 287100 35430
rect 288452 16574 288480 76706
rect 296720 76696 296772 76702
rect 296720 76638 296772 76644
rect 291200 72684 291252 72690
rect 291200 72626 291252 72632
rect 289820 31340 289872 31346
rect 289820 31282 289872 31288
rect 284404 16546 284984 16574
rect 285692 16546 286640 16574
rect 287072 16546 287376 16574
rect 288452 16546 289032 16574
rect 281878 354 281990 480
rect 281552 326 281990 354
rect 281878 -960 281990 326
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 284956 354 284984 16546
rect 286612 480 286640 16546
rect 285374 354 285486 480
rect 284956 326 285486 354
rect 285374 -960 285486 326
rect 286570 -960 286682 480
rect 287348 354 287376 16546
rect 289004 480 289032 16546
rect 287766 354 287878 480
rect 287348 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 289832 354 289860 31282
rect 291212 16574 291240 72626
rect 292580 64388 292632 64394
rect 292580 64330 292632 64336
rect 291212 16546 291424 16574
rect 291396 480 291424 16546
rect 292592 480 292620 64330
rect 293960 35420 294012 35426
rect 293960 35362 294012 35368
rect 292672 24472 292724 24478
rect 292672 24414 292724 24420
rect 292684 16574 292712 24414
rect 293972 16574 294000 35362
rect 296732 16574 296760 76638
rect 318800 73976 318852 73982
rect 318800 73918 318852 73924
rect 311900 72616 311952 72622
rect 311900 72558 311952 72564
rect 298098 72448 298154 72457
rect 298098 72383 298154 72392
rect 292684 16546 293264 16574
rect 293972 16546 294920 16574
rect 296732 16546 297312 16574
rect 290158 354 290270 480
rect 289832 326 290270 354
rect 290158 -960 290270 326
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 354 293264 16546
rect 294892 480 294920 16546
rect 295616 10600 295668 10606
rect 295616 10542 295668 10548
rect 293654 354 293766 480
rect 293236 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 295628 354 295656 10542
rect 297284 480 297312 16546
rect 296046 354 296158 480
rect 295628 326 296158 354
rect 296046 -960 296158 326
rect 297242 -960 297354 480
rect 298112 354 298140 72383
rect 306380 67312 306432 67318
rect 306380 67254 306432 67260
rect 305000 35352 305052 35358
rect 305000 35294 305052 35300
rect 303620 23384 303672 23390
rect 303620 23326 303672 23332
rect 303632 16574 303660 23326
rect 305012 16574 305040 35294
rect 303632 16546 303936 16574
rect 305012 16546 305592 16574
rect 301502 13288 301558 13297
rect 301502 13223 301558 13232
rect 299662 10432 299718 10441
rect 299662 10367 299718 10376
rect 299676 480 299704 10367
rect 300766 9072 300822 9081
rect 300766 9007 300822 9016
rect 300780 480 300808 9007
rect 298438 354 298550 480
rect 298112 326 298550 354
rect 298438 -960 298550 326
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 354 301544 13223
rect 303160 3868 303212 3874
rect 303160 3810 303212 3816
rect 303172 480 303200 3810
rect 301934 354 302046 480
rect 301516 326 302046 354
rect 301934 -960 302046 326
rect 303130 -960 303242 480
rect 303908 354 303936 16546
rect 305564 480 305592 16546
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306392 354 306420 67254
rect 309140 63096 309192 63102
rect 309140 63038 309192 63044
rect 307760 35284 307812 35290
rect 307760 35226 307812 35232
rect 307772 3262 307800 35226
rect 307852 25900 307904 25906
rect 307852 25842 307904 25848
rect 307864 16574 307892 25842
rect 309152 16574 309180 63038
rect 310520 27056 310572 27062
rect 310520 26998 310572 27004
rect 310532 16574 310560 26998
rect 311912 16574 311940 72558
rect 316038 53136 316094 53145
rect 316038 53071 316094 53080
rect 307864 16546 307984 16574
rect 309152 16546 309824 16574
rect 310532 16546 311480 16574
rect 311912 16546 312216 16574
rect 307760 3256 307812 3262
rect 307760 3198 307812 3204
rect 307956 480 307984 16546
rect 309048 3256 309100 3262
rect 309048 3198 309100 3204
rect 309060 480 309088 3198
rect 306718 354 306830 480
rect 306392 326 306830 354
rect 306718 -960 306830 326
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 354 309824 16546
rect 311452 480 311480 16546
rect 310214 354 310326 480
rect 309796 326 310326 354
rect 310214 -960 310326 326
rect 311410 -960 311522 480
rect 312188 354 312216 16546
rect 313832 11960 313884 11966
rect 313832 11902 313884 11908
rect 313844 480 313872 11902
rect 315026 5128 315082 5137
rect 315026 5063 315082 5072
rect 315040 480 315068 5063
rect 316052 3262 316080 53071
rect 317418 29608 317474 29617
rect 317418 29543 317474 29552
rect 317432 16574 317460 29543
rect 318812 16574 318840 73918
rect 320180 68536 320232 68542
rect 320180 68478 320232 68484
rect 319442 21720 319498 21729
rect 319442 21655 319498 21664
rect 317432 16546 318104 16574
rect 318812 16546 319392 16574
rect 316222 16280 316278 16289
rect 316222 16215 316278 16224
rect 316040 3256 316092 3262
rect 316040 3198 316092 3204
rect 316236 480 316264 16215
rect 317328 3256 317380 3262
rect 317328 3198 317380 3204
rect 317340 480 317368 3198
rect 312606 354 312718 480
rect 312188 326 312718 354
rect 312606 -960 312718 326
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 16546
rect 319364 3482 319392 16546
rect 319456 3874 319484 21655
rect 320192 16574 320220 68478
rect 322216 28286 322244 78134
rect 324412 76628 324464 76634
rect 324412 76570 324464 76576
rect 322204 28280 322256 28286
rect 322204 28222 322256 28228
rect 320192 16546 320496 16574
rect 319444 3868 319496 3874
rect 319444 3810 319496 3816
rect 319364 3454 319760 3482
rect 319732 480 319760 3454
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320468 354 320496 16546
rect 323308 6792 323360 6798
rect 323308 6734 323360 6740
rect 322112 3392 322164 3398
rect 322112 3334 322164 3340
rect 322124 480 322152 3334
rect 323320 480 323348 6734
rect 324424 480 324452 76570
rect 396080 75608 396132 75614
rect 396080 75550 396132 75556
rect 354680 73908 354732 73914
rect 354680 73850 354732 73856
rect 340880 72548 340932 72554
rect 340880 72490 340932 72496
rect 338120 64320 338172 64326
rect 338120 64262 338172 64268
rect 332600 31272 332652 31278
rect 332600 31214 332652 31220
rect 332612 16574 332640 31214
rect 338132 16574 338160 64262
rect 339500 26988 339552 26994
rect 339500 26930 339552 26936
rect 332612 16546 332732 16574
rect 338132 16546 338712 16574
rect 326804 6724 326856 6730
rect 326804 6666 326856 6672
rect 325608 4140 325660 4146
rect 325608 4082 325660 4088
rect 325620 480 325648 4082
rect 326816 480 326844 6666
rect 329196 6656 329248 6662
rect 329196 6598 329248 6604
rect 328000 4072 328052 4078
rect 328000 4014 328052 4020
rect 328012 480 328040 4014
rect 329208 480 329236 6598
rect 330392 6588 330444 6594
rect 330392 6530 330444 6536
rect 330404 480 330432 6530
rect 331588 4004 331640 4010
rect 331588 3946 331640 3952
rect 331600 480 331628 3946
rect 332704 480 332732 16546
rect 336278 6488 336334 6497
rect 336278 6423 336334 6432
rect 333886 6216 333942 6225
rect 333886 6151 333942 6160
rect 333900 480 333928 6151
rect 335082 3632 335138 3641
rect 335082 3567 335138 3576
rect 335096 480 335124 3567
rect 336292 480 336320 6423
rect 337474 6352 337530 6361
rect 337474 6287 337530 6296
rect 337488 480 337516 6287
rect 338684 480 338712 16546
rect 320886 354 320998 480
rect 320468 326 320998 354
rect 320886 -960 320998 326
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339512 354 339540 26930
rect 340892 3210 340920 72490
rect 353298 71224 353354 71233
rect 353298 71159 353354 71168
rect 347780 67244 347832 67250
rect 347780 67186 347832 67192
rect 340972 67176 341024 67182
rect 340972 67118 341024 67124
rect 340984 3398 341012 67118
rect 346400 25832 346452 25838
rect 346400 25774 346452 25780
rect 343640 21684 343692 21690
rect 343640 21626 343692 21632
rect 343652 16574 343680 21626
rect 346412 16574 346440 25774
rect 347792 16574 347820 67186
rect 351918 47560 351974 47569
rect 351918 47495 351974 47504
rect 350538 18864 350594 18873
rect 350538 18799 350594 18808
rect 350552 16574 350580 18799
rect 351932 16574 351960 47495
rect 353312 16574 353340 71159
rect 354692 16574 354720 73850
rect 375380 73840 375432 73846
rect 375380 73782 375432 73788
rect 357440 72480 357492 72486
rect 357440 72422 357492 72428
rect 343652 16546 344600 16574
rect 346412 16546 346992 16574
rect 347792 16546 348096 16574
rect 350552 16546 351224 16574
rect 351932 16546 352880 16574
rect 353312 16546 353616 16574
rect 354692 16546 355272 16574
rect 343364 9172 343416 9178
rect 343364 9114 343416 9120
rect 340972 3392 341024 3398
rect 340972 3334 341024 3340
rect 342168 3392 342220 3398
rect 342168 3334 342220 3340
rect 340892 3182 341012 3210
rect 340984 480 341012 3182
rect 342180 480 342208 3334
rect 343376 480 343404 9114
rect 344572 480 344600 16546
rect 345296 13456 345348 13462
rect 345296 13398 345348 13404
rect 339838 354 339950 480
rect 339512 326 339950 354
rect 339838 -960 339950 326
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345308 354 345336 13398
rect 346964 480 346992 16546
rect 348068 480 348096 16546
rect 349160 13388 349212 13394
rect 349160 13330 349212 13336
rect 349172 3210 349200 13330
rect 349250 13152 349306 13161
rect 349250 13087 349306 13096
rect 349264 3398 349292 13087
rect 349252 3392 349304 3398
rect 349252 3334 349304 3340
rect 350448 3392 350500 3398
rect 350448 3334 350500 3340
rect 349172 3182 349292 3210
rect 349264 480 349292 3182
rect 350460 480 350488 3334
rect 345726 354 345838 480
rect 345308 326 345838 354
rect 345726 -960 345838 326
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351196 354 351224 16546
rect 352852 480 352880 16546
rect 351614 354 351726 480
rect 351196 326 351726 354
rect 351614 -960 351726 326
rect 352810 -960 352922 480
rect 353588 354 353616 16546
rect 355244 480 355272 16546
rect 356336 3936 356388 3942
rect 356336 3878 356388 3884
rect 356348 480 356376 3878
rect 357452 3398 357480 72422
rect 362960 68468 363012 68474
rect 362960 68410 363012 68416
rect 358820 65612 358872 65618
rect 358820 65554 358872 65560
rect 357532 31204 357584 31210
rect 357532 31146 357584 31152
rect 357440 3392 357492 3398
rect 357440 3334 357492 3340
rect 357544 480 357572 31146
rect 358832 16574 358860 65554
rect 360200 23248 360252 23254
rect 360200 23190 360252 23196
rect 360212 16574 360240 23190
rect 362972 16574 363000 68410
rect 368480 64252 368532 64258
rect 368480 64194 368532 64200
rect 367098 40624 367154 40633
rect 367098 40559 367154 40568
rect 367112 16574 367140 40559
rect 368492 16574 368520 64194
rect 374000 63028 374052 63034
rect 374000 62970 374052 62976
rect 372618 35184 372674 35193
rect 372618 35119 372674 35128
rect 372632 16574 372660 35119
rect 358832 16546 359504 16574
rect 360212 16546 361160 16574
rect 362972 16546 363552 16574
rect 367112 16546 367784 16574
rect 368492 16546 369440 16574
rect 372632 16546 372936 16574
rect 358728 3392 358780 3398
rect 358728 3334 358780 3340
rect 358740 480 358768 3334
rect 354006 354 354118 480
rect 353588 326 354118 354
rect 354006 -960 354118 326
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359476 354 359504 16546
rect 361132 480 361160 16546
rect 362316 3324 362368 3330
rect 362316 3266 362368 3272
rect 362328 480 362356 3266
rect 363524 480 363552 16546
rect 365720 13320 365772 13326
rect 365720 13262 365772 13268
rect 364616 10532 364668 10538
rect 364616 10474 364668 10480
rect 364628 480 364656 10474
rect 365732 3398 365760 13262
rect 365812 5092 365864 5098
rect 365812 5034 365864 5040
rect 365720 3392 365772 3398
rect 365720 3334 365772 3340
rect 365824 480 365852 5034
rect 367008 3392 367060 3398
rect 367008 3334 367060 3340
rect 367020 480 367048 3334
rect 359894 354 360006 480
rect 359476 326 360006 354
rect 359894 -960 360006 326
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 354 367784 16546
rect 369412 480 369440 16546
rect 371238 16144 371294 16153
rect 371238 16079 371294 16088
rect 370134 14784 370190 14793
rect 370134 14719 370190 14728
rect 368174 354 368286 480
rect 367756 326 368286 354
rect 368174 -960 368286 326
rect 369370 -960 369482 480
rect 370148 354 370176 14719
rect 370566 354 370678 480
rect 370148 326 370678 354
rect 371252 354 371280 16079
rect 372908 480 372936 16546
rect 374012 1170 374040 62970
rect 374092 24404 374144 24410
rect 374092 24346 374144 24352
rect 374104 3398 374132 24346
rect 375392 16574 375420 73782
rect 382280 70032 382332 70038
rect 382280 69974 382332 69980
rect 376760 65544 376812 65550
rect 376760 65486 376812 65492
rect 376772 16574 376800 65486
rect 379520 23180 379572 23186
rect 379520 23122 379572 23128
rect 375392 16546 376064 16574
rect 376772 16546 377720 16574
rect 374092 3392 374144 3398
rect 374092 3334 374144 3340
rect 375288 3392 375340 3398
rect 375288 3334 375340 3340
rect 374012 1142 374132 1170
rect 374104 480 374132 1142
rect 375300 480 375328 3334
rect 371670 354 371782 480
rect 371252 326 371782 354
rect 370566 -960 370678 326
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 354 376064 16546
rect 377692 480 377720 16546
rect 378416 16176 378468 16182
rect 378416 16118 378468 16124
rect 376454 354 376566 480
rect 376036 326 376566 354
rect 376454 -960 376566 326
rect 377650 -960 377762 480
rect 378428 354 378456 16118
rect 378846 354 378958 480
rect 378428 326 378958 354
rect 379532 354 379560 23122
rect 381176 14748 381228 14754
rect 381176 14690 381228 14696
rect 381188 480 381216 14690
rect 382292 3210 382320 69974
rect 390560 69964 390612 69970
rect 390560 69906 390612 69912
rect 382372 35216 382424 35222
rect 382372 35158 382424 35164
rect 382384 3398 382412 35158
rect 389180 31136 389232 31142
rect 389180 31078 389232 31084
rect 386418 25528 386474 25537
rect 386418 25463 386474 25472
rect 386432 16574 386460 25463
rect 389192 16574 389220 31078
rect 386432 16546 386736 16574
rect 389192 16546 389496 16574
rect 384304 14680 384356 14686
rect 384304 14622 384356 14628
rect 382372 3392 382424 3398
rect 382372 3334 382424 3340
rect 383568 3392 383620 3398
rect 383568 3334 383620 3340
rect 382292 3182 382412 3210
rect 382384 480 382412 3182
rect 383580 480 383608 3334
rect 379950 354 380062 480
rect 379532 326 380062 354
rect 378846 -960 378958 326
rect 379950 -960 380062 326
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384316 354 384344 14622
rect 385960 14612 386012 14618
rect 385960 14554 386012 14560
rect 385972 480 386000 14554
rect 384734 354 384846 480
rect 384316 326 384846 354
rect 384734 -960 384846 326
rect 385930 -960 386042 480
rect 386708 354 386736 16546
rect 387798 16008 387854 16017
rect 387798 15943 387854 15952
rect 387126 354 387238 480
rect 386708 326 387238 354
rect 387812 354 387840 15943
rect 389468 480 389496 16546
rect 390572 1290 390600 69906
rect 390652 42084 390704 42090
rect 390652 42026 390704 42032
rect 390560 1284 390612 1290
rect 390560 1226 390612 1232
rect 390664 480 390692 42026
rect 391940 32768 391992 32774
rect 391940 32710 391992 32716
rect 391952 16574 391980 32710
rect 391952 16546 392624 16574
rect 391848 1284 391900 1290
rect 391848 1226 391900 1232
rect 391860 480 391888 1226
rect 388230 354 388342 480
rect 387812 326 388342 354
rect 387126 -960 387238 326
rect 388230 -960 388342 326
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 354 392624 16546
rect 395344 16108 395396 16114
rect 395344 16050 395396 16056
rect 394240 10464 394292 10470
rect 394240 10406 394292 10412
rect 394252 480 394280 10406
rect 395356 480 395384 16050
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 75550
rect 402978 75440 403034 75449
rect 402978 75375 403034 75384
rect 401600 58676 401652 58682
rect 401600 58618 401652 58624
rect 397460 37936 397512 37942
rect 397460 37878 397512 37884
rect 397472 16574 397500 37878
rect 401612 16574 401640 58618
rect 402992 16574 403020 75375
rect 426440 69896 426492 69902
rect 426440 69838 426492 69844
rect 408500 62960 408552 62966
rect 408500 62902 408552 62908
rect 404360 39364 404412 39370
rect 404360 39306 404412 39312
rect 397472 16546 397776 16574
rect 401612 16546 402560 16574
rect 402992 16546 403664 16574
rect 397748 480 397776 16546
rect 398840 16040 398892 16046
rect 398840 15982 398892 15988
rect 398852 3210 398880 15982
rect 398932 10396 398984 10402
rect 398932 10338 398984 10344
rect 398944 3398 398972 10338
rect 401324 7812 401376 7818
rect 401324 7754 401376 7760
rect 398932 3392 398984 3398
rect 398932 3334 398984 3340
rect 400128 3392 400180 3398
rect 400128 3334 400180 3340
rect 398852 3182 398972 3210
rect 398944 480 398972 3182
rect 400140 480 400168 3334
rect 401336 480 401364 7754
rect 402532 480 402560 16546
rect 403636 480 403664 16546
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404372 354 404400 39306
rect 405738 17368 405794 17377
rect 405738 17303 405794 17312
rect 405752 16574 405780 17303
rect 408512 16574 408540 62902
rect 412640 61464 412692 61470
rect 412640 61406 412692 61412
rect 411260 43444 411312 43450
rect 411260 43386 411312 43392
rect 411272 16574 411300 43386
rect 405752 16546 406056 16574
rect 408512 16546 409184 16574
rect 411272 16546 411944 16574
rect 406028 480 406056 16546
rect 407210 14648 407266 14657
rect 407210 14583 407266 14592
rect 407224 480 407252 14583
rect 408406 8936 408462 8945
rect 408406 8871 408462 8880
rect 408420 480 408448 8871
rect 404790 354 404902 480
rect 404372 326 404902 354
rect 404790 -960 404902 326
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 354 409184 16546
rect 410800 6520 410852 6526
rect 410800 6462 410852 6468
rect 410812 480 410840 6462
rect 411916 480 411944 16546
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 354 412680 61406
rect 418160 40724 418212 40730
rect 418160 40666 418212 40672
rect 415400 17604 415452 17610
rect 415400 17546 415452 17552
rect 414296 11892 414348 11898
rect 414296 11834 414348 11840
rect 414308 480 414336 11834
rect 415412 3398 415440 17546
rect 418172 16574 418200 40666
rect 422298 24168 422354 24177
rect 422298 24103 422354 24112
rect 419540 17536 419592 17542
rect 419540 17478 419592 17484
rect 419552 16574 419580 17478
rect 422312 16574 422340 24103
rect 423678 18728 423734 18737
rect 423678 18663 423734 18672
rect 418172 16546 418568 16574
rect 419552 16546 420224 16574
rect 422312 16546 422616 16574
rect 417424 13252 417476 13258
rect 417424 13194 417476 13200
rect 415492 11824 415544 11830
rect 415492 11766 415544 11772
rect 415400 3392 415452 3398
rect 415400 3334 415452 3340
rect 415504 480 415532 11766
rect 416688 3392 416740 3398
rect 416688 3334 416740 3340
rect 416700 480 416728 3334
rect 413070 354 413182 480
rect 412652 326 413182 354
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 13194
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 418540 354 418568 16546
rect 420196 480 420224 16546
rect 420918 15872 420974 15881
rect 420918 15807 420974 15816
rect 418958 354 419070 480
rect 418540 326 419070 354
rect 417854 -960 417966 326
rect 418958 -960 419070 326
rect 420154 -960 420266 480
rect 420932 354 420960 15807
rect 422588 480 422616 16546
rect 423692 3210 423720 18663
rect 426452 16574 426480 69838
rect 427820 68400 427872 68406
rect 427820 68342 427872 68348
rect 427832 16574 427860 68342
rect 430592 16574 430620 80135
rect 444380 78804 444432 78810
rect 444380 78746 444432 78752
rect 431960 75540 432012 75546
rect 431960 75482 432012 75488
rect 431972 16574 432000 75482
rect 438860 75472 438912 75478
rect 438860 75414 438912 75420
rect 437480 67108 437532 67114
rect 437480 67050 437532 67056
rect 433340 60036 433392 60042
rect 433340 59978 433392 59984
rect 433352 16574 433380 59978
rect 434720 32700 434772 32706
rect 434720 32642 434772 32648
rect 434732 16574 434760 32642
rect 426452 16546 426848 16574
rect 427832 16546 428504 16574
rect 430592 16546 430896 16574
rect 431972 16546 432092 16574
rect 433352 16546 434024 16574
rect 434732 16546 435128 16574
rect 425704 15972 425756 15978
rect 425704 15914 425756 15920
rect 423770 11792 423826 11801
rect 423770 11727 423826 11736
rect 423784 3398 423812 11727
rect 423772 3392 423824 3398
rect 423772 3334 423824 3340
rect 424968 3392 425020 3398
rect 424968 3334 425020 3340
rect 423692 3182 423812 3210
rect 423784 480 423812 3182
rect 424980 480 425008 3334
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 425716 354 425744 15914
rect 426134 354 426246 480
rect 425716 326 426246 354
rect 426820 354 426848 16546
rect 428476 480 428504 16546
rect 429200 13184 429252 13190
rect 429200 13126 429252 13132
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 426134 -960 426246 326
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429212 354 429240 13126
rect 430868 480 430896 16546
rect 432064 480 432092 16546
rect 433248 6452 433300 6458
rect 433248 6394 433300 6400
rect 433260 480 433288 6394
rect 429630 354 429742 480
rect 429212 326 429742 354
rect 429630 -960 429742 326
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 433996 354 434024 16546
rect 434414 354 434526 480
rect 433996 326 434526 354
rect 435100 354 435128 16546
rect 436744 14544 436796 14550
rect 436744 14486 436796 14492
rect 436756 480 436784 14486
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 434414 -960 434526 326
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437492 354 437520 67050
rect 438872 16574 438900 75414
rect 442998 21584 443054 21593
rect 442998 21519 443054 21528
rect 440240 17468 440292 17474
rect 440240 17410 440292 17416
rect 440252 16574 440280 17410
rect 443012 16574 443040 21519
rect 444392 16574 444420 78746
rect 462332 78713 462360 703520
rect 478524 702434 478552 703520
rect 477512 702406 478552 702434
rect 477512 144226 477540 702406
rect 494808 700398 494836 703520
rect 494796 700392 494848 700398
rect 494796 700334 494848 700340
rect 477500 144220 477552 144226
rect 477500 144162 477552 144168
rect 462318 78704 462374 78713
rect 462318 78639 462374 78648
rect 471980 78124 472032 78130
rect 471980 78066 472032 78072
rect 454040 76560 454092 76566
rect 454040 76502 454092 76508
rect 447140 21616 447192 21622
rect 447140 21558 447192 21564
rect 447152 16574 447180 21558
rect 448520 18896 448572 18902
rect 448520 18838 448572 18844
rect 438872 16546 439176 16574
rect 440252 16546 440372 16574
rect 443012 16546 443408 16574
rect 444392 16546 445064 16574
rect 447152 16546 447456 16574
rect 439148 480 439176 16546
rect 440344 480 440372 16546
rect 441528 6384 441580 6390
rect 441528 6326 441580 6332
rect 441540 480 441568 6326
rect 442630 4992 442686 5001
rect 442630 4927 442686 4936
rect 442644 480 442672 4927
rect 437910 354 438022 480
rect 437492 326 438022 354
rect 437910 -960 438022 326
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443380 354 443408 16546
rect 445036 480 445064 16546
rect 446220 7744 446272 7750
rect 446220 7686 446272 7692
rect 446232 480 446260 7686
rect 447428 480 447456 16546
rect 448532 3210 448560 18838
rect 451280 18828 451332 18834
rect 451280 18770 451332 18776
rect 448612 17400 448664 17406
rect 448612 17342 448664 17348
rect 448624 3398 448652 17342
rect 451292 16574 451320 18770
rect 451292 16546 451688 16574
rect 450912 5024 450964 5030
rect 450912 4966 450964 4972
rect 448612 3392 448664 3398
rect 448612 3334 448664 3340
rect 449808 3392 449860 3398
rect 449808 3334 449860 3340
rect 448532 3182 448652 3210
rect 448624 480 448652 3182
rect 449820 480 449848 3334
rect 450924 480 450952 4966
rect 443798 354 443910 480
rect 443380 326 443910 354
rect 443798 -960 443910 326
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 451660 354 451688 16546
rect 453304 13116 453356 13122
rect 453304 13058 453356 13064
rect 453316 480 453344 13058
rect 452078 354 452190 480
rect 451660 326 452190 354
rect 452078 -960 452190 326
rect 453274 -960 453386 480
rect 454052 354 454080 76502
rect 467840 75404 467892 75410
rect 467840 75346 467892 75352
rect 462320 67040 462372 67046
rect 462320 66982 462372 66988
rect 459558 61432 459614 61441
rect 459558 61367 459614 61376
rect 456800 20188 456852 20194
rect 456800 20130 456852 20136
rect 455420 20052 455472 20058
rect 455420 19994 455472 20000
rect 455432 16574 455460 19994
rect 455432 16546 455736 16574
rect 455708 480 455736 16546
rect 456812 3398 456840 20130
rect 458178 20088 458234 20097
rect 458178 20023 458234 20032
rect 456890 17232 456946 17241
rect 456890 17167 456946 17176
rect 456800 3392 456852 3398
rect 456800 3334 456852 3340
rect 456904 480 456932 17167
rect 458192 16574 458220 20023
rect 459572 16574 459600 61367
rect 460938 21448 460994 21457
rect 460938 21383 460994 21392
rect 460952 16574 460980 21383
rect 458192 16546 459232 16574
rect 459572 16546 459968 16574
rect 460952 16546 461624 16574
rect 458088 3392 458140 3398
rect 458088 3334 458140 3340
rect 458100 480 458128 3334
rect 459204 480 459232 16546
rect 454470 354 454582 480
rect 454052 326 454582 354
rect 454470 -960 454582 326
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 16546
rect 461596 480 461624 16546
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462332 354 462360 66982
rect 463700 32632 463752 32638
rect 463700 32574 463752 32580
rect 463712 16574 463740 32574
rect 467104 24336 467156 24342
rect 467104 24278 467156 24284
rect 465080 20120 465132 20126
rect 465080 20062 465132 20068
rect 463712 16546 464016 16574
rect 463988 480 464016 16546
rect 465092 6914 465120 20062
rect 465172 19984 465224 19990
rect 465172 19926 465224 19932
rect 465184 16574 465212 19926
rect 465184 16546 465856 16574
rect 465092 6886 465212 6914
rect 465184 480 465212 6886
rect 462750 354 462862 480
rect 462332 326 462862 354
rect 462750 -960 462862 326
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 465828 354 465856 16546
rect 467116 3942 467144 24278
rect 467852 16574 467880 75346
rect 471992 16574 472020 78066
rect 480260 78056 480312 78062
rect 478878 78024 478934 78033
rect 480260 77998 480312 78004
rect 478878 77959 478934 77968
rect 473360 21548 473412 21554
rect 473360 21490 473412 21496
rect 473372 16574 473400 21490
rect 476118 21312 476174 21321
rect 476118 21247 476174 21256
rect 476132 16574 476160 21247
rect 467852 16546 468248 16574
rect 471992 16546 472296 16574
rect 473372 16546 473492 16574
rect 476132 16546 476528 16574
rect 467472 6316 467524 6322
rect 467472 6258 467524 6264
rect 467104 3936 467156 3942
rect 467104 3878 467156 3884
rect 467484 480 467512 6258
rect 466246 354 466358 480
rect 465828 326 466358 354
rect 466246 -960 466358 326
rect 467442 -960 467554 480
rect 468220 354 468248 16546
rect 471060 9104 471112 9110
rect 471060 9046 471112 9052
rect 469864 7676 469916 7682
rect 469864 7618 469916 7624
rect 469876 480 469904 7618
rect 471072 480 471100 9046
rect 472268 480 472296 16546
rect 473464 480 473492 16546
rect 474094 11656 474150 11665
rect 474094 11591 474150 11600
rect 468638 354 468750 480
rect 468220 326 468750 354
rect 468638 -960 468750 326
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474108 354 474136 11591
rect 475752 3800 475804 3806
rect 475752 3742 475804 3748
rect 475764 480 475792 3742
rect 474526 354 474638 480
rect 474108 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476500 354 476528 16546
rect 478142 14512 478198 14521
rect 478142 14447 478198 14456
rect 478156 480 478184 14447
rect 476918 354 477030 480
rect 476500 326 477030 354
rect 476918 -960 477030 326
rect 478114 -960 478226 480
rect 478892 354 478920 77959
rect 480272 16574 480300 77998
rect 498200 77988 498252 77994
rect 498200 77930 498252 77936
rect 483018 77888 483074 77897
rect 483018 77823 483074 77832
rect 481640 57316 481692 57322
rect 481640 57258 481692 57264
rect 480272 16546 480576 16574
rect 480548 480 480576 16546
rect 481652 6914 481680 57258
rect 481732 32564 481784 32570
rect 481732 32506 481784 32512
rect 481744 16574 481772 32506
rect 483032 16574 483060 77823
rect 490012 75336 490064 75342
rect 490012 75278 490064 75284
rect 496818 75304 496874 75313
rect 488540 62892 488592 62898
rect 488540 62834 488592 62840
rect 484400 21480 484452 21486
rect 484400 21422 484452 21428
rect 484412 16574 484440 21422
rect 488552 16574 488580 62834
rect 481744 16546 482416 16574
rect 483032 16546 484072 16574
rect 484412 16546 484808 16574
rect 488552 16546 488856 16574
rect 481652 6886 481772 6914
rect 481744 480 481772 6886
rect 479310 354 479422 480
rect 478892 326 479422 354
rect 479310 -960 479422 326
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482388 354 482416 16546
rect 484044 480 484072 16546
rect 482806 354 482918 480
rect 482388 326 482918 354
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 484780 354 484808 16546
rect 486424 10328 486476 10334
rect 486424 10270 486476 10276
rect 486436 480 486464 10270
rect 487620 4956 487672 4962
rect 487620 4898 487672 4904
rect 487632 480 487660 4898
rect 488828 480 488856 16546
rect 490024 6914 490052 75278
rect 496818 75239 496874 75248
rect 494058 71088 494114 71097
rect 494058 71023 494114 71032
rect 492680 17332 492732 17338
rect 492680 17274 492732 17280
rect 492692 16574 492720 17274
rect 494072 16574 494100 71023
rect 495438 19952 495494 19961
rect 495438 19887 495494 19896
rect 492692 16546 493088 16574
rect 494072 16546 494744 16574
rect 492312 9036 492364 9042
rect 492312 8978 492364 8984
rect 489932 6886 490052 6914
rect 489932 480 489960 6886
rect 491116 3732 491168 3738
rect 491116 3674 491168 3680
rect 491128 480 491156 3674
rect 492324 480 492352 8978
rect 485198 354 485310 480
rect 484780 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493060 354 493088 16546
rect 494716 480 494744 16546
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495452 354 495480 19887
rect 496832 16574 496860 75239
rect 496832 16546 497136 16574
rect 497108 480 497136 16546
rect 498212 480 498240 77930
rect 527192 77246 527220 703520
rect 543476 702434 543504 703520
rect 542372 702406 543504 702434
rect 542372 141574 542400 702406
rect 559668 700330 559696 703520
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 580262 683904 580318 683913
rect 580262 683839 580318 683848
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 579710 617536 579766 617545
rect 579710 617471 579766 617480
rect 579724 616894 579752 617471
rect 579712 616888 579764 616894
rect 579712 616830 579764 616836
rect 580170 564360 580226 564369
rect 580170 564295 580226 564304
rect 580184 563106 580212 564295
rect 580172 563100 580224 563106
rect 580172 563042 580224 563048
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 579986 431624 580042 431633
rect 579986 431559 580042 431568
rect 580000 430642 580028 431559
rect 579988 430636 580040 430642
rect 579988 430578 580040 430584
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580184 418198 580212 418231
rect 580172 418192 580224 418198
rect 580172 418134 580224 418140
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 579802 378448 579858 378457
rect 579802 378383 579858 378392
rect 579816 378214 579844 378383
rect 579804 378208 579856 378214
rect 579804 378150 579856 378156
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580080 351960 580132 351966
rect 580078 351928 580080 351937
rect 580132 351928 580134 351937
rect 580078 351863 580134 351872
rect 580078 325272 580134 325281
rect 580078 325207 580134 325216
rect 580092 324358 580120 325207
rect 580080 324352 580132 324358
rect 580080 324294 580132 324300
rect 580078 312080 580134 312089
rect 580078 312015 580134 312024
rect 580092 311914 580120 312015
rect 580080 311908 580132 311914
rect 580080 311850 580132 311856
rect 580078 298752 580134 298761
rect 580078 298687 580134 298696
rect 580092 298178 580120 298687
rect 580080 298172 580132 298178
rect 580080 298114 580132 298120
rect 579802 272232 579858 272241
rect 579802 272167 579858 272176
rect 579816 271930 579844 272167
rect 579804 271924 579856 271930
rect 579804 271866 579856 271872
rect 579986 258904 580042 258913
rect 579986 258839 580042 258848
rect 580000 258126 580028 258839
rect 579988 258120 580040 258126
rect 579988 258062 580040 258068
rect 579986 245576 580042 245585
rect 579986 245511 580042 245520
rect 580000 244322 580028 245511
rect 579988 244316 580040 244322
rect 579988 244258 580040 244264
rect 580078 232384 580134 232393
rect 580078 232319 580134 232328
rect 580092 231878 580120 232319
rect 580080 231872 580132 231878
rect 580080 231814 580132 231820
rect 580184 222902 580212 365055
rect 580172 222896 580224 222902
rect 580172 222838 580224 222844
rect 579986 219056 580042 219065
rect 579986 218991 580042 219000
rect 580000 218074 580028 218991
rect 579988 218068 580040 218074
rect 579988 218010 580040 218016
rect 580170 205728 580226 205737
rect 580170 205663 580172 205672
rect 580224 205663 580226 205672
rect 580172 205634 580224 205640
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580184 191894 580212 192471
rect 580172 191888 580224 191894
rect 580172 191830 580224 191836
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580184 178090 580212 179143
rect 580172 178084 580224 178090
rect 580172 178026 580224 178032
rect 580276 167686 580304 683839
rect 580446 630864 580502 630873
rect 580446 630799 580502 630808
rect 580354 591016 580410 591025
rect 580354 590951 580410 590960
rect 580264 167680 580316 167686
rect 580264 167622 580316 167628
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580184 165646 580212 165815
rect 580172 165640 580224 165646
rect 580172 165582 580224 165588
rect 580170 152688 580226 152697
rect 580170 152623 580226 152632
rect 580184 151842 580212 152623
rect 580172 151836 580224 151842
rect 580172 151778 580224 151784
rect 542360 141568 542412 141574
rect 542360 141510 542412 141516
rect 580172 139460 580224 139466
rect 580172 139402 580224 139408
rect 580184 139369 580212 139402
rect 580170 139360 580226 139369
rect 580170 139295 580226 139304
rect 580078 126032 580134 126041
rect 580078 125967 580134 125976
rect 580092 125662 580120 125967
rect 580080 125656 580132 125662
rect 580080 125598 580132 125604
rect 580170 112840 580226 112849
rect 580170 112775 580226 112784
rect 580184 111858 580212 112775
rect 580172 111852 580224 111858
rect 580172 111794 580224 111800
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580184 99414 580212 99447
rect 580172 99408 580224 99414
rect 580172 99350 580224 99356
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 580184 85610 580212 86119
rect 580172 85604 580224 85610
rect 580172 85546 580224 85552
rect 555424 81456 555476 81462
rect 555424 81398 555476 81404
rect 554780 78736 554832 78742
rect 554780 78678 554832 78684
rect 527180 77240 527232 77246
rect 527180 77182 527232 77188
rect 549258 76664 549314 76673
rect 549258 76599 549314 76608
rect 499580 75268 499632 75274
rect 499580 75210 499632 75216
rect 498292 23112 498344 23118
rect 498292 23054 498344 23060
rect 498304 16574 498332 23054
rect 499592 16574 499620 75210
rect 528558 75168 528614 75177
rect 528558 75103 528614 75112
rect 505100 69828 505152 69834
rect 505100 69770 505152 69776
rect 505112 16574 505140 69770
rect 518900 69760 518952 69766
rect 518900 69702 518952 69708
rect 511998 68232 512054 68241
rect 511998 68167 512054 68176
rect 507860 57248 507912 57254
rect 507860 57190 507912 57196
rect 506480 26920 506532 26926
rect 506480 26862 506532 26868
rect 498304 16546 498976 16574
rect 499592 16546 500632 16574
rect 505112 16546 505416 16574
rect 495870 354 495982 480
rect 495452 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 498948 354 498976 16546
rect 500604 480 500632 16546
rect 502984 14476 503036 14482
rect 502984 14418 503036 14424
rect 501788 3664 501840 3670
rect 501788 3606 501840 3612
rect 501800 480 501828 3606
rect 502996 480 503024 14418
rect 504180 7608 504232 7614
rect 504180 7550 504232 7556
rect 504192 480 504220 7550
rect 505388 480 505416 16546
rect 506492 3398 506520 26862
rect 506572 21412 506624 21418
rect 506572 21354 506624 21360
rect 506480 3392 506532 3398
rect 506480 3334 506532 3340
rect 506584 3210 506612 21354
rect 507872 16574 507900 57190
rect 510618 27024 510674 27033
rect 510618 26959 510674 26968
rect 509240 23044 509292 23050
rect 509240 22986 509292 22992
rect 509252 16574 509280 22986
rect 510632 16574 510660 26959
rect 507872 16546 508912 16574
rect 509252 16546 509648 16574
rect 510632 16546 511304 16574
rect 507308 3392 507360 3398
rect 507308 3334 507360 3340
rect 506492 3182 506612 3210
rect 506492 480 506520 3182
rect 499366 354 499478 480
rect 498948 326 499478 354
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507320 354 507348 3334
rect 508884 480 508912 16546
rect 507646 354 507758 480
rect 507320 326 507758 354
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 509620 354 509648 16546
rect 511276 480 511304 16546
rect 510038 354 510150 480
rect 509620 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512012 354 512040 68167
rect 514850 28248 514906 28257
rect 514850 28183 514906 28192
rect 513378 10296 513434 10305
rect 513378 10231 513434 10240
rect 512430 354 512542 480
rect 512012 326 512542 354
rect 513392 354 513420 10231
rect 514864 6914 514892 28183
rect 517520 25764 517572 25770
rect 517520 25706 517572 25712
rect 516140 22976 516192 22982
rect 516140 22918 516192 22924
rect 516152 16574 516180 22918
rect 517532 16574 517560 25706
rect 518912 16574 518940 69702
rect 525800 61396 525852 61402
rect 525800 61338 525852 61344
rect 524420 31068 524472 31074
rect 524420 31010 524472 31016
rect 521660 29708 521712 29714
rect 521660 29650 521712 29656
rect 520280 22908 520332 22914
rect 520280 22850 520332 22856
rect 516152 16546 517192 16574
rect 517532 16546 517928 16574
rect 518912 16546 519584 16574
rect 514772 6886 514892 6914
rect 514772 480 514800 6886
rect 515956 3596 516008 3602
rect 515956 3538 516008 3544
rect 515968 480 515996 3538
rect 517164 480 517192 16546
rect 513534 354 513646 480
rect 513392 326 513646 354
rect 512430 -960 512542 326
rect 513534 -960 513646 326
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 517900 354 517928 16546
rect 519556 480 519584 16546
rect 518318 354 518430 480
rect 517900 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520292 354 520320 22850
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 521672 354 521700 29650
rect 524432 16574 524460 31010
rect 525812 16574 525840 61338
rect 524432 16546 525472 16574
rect 525812 16546 526208 16574
rect 523776 11756 523828 11762
rect 523776 11698 523828 11704
rect 523040 4888 523092 4894
rect 523040 4830 523092 4836
rect 523052 480 523080 4830
rect 521814 354 521926 480
rect 521672 326 521926 354
rect 520710 -960 520822 326
rect 521814 -960 521926 326
rect 523010 -960 523122 480
rect 523788 354 523816 11698
rect 525444 480 525472 16546
rect 524206 354 524318 480
rect 523788 326 524318 354
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 526180 354 526208 16546
rect 527824 4820 527876 4826
rect 527824 4762 527876 4768
rect 527836 480 527864 4762
rect 526598 354 526710 480
rect 526180 326 526710 354
rect 526598 -960 526710 326
rect 527794 -960 527906 480
rect 528572 354 528600 75103
rect 539600 66972 539652 66978
rect 539600 66914 539652 66920
rect 529938 62928 529994 62937
rect 529938 62863 529994 62872
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 529952 354 529980 62863
rect 531318 32600 531374 32609
rect 531318 32535 531374 32544
rect 531332 3534 531360 32535
rect 535460 24268 535512 24274
rect 535460 24210 535512 24216
rect 535472 16574 535500 24210
rect 538220 24200 538272 24206
rect 538220 24142 538272 24148
rect 535472 16546 536144 16574
rect 531410 13016 531466 13025
rect 531410 12951 531466 12960
rect 531320 3528 531372 3534
rect 531320 3470 531372 3476
rect 531424 3346 531452 12951
rect 534908 3936 534960 3942
rect 534908 3878 534960 3884
rect 532148 3528 532200 3534
rect 532148 3470 532200 3476
rect 531332 3318 531452 3346
rect 531332 480 531360 3318
rect 530094 354 530206 480
rect 529952 326 530206 354
rect 528990 -960 529102 326
rect 530094 -960 530206 326
rect 531290 -960 531402 480
rect 532160 354 532188 3470
rect 533712 3460 533764 3466
rect 533712 3402 533764 3408
rect 533724 480 533752 3402
rect 534920 480 534948 3878
rect 536116 480 536144 16546
rect 537208 3392 537260 3398
rect 537208 3334 537260 3340
rect 537220 480 537248 3334
rect 532486 354 532598 480
rect 532160 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538232 354 538260 24142
rect 539612 3534 539640 66914
rect 543740 66904 543792 66910
rect 543740 66846 543792 66852
rect 539692 32496 539744 32502
rect 539692 32438 539744 32444
rect 539600 3528 539652 3534
rect 539600 3470 539652 3476
rect 539704 3346 539732 32438
rect 542360 29640 542412 29646
rect 542360 29582 542412 29588
rect 542372 16574 542400 29582
rect 543752 16574 543780 66846
rect 546498 30968 546554 30977
rect 546498 30903 546554 30912
rect 545120 17264 545172 17270
rect 545120 17206 545172 17212
rect 545132 16574 545160 17206
rect 542372 16546 542768 16574
rect 543752 16546 544424 16574
rect 545132 16546 545528 16574
rect 541992 15904 542044 15910
rect 541992 15846 542044 15852
rect 540428 3528 540480 3534
rect 540428 3470 540480 3476
rect 539612 3318 539732 3346
rect 539612 480 539640 3318
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 538374 -960 538486 326
rect 539570 -960 539682 480
rect 540440 354 540468 3470
rect 542004 480 542032 15846
rect 540766 354 540878 480
rect 540440 326 540878 354
rect 540766 -960 540878 326
rect 541962 -960 542074 480
rect 542740 354 542768 16546
rect 544396 480 544424 16546
rect 545500 480 545528 16546
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546512 354 546540 30903
rect 547878 18592 547934 18601
rect 547878 18527 547934 18536
rect 547892 16574 547920 18527
rect 549272 16574 549300 76599
rect 550638 62792 550694 62801
rect 550638 62727 550694 62736
rect 550652 16574 550680 62727
rect 552020 24132 552072 24138
rect 552020 24074 552072 24080
rect 552032 16574 552060 24074
rect 553400 18760 553452 18766
rect 553400 18702 553452 18708
rect 553412 16574 553440 18702
rect 547892 16546 548656 16574
rect 549272 16546 550312 16574
rect 550652 16546 551048 16574
rect 552032 16546 552704 16574
rect 553412 16546 553808 16574
rect 547878 4856 547934 4865
rect 547878 4791 547934 4800
rect 547892 480 547920 4791
rect 546654 354 546766 480
rect 546512 326 546766 354
rect 546654 -960 546766 326
rect 547850 -960 547962 480
rect 548628 354 548656 16546
rect 550284 480 550312 16546
rect 549046 354 549158 480
rect 548628 326 549158 354
rect 549046 -960 549158 326
rect 550242 -960 550354 480
rect 551020 354 551048 16546
rect 552676 480 552704 16546
rect 553780 480 553808 16546
rect 551438 354 551550 480
rect 551020 326 551550 354
rect 551438 -960 551550 326
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554792 354 554820 78678
rect 555436 6866 555464 81398
rect 580368 80714 580396 590951
rect 580460 160750 580488 630799
rect 580630 577688 580686 577697
rect 580630 577623 580686 577632
rect 580538 537840 580594 537849
rect 580538 537775 580594 537784
rect 580448 160744 580500 160750
rect 580448 160686 580500 160692
rect 580356 80708 580408 80714
rect 580356 80650 580408 80656
rect 580552 79354 580580 537775
rect 580644 153882 580672 577623
rect 580814 524512 580870 524521
rect 580814 524447 580870 524456
rect 580722 484664 580778 484673
rect 580722 484599 580778 484608
rect 580632 153876 580684 153882
rect 580632 153818 580684 153824
rect 580540 79348 580592 79354
rect 580540 79290 580592 79296
rect 580736 77586 580764 484599
rect 580828 141506 580856 524447
rect 580906 471472 580962 471481
rect 580906 471407 580962 471416
rect 580816 141500 580868 141506
rect 580816 141442 580868 141448
rect 580920 141438 580948 471407
rect 580908 141432 580960 141438
rect 580908 141374 580960 141380
rect 580724 77580 580776 77586
rect 580724 77522 580776 77528
rect 565818 76528 565874 76537
rect 565818 76463 565874 76472
rect 564440 75200 564492 75206
rect 564440 75142 564492 75148
rect 561680 64184 561732 64190
rect 561680 64126 561732 64132
rect 557540 62824 557592 62830
rect 557540 62766 557592 62772
rect 556160 22840 556212 22846
rect 556160 22782 556212 22788
rect 555424 6860 555476 6866
rect 555424 6802 555476 6808
rect 556172 480 556200 22782
rect 556252 18692 556304 18698
rect 556252 18634 556304 18640
rect 556264 16574 556292 18634
rect 557552 16574 557580 62766
rect 558920 25696 558972 25702
rect 558920 25638 558972 25644
rect 558932 16574 558960 25638
rect 560300 18624 560352 18630
rect 560300 18566 560352 18572
rect 560312 16574 560340 18566
rect 561692 16574 561720 64126
rect 563060 25628 563112 25634
rect 563060 25570 563112 25576
rect 556264 16546 556936 16574
rect 557552 16546 558592 16574
rect 558932 16546 559328 16574
rect 560312 16546 560432 16574
rect 561692 16546 562088 16574
rect 554934 354 555046 480
rect 554792 326 555046 354
rect 554934 -960 555046 326
rect 556130 -960 556242 480
rect 556908 354 556936 16546
rect 558564 480 558592 16546
rect 557326 354 557438 480
rect 556908 326 557438 354
rect 557326 -960 557438 326
rect 558522 -960 558634 480
rect 559300 354 559328 16546
rect 559718 354 559830 480
rect 559300 326 559830 354
rect 560404 354 560432 16546
rect 562060 480 562088 16546
rect 560822 354 560934 480
rect 560404 326 560934 354
rect 559718 -960 559830 326
rect 560822 -960 560934 326
rect 562018 -960 562130 480
rect 563072 354 563100 25570
rect 564452 480 564480 75142
rect 564532 68332 564584 68338
rect 564532 68274 564584 68280
rect 564544 16574 564572 68274
rect 565832 16574 565860 76463
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 568580 69692 568632 69698
rect 568580 69634 568632 69640
rect 567198 32464 567254 32473
rect 567198 32399 567254 32408
rect 567212 16574 567240 32399
rect 568592 16574 568620 69634
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 578238 33824 578294 33833
rect 578238 33759 578294 33768
rect 574100 32428 574152 32434
rect 574100 32370 574152 32376
rect 572720 25560 572772 25566
rect 572720 25502 572772 25508
rect 572732 16574 572760 25502
rect 574112 16574 574140 32370
rect 576858 26888 576914 26897
rect 576858 26823 576914 26832
rect 576872 16574 576900 26823
rect 578252 16574 578280 33759
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 581000 28280 581052 28286
rect 581000 28222 581052 28228
rect 580172 22772 580224 22778
rect 580172 22714 580224 22720
rect 580184 19825 580212 22714
rect 580170 19816 580226 19825
rect 580170 19751 580226 19760
rect 581012 16574 581040 28222
rect 564544 16546 565216 16574
rect 565832 16546 566872 16574
rect 567212 16546 567608 16574
rect 568592 16546 568712 16574
rect 572732 16546 573496 16574
rect 574112 16546 575152 16574
rect 576872 16546 576992 16574
rect 578252 16546 578648 16574
rect 581012 16546 581776 16574
rect 563214 354 563326 480
rect 563072 326 563326 354
rect 563214 -960 563326 326
rect 564410 -960 564522 480
rect 565188 354 565216 16546
rect 566844 480 566872 16546
rect 565606 354 565718 480
rect 565188 326 565718 354
rect 565606 -960 565718 326
rect 566802 -960 566914 480
rect 567580 354 567608 16546
rect 567998 354 568110 480
rect 567580 326 568110 354
rect 568684 354 568712 16546
rect 571524 8968 571576 8974
rect 571524 8910 571576 8916
rect 570326 3496 570382 3505
rect 570326 3431 570382 3440
rect 570340 480 570368 3431
rect 571536 480 571564 8910
rect 572720 6248 572772 6254
rect 572720 6190 572772 6196
rect 572732 480 572760 6190
rect 569102 354 569214 480
rect 568684 326 569214 354
rect 567998 -960 568110 326
rect 569102 -960 569214 326
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573468 354 573496 16546
rect 575124 480 575152 16546
rect 576308 6180 576360 6186
rect 576308 6122 576360 6128
rect 576320 480 576348 6122
rect 573886 354 573998 480
rect 573468 326 573998 354
rect 573886 -960 573998 326
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 576964 354 576992 16546
rect 578620 480 578648 16546
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 580998 3360 581054 3369
rect 580998 3295 581054 3304
rect 581012 480 581040 3295
rect 577382 354 577494 480
rect 576964 326 577494 354
rect 577382 -960 577494 326
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 581748 354 581776 16546
rect 583392 3868 583444 3874
rect 583392 3810 583444 3816
rect 583404 480 583432 3810
rect 582166 354 582278 480
rect 581748 326 582278 354
rect 582166 -960 582278 326
rect 583362 -960 583474 480
<< via2 >>
rect 2778 684256 2834 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 2778 632068 2780 632088
rect 2780 632068 2832 632088
rect 2832 632068 2834 632088
rect 2778 632032 2834 632068
rect 3054 566888 3110 566944
rect 3330 514820 3386 514856
rect 3330 514800 3332 514820
rect 3332 514800 3384 514820
rect 3384 514800 3386 514820
rect 2778 462596 2834 462632
rect 2778 462576 2780 462596
rect 2780 462576 2832 462596
rect 2832 462576 2834 462596
rect 3146 423544 3202 423600
rect 3330 410488 3386 410544
rect 3330 371320 3386 371376
rect 3330 358400 3386 358456
rect 2778 345344 2834 345400
rect 3146 319232 3202 319288
rect 3238 306176 3294 306232
rect 3146 267144 3202 267200
rect 3146 254088 3202 254144
rect 2778 241032 2834 241088
rect 3146 227976 3202 228032
rect 3146 214920 3202 214976
rect 3146 201884 3202 201920
rect 3146 201864 3148 201884
rect 3148 201864 3200 201884
rect 3200 201864 3202 201884
rect 2778 188808 2834 188864
rect 3146 162868 3148 162888
rect 3148 162868 3200 162888
rect 3200 162868 3202 162888
rect 3146 162832 3202 162868
rect 3330 293120 3386 293176
rect 3238 136740 3294 136776
rect 3238 136720 3240 136740
rect 3240 136720 3292 136740
rect 3292 136720 3294 136740
rect 3146 110608 3202 110664
rect 3238 97552 3294 97608
rect 3514 619112 3570 619168
rect 3606 606056 3662 606112
rect 3514 579944 3570 580000
rect 3514 553832 3570 553888
rect 3882 527856 3938 527912
rect 3790 501744 3846 501800
rect 3698 449520 3754 449576
rect 3514 81096 3570 81152
rect 4066 475632 4122 475688
rect 3974 397432 4030 397488
rect 3882 149776 3938 149832
rect 3698 81232 3754 81288
rect 3790 79328 3846 79384
rect 3606 79192 3662 79248
rect 3422 79056 3478 79112
rect 3238 78920 3294 78976
rect 1398 76472 1454 76528
rect 2778 75112 2834 75168
rect 3422 71576 3478 71632
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 3422 32408 3478 32464
rect 3974 84632 4030 84688
rect 117318 136856 117374 136912
rect 6918 79464 6974 79520
rect 117318 135360 117374 135416
rect 117318 133900 117320 133920
rect 117320 133900 117372 133920
rect 117372 133900 117374 133920
rect 117318 133864 117374 133900
rect 117318 132404 117320 132424
rect 117320 132404 117372 132424
rect 117372 132404 117374 132424
rect 117318 132368 117374 132404
rect 117318 130872 117374 130928
rect 117318 129376 117374 129432
rect 117318 127880 117374 127936
rect 117318 126384 117374 126440
rect 117318 124888 117374 124944
rect 117318 123392 117374 123448
rect 117318 121896 117374 121952
rect 117318 120400 117374 120456
rect 117318 118904 117374 118960
rect 117318 117408 117374 117464
rect 117318 115912 117374 115968
rect 117318 114452 117320 114472
rect 117320 114452 117372 114472
rect 117372 114452 117374 114472
rect 117318 114416 117374 114452
rect 117318 112920 117374 112976
rect 117318 111424 117374 111480
rect 117318 109928 117374 109984
rect 118054 94968 118110 95024
rect 118146 91976 118202 92032
rect 118238 90480 118294 90536
rect 118422 108432 118478 108488
rect 138110 195916 138112 195936
rect 138112 195916 138164 195936
rect 138164 195916 138166 195936
rect 138110 195880 138166 195916
rect 140410 195880 140466 195936
rect 158810 195872 158866 195928
rect 160098 195916 160100 195936
rect 160100 195916 160152 195936
rect 160152 195916 160154 195936
rect 160098 195880 160154 195916
rect 140778 195608 140834 195664
rect 139398 195472 139454 195528
rect 140870 191800 140926 191856
rect 140778 190848 140834 190904
rect 140962 191528 141018 191584
rect 140870 184320 140926 184376
rect 140778 184184 140834 184240
rect 144458 190984 144514 191040
rect 145838 188944 145894 189000
rect 140962 184048 141018 184104
rect 118790 102448 118846 102504
rect 118882 100952 118938 101008
rect 118974 99456 119030 99512
rect 144642 181056 144698 181112
rect 144734 180920 144790 180976
rect 144872 180956 144920 180976
rect 144920 180956 144928 180976
rect 144872 180920 144928 180956
rect 157798 179968 157854 180024
rect 144090 178880 144146 178936
rect 141606 178744 141662 178800
rect 143078 178744 143134 178800
rect 159454 179968 159510 180024
rect 158626 176432 158682 176488
rect 142526 172896 142582 172952
rect 154486 175344 154542 175400
rect 158442 172896 158498 172952
rect 171506 142704 171562 142760
rect 179602 135496 179658 135552
rect 179510 131960 179566 132016
rect 179418 122848 179474 122904
rect 119342 106936 119398 106992
rect 119250 105440 119306 105496
rect 119158 97960 119214 98016
rect 119066 96464 119122 96520
rect 118698 93472 118754 93528
rect 118606 88984 118662 89040
rect 118514 87488 118570 87544
rect 118330 85992 118386 86048
rect 118514 83000 118570 83056
rect 118422 81504 118478 81560
rect 20718 76608 20774 76664
rect 4066 58520 4122 58576
rect 3882 19352 3938 19408
rect 22098 43424 22154 43480
rect 3422 6432 3478 6488
rect 4066 4800 4122 4856
rect 20626 3304 20682 3360
rect 35898 75248 35954 75304
rect 40038 73752 40094 73808
rect 38382 7520 38438 7576
rect 41878 7656 41934 7712
rect 53838 75384 53894 75440
rect 57150 8880 57206 8936
rect 56046 7792 56102 7848
rect 57978 75520 58034 75576
rect 111798 76880 111854 76936
rect 93858 76744 93914 76800
rect 91098 44784 91154 44840
rect 73802 6160 73858 6216
rect 72606 3440 72662 3496
rect 78586 9016 78642 9072
rect 92478 10240 92534 10296
rect 120630 104488 120686 104544
rect 120630 84224 120686 84280
rect 120630 81368 120686 81424
rect 110510 10376 110566 10432
rect 109314 7928 109370 7984
rect 111614 6296 111670 6352
rect 178498 80960 178554 81016
rect 125736 79872 125792 79928
rect 126196 79872 126252 79928
rect 126656 79906 126712 79962
rect 125782 78784 125838 78840
rect 125598 76472 125654 76528
rect 125874 78648 125930 78704
rect 125874 77560 125930 77616
rect 126518 79600 126574 79656
rect 127208 79838 127264 79894
rect 127070 79600 127126 79656
rect 127162 77424 127218 77480
rect 127346 79600 127402 79656
rect 127668 79906 127724 79962
rect 128128 79872 128184 79928
rect 127806 79736 127862 79792
rect 127254 77288 127310 77344
rect 127070 76608 127126 76664
rect 127070 44920 127126 44976
rect 127714 79600 127770 79656
rect 128312 79736 128368 79792
rect 128772 79872 128828 79928
rect 129048 79872 129104 79928
rect 128174 79600 128230 79656
rect 129002 79736 129058 79792
rect 128726 79636 128728 79656
rect 128728 79636 128780 79656
rect 128780 79636 128782 79656
rect 128726 79600 128782 79636
rect 128542 78784 128598 78840
rect 128358 75248 128414 75304
rect 128818 78512 128874 78568
rect 129416 79872 129472 79928
rect 129784 79838 129840 79894
rect 129968 79906 130024 79962
rect 130520 79872 130576 79928
rect 129370 78512 129426 78568
rect 130566 79736 130622 79792
rect 131348 79824 131404 79826
rect 130014 78784 130070 78840
rect 129830 78648 129886 78704
rect 131348 79772 131350 79824
rect 131350 79772 131402 79824
rect 131402 79772 131404 79824
rect 131348 79770 131404 79772
rect 130382 74432 130438 74488
rect 131624 79906 131680 79962
rect 131578 79736 131634 79792
rect 131302 77016 131358 77072
rect 131210 73208 131266 73264
rect 131900 79906 131956 79962
rect 132360 79872 132416 79928
rect 132544 79906 132600 79962
rect 132728 79872 132784 79928
rect 132912 79906 132968 79962
rect 131762 78784 131818 78840
rect 131762 78376 131818 78432
rect 132222 79600 132278 79656
rect 132498 79600 132554 79656
rect 132774 79600 132830 79656
rect 133740 79872 133796 79928
rect 134016 79872 134072 79928
rect 134292 79872 134348 79928
rect 134476 79906 134532 79962
rect 134936 79872 134992 79928
rect 132774 76608 132830 76664
rect 132682 75792 132738 75848
rect 133970 76608 134026 76664
rect 134246 77016 134302 77072
rect 134614 76608 134670 76664
rect 135488 79872 135544 79928
rect 135856 79906 135912 79962
rect 136408 79906 136464 79962
rect 136592 79906 136648 79962
rect 135626 79600 135682 79656
rect 135258 74432 135314 74488
rect 135534 76608 135590 76664
rect 136546 79736 136602 79792
rect 137052 79906 137108 79962
rect 137696 79906 137752 79962
rect 138248 79906 138304 79962
rect 138616 79906 138672 79962
rect 139352 79906 139408 79962
rect 139536 79872 139592 79928
rect 136914 78104 136970 78160
rect 138202 79600 138258 79656
rect 137834 76744 137890 76800
rect 137926 76608 137982 76664
rect 138018 76472 138074 76528
rect 138984 79736 139040 79792
rect 139122 79736 139178 79792
rect 138938 79600 138994 79656
rect 139122 78648 139178 78704
rect 139352 79736 139408 79792
rect 139490 79736 139546 79792
rect 139720 79872 139776 79928
rect 140548 79906 140604 79962
rect 139306 78512 139362 78568
rect 140456 79736 140512 79792
rect 141284 79872 141340 79928
rect 140134 76336 140190 76392
rect 140410 76608 140466 76664
rect 140594 74024 140650 74080
rect 141238 79736 141294 79792
rect 141836 79872 141892 79928
rect 141146 79600 141202 79656
rect 141974 79600 142030 79656
rect 141974 78512 142030 78568
rect 142158 77016 142214 77072
rect 142066 75928 142122 75984
rect 142756 79872 142812 79928
rect 142756 79736 142812 79792
rect 141974 75520 142030 75576
rect 143400 79906 143456 79962
rect 143124 79770 143180 79826
rect 143170 79600 143226 79656
rect 143262 75928 143318 75984
rect 143630 79736 143686 79792
rect 143860 79872 143916 79928
rect 143354 75792 143410 75848
rect 143538 73888 143594 73944
rect 144458 79636 144460 79656
rect 144460 79636 144512 79656
rect 144512 79636 144514 79656
rect 144458 79600 144514 79636
rect 144366 78784 144422 78840
rect 144872 79906 144928 79962
rect 145056 79906 145112 79962
rect 145010 79736 145066 79792
rect 144826 76880 144882 76936
rect 144642 76064 144698 76120
rect 146160 79872 146216 79928
rect 146344 79872 146400 79928
rect 146712 79906 146768 79962
rect 147080 79872 147136 79928
rect 146206 79620 146262 79656
rect 146206 79600 146208 79620
rect 146208 79600 146260 79620
rect 146260 79600 146262 79620
rect 146114 75928 146170 75984
rect 146298 78512 146354 78568
rect 146758 78784 146814 78840
rect 147816 79872 147872 79928
rect 146942 78784 146998 78840
rect 146666 77968 146722 78024
rect 146206 73752 146262 73808
rect 146942 77968 146998 78024
rect 147310 77968 147366 78024
rect 147402 77288 147458 77344
rect 147770 79600 147826 79656
rect 147494 76744 147550 76800
rect 147678 77560 147734 77616
rect 147862 75928 147918 75984
rect 147586 72528 147642 72584
rect 148644 79872 148700 79928
rect 148920 79906 148976 79962
rect 149196 79872 149252 79928
rect 148874 79600 148930 79656
rect 148782 77832 148838 77888
rect 149150 79736 149206 79792
rect 149058 78376 149114 78432
rect 148966 75928 149022 75984
rect 150116 79736 150172 79792
rect 150300 79906 150356 79962
rect 149978 78648 150034 78704
rect 150760 79872 150816 79928
rect 150254 78512 150310 78568
rect 151404 79872 151460 79928
rect 151772 79736 151828 79792
rect 151956 79872 152012 79928
rect 152002 79736 152058 79792
rect 151634 76608 151690 76664
rect 151726 76472 151782 76528
rect 152600 79872 152656 79928
rect 152784 79872 152840 79928
rect 153152 79906 153208 79962
rect 152462 79600 152518 79656
rect 152738 78512 152794 78568
rect 152830 76472 152886 76528
rect 153106 79736 153162 79792
rect 153198 79600 153254 79656
rect 153704 79872 153760 79928
rect 153014 76608 153070 76664
rect 153382 77016 153438 77072
rect 153382 76608 153438 76664
rect 154072 79872 154128 79928
rect 154164 79736 154220 79792
rect 154440 79872 154496 79928
rect 154210 76336 154266 76392
rect 154394 76608 154450 76664
rect 154716 79872 154772 79928
rect 154578 79600 154634 79656
rect 154486 76472 154542 76528
rect 155452 79872 155508 79928
rect 155406 79736 155462 79792
rect 155728 79872 155784 79928
rect 156096 79872 156152 79928
rect 156556 79872 156612 79928
rect 155038 78240 155094 78296
rect 155038 78104 155094 78160
rect 155590 76608 155646 76664
rect 156510 79736 156566 79792
rect 157108 79872 157164 79928
rect 155958 77560 156014 77616
rect 156418 79600 156474 79656
rect 156418 76608 156474 76664
rect 157200 79736 157256 79792
rect 157752 79872 157808 79928
rect 157062 78104 157118 78160
rect 156970 77832 157026 77888
rect 157246 76608 157302 76664
rect 157522 76608 157578 76664
rect 158304 79736 158360 79792
rect 158488 79872 158544 79928
rect 157982 75384 158038 75440
rect 158258 79600 158314 79656
rect 158534 76608 158590 76664
rect 158442 76472 158498 76528
rect 159040 79906 159096 79962
rect 158994 79600 159050 79656
rect 159960 79872 160016 79928
rect 159730 77968 159786 78024
rect 159914 79620 159970 79656
rect 159914 79600 159916 79620
rect 159916 79600 159968 79620
rect 159968 79600 159970 79620
rect 160696 79906 160752 79962
rect 160880 79872 160936 79928
rect 160098 78784 160154 78840
rect 160374 79620 160430 79656
rect 160374 79600 160376 79620
rect 160376 79600 160428 79620
rect 160428 79600 160430 79620
rect 160374 79056 160430 79112
rect 160282 77288 160338 77344
rect 160006 76200 160062 76256
rect 160374 76336 160430 76392
rect 160742 79600 160798 79656
rect 161248 79872 161304 79928
rect 161616 79872 161672 79928
rect 161386 76608 161442 76664
rect 161110 76472 161166 76528
rect 160558 19896 160614 19952
rect 158902 4800 158958 4856
rect 161938 79736 161994 79792
rect 162444 79872 162500 79928
rect 162214 79600 162270 79656
rect 162628 79736 162684 79792
rect 162904 79736 162960 79792
rect 163272 79872 163328 79928
rect 163318 79736 163374 79792
rect 162674 79636 162676 79656
rect 162676 79636 162728 79656
rect 162728 79636 162730 79656
rect 162674 79600 162730 79636
rect 162766 78512 162822 78568
rect 162674 77560 162730 77616
rect 162858 72664 162914 72720
rect 161294 3304 161350 3360
rect 164008 79872 164064 79928
rect 163410 78648 163466 78704
rect 163962 79600 164018 79656
rect 164560 79872 164616 79928
rect 164146 79600 164202 79656
rect 164054 79056 164110 79112
rect 164422 79328 164478 79384
rect 164422 79056 164478 79112
rect 164422 76608 164478 76664
rect 164928 79872 164984 79928
rect 164790 79192 164846 79248
rect 164790 78240 164846 78296
rect 165296 79736 165352 79792
rect 165572 79872 165628 79928
rect 165250 79600 165306 79656
rect 165158 78240 165214 78296
rect 165158 77832 165214 77888
rect 165434 76608 165490 76664
rect 165940 79872 165996 79928
rect 165894 79736 165950 79792
rect 165526 76472 165582 76528
rect 166078 79600 166134 79656
rect 166768 79872 166824 79928
rect 166354 78804 166410 78840
rect 166354 78784 166356 78804
rect 166356 78784 166408 78804
rect 166408 78784 166410 78804
rect 166630 79600 166686 79656
rect 166952 79736 167008 79792
rect 167136 79872 167192 79928
rect 167320 79872 167376 79928
rect 166814 76608 166870 76664
rect 166906 75112 166962 75168
rect 167182 79600 167238 79656
rect 167504 79906 167560 79962
rect 168424 79906 168480 79962
rect 167550 76336 167606 76392
rect 168562 79736 168618 79792
rect 168102 78648 168158 78704
rect 168286 79600 168342 79656
rect 168194 76608 168250 76664
rect 169344 79872 169400 79928
rect 168838 76472 168894 76528
rect 169988 79872 170044 79928
rect 169390 78784 169446 78840
rect 169390 76608 169446 76664
rect 169574 76472 169630 76528
rect 169758 76064 169814 76120
rect 170816 79872 170872 79928
rect 169942 79600 169998 79656
rect 169850 75928 169906 75984
rect 169758 75792 169814 75848
rect 170264 79736 170320 79792
rect 170586 79736 170642 79792
rect 170126 78648 170182 78704
rect 170402 79600 170458 79656
rect 170310 76200 170366 76256
rect 170678 78784 170734 78840
rect 171046 79600 171102 79656
rect 171552 79872 171608 79928
rect 171736 79872 171792 79928
rect 171920 79872 171976 79928
rect 171138 78784 171194 78840
rect 170954 78648 171010 78704
rect 171322 78240 171378 78296
rect 171138 78104 171194 78160
rect 171506 77832 171562 77888
rect 171322 77560 171378 77616
rect 171138 77424 171194 77480
rect 170862 75792 170918 75848
rect 172380 79872 172436 79928
rect 172564 79872 172620 79928
rect 172058 78376 172114 78432
rect 172242 78104 172298 78160
rect 171966 77696 172022 77752
rect 172150 77560 172206 77616
rect 172334 77424 172390 77480
rect 173208 79736 173264 79792
rect 172978 79464 173034 79520
rect 173070 78920 173126 78976
rect 173622 79636 173624 79656
rect 173624 79636 173676 79656
rect 173676 79636 173678 79656
rect 173622 79600 173678 79636
rect 173346 79464 173402 79520
rect 173254 79328 173310 79384
rect 173438 79056 173494 79112
rect 173162 78784 173218 78840
rect 173990 79192 174046 79248
rect 172518 60016 172574 60072
rect 173254 77152 173310 77208
rect 173898 75656 173954 75712
rect 175094 79736 175150 79792
rect 176658 79872 176714 79928
rect 176566 78784 176622 78840
rect 175278 69536 175334 69592
rect 178590 80824 178646 80880
rect 178498 80008 178554 80064
rect 177302 76064 177358 76120
rect 176658 75520 176714 75576
rect 178682 72664 178738 72720
rect 180982 138624 181038 138680
rect 180890 133048 180946 133104
rect 180798 124072 180854 124128
rect 180154 81096 180210 81152
rect 181258 137536 181314 137592
rect 181166 116592 181222 116648
rect 181074 115096 181130 115152
rect 180982 88168 181038 88224
rect 180338 81368 180394 81424
rect 182178 130056 182234 130112
rect 182362 134544 182418 134600
rect 182270 128560 182326 128616
rect 182546 127064 182602 127120
rect 182454 125568 182510 125624
rect 182638 121080 182694 121136
rect 182730 119584 182786 119640
rect 182362 118088 182418 118144
rect 182270 113600 182326 113656
rect 182178 112104 182234 112160
rect 183282 110608 183338 110664
rect 183466 109112 183522 109168
rect 182270 107616 182326 107672
rect 183466 106120 183522 106176
rect 183466 104624 183522 104680
rect 183466 103128 183522 103184
rect 182914 101632 182970 101688
rect 182914 100136 182970 100192
rect 183098 98640 183154 98696
rect 183466 97144 183522 97200
rect 183190 95648 183246 95704
rect 183282 94152 183338 94208
rect 183282 92656 183338 92712
rect 183466 91160 183522 91216
rect 182178 89684 182234 89720
rect 182178 89664 182180 89684
rect 182180 89664 182232 89684
rect 182232 89664 182234 89684
rect 182178 86708 182180 86728
rect 182180 86708 182232 86728
rect 182232 86708 182234 86728
rect 182178 86672 182234 86708
rect 182638 85176 182694 85232
rect 182822 83680 182878 83736
rect 182454 82184 182510 82240
rect 194598 74024 194654 74080
rect 193218 65456 193274 65512
rect 191838 18944 191894 19000
rect 193310 28464 193366 28520
rect 213366 10648 213422 10704
rect 230478 73888 230534 73944
rect 227718 59880 227774 59936
rect 226430 34040 226486 34096
rect 229098 28328 229154 28384
rect 247038 76880 247094 76936
rect 244278 73752 244334 73808
rect 248418 20168 248474 20224
rect 246394 7656 246450 7712
rect 266358 33904 266414 33960
rect 264150 9152 264206 9208
rect 265346 7520 265402 7576
rect 396722 80960 396778 81016
rect 396906 80824 396962 80880
rect 397090 80688 397146 80744
rect 430578 80144 430634 80200
rect 397458 78784 397514 78840
rect 282918 76744 282974 76800
rect 280158 44784 280214 44840
rect 284298 72528 284354 72584
rect 281538 10512 281594 10568
rect 298098 72392 298154 72448
rect 301502 13232 301558 13288
rect 299662 10376 299718 10432
rect 300766 9016 300822 9072
rect 316038 53080 316094 53136
rect 315026 5072 315082 5128
rect 317418 29552 317474 29608
rect 319442 21664 319498 21720
rect 316222 16224 316278 16280
rect 336278 6432 336334 6488
rect 333886 6160 333942 6216
rect 335082 3576 335138 3632
rect 337474 6296 337530 6352
rect 353298 71168 353354 71224
rect 351918 47504 351974 47560
rect 350538 18808 350594 18864
rect 349250 13096 349306 13152
rect 367098 40568 367154 40624
rect 372618 35128 372674 35184
rect 371238 16088 371294 16144
rect 370134 14728 370190 14784
rect 386418 25472 386474 25528
rect 387798 15952 387854 16008
rect 402978 75384 403034 75440
rect 405738 17312 405794 17368
rect 407210 14592 407266 14648
rect 408406 8880 408462 8936
rect 422298 24112 422354 24168
rect 423678 18672 423734 18728
rect 420918 15816 420974 15872
rect 423770 11736 423826 11792
rect 442998 21528 443054 21584
rect 462318 78648 462374 78704
rect 442630 4936 442686 4992
rect 459558 61376 459614 61432
rect 458178 20032 458234 20088
rect 456890 17176 456946 17232
rect 460938 21392 460994 21448
rect 478878 77968 478934 78024
rect 476118 21256 476174 21312
rect 474094 11600 474150 11656
rect 478142 14456 478198 14512
rect 483018 77832 483074 77888
rect 496818 75248 496874 75304
rect 494058 71032 494114 71088
rect 495438 19896 495494 19952
rect 580262 683848 580318 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 579710 617480 579766 617536
rect 580170 564304 580226 564360
rect 580170 511264 580226 511320
rect 580170 458088 580226 458144
rect 579986 431568 580042 431624
rect 580170 418240 580226 418296
rect 580170 404912 580226 404968
rect 579802 378392 579858 378448
rect 580170 365064 580226 365120
rect 580078 351908 580080 351928
rect 580080 351908 580132 351928
rect 580132 351908 580134 351928
rect 580078 351872 580134 351908
rect 580078 325216 580134 325272
rect 580078 312024 580134 312080
rect 580078 298696 580134 298752
rect 579802 272176 579858 272232
rect 579986 258848 580042 258904
rect 579986 245520 580042 245576
rect 580078 232328 580134 232384
rect 579986 219000 580042 219056
rect 580170 205692 580226 205728
rect 580170 205672 580172 205692
rect 580172 205672 580224 205692
rect 580224 205672 580226 205692
rect 580170 192480 580226 192536
rect 580170 179152 580226 179208
rect 580446 630808 580502 630864
rect 580354 590960 580410 591016
rect 580170 165824 580226 165880
rect 580170 152632 580226 152688
rect 580170 139304 580226 139360
rect 580078 125976 580134 126032
rect 580170 112784 580226 112840
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 549258 76608 549314 76664
rect 528558 75112 528614 75168
rect 511998 68176 512054 68232
rect 510618 26968 510674 27024
rect 514850 28192 514906 28248
rect 513378 10240 513434 10296
rect 529938 62872 529994 62928
rect 531318 32544 531374 32600
rect 531410 12960 531466 13016
rect 546498 30912 546554 30968
rect 547878 18536 547934 18592
rect 550638 62736 550694 62792
rect 547878 4800 547934 4856
rect 580630 577632 580686 577688
rect 580538 537784 580594 537840
rect 580814 524456 580870 524512
rect 580722 484608 580778 484664
rect 580906 471416 580962 471472
rect 565818 76472 565874 76528
rect 580170 72936 580226 72992
rect 567198 32408 567254 32464
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 578238 33768 578294 33824
rect 576858 26832 576914 26888
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 580170 19760 580226 19816
rect 570326 3440 570382 3496
rect 580170 6568 580226 6624
rect 580998 3304 581054 3360
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697234 584960 697324
rect 567150 697174 584960 697234
rect 396574 696900 396580 696964
rect 396644 696962 396650 696964
rect 567150 696962 567210 697174
rect 583520 697084 584960 697174
rect 396644 696902 567210 696962
rect 396644 696900 396650 696902
rect -960 684314 480 684404
rect 2773 684314 2839 684317
rect -960 684312 2839 684314
rect -960 684256 2778 684312
rect 2834 684256 2839 684312
rect -960 684254 2839 684256
rect -960 684164 480 684254
rect 2773 684251 2839 684254
rect 580257 683906 580323 683909
rect 583520 683906 584960 683996
rect 580257 683904 584960 683906
rect 580257 683848 580262 683904
rect 580318 683848 584960 683904
rect 580257 683846 584960 683848
rect 580257 683843 580323 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 644058 584960 644148
rect 583342 643998 584960 644058
rect 583342 643922 583402 643998
rect 583520 643922 584960 643998
rect 583342 643908 584960 643922
rect 583342 643862 583586 643908
rect 396758 643180 396764 643244
rect 396828 643242 396834 643244
rect 583526 643242 583586 643862
rect 396828 643182 583586 643242
rect 396828 643180 396834 643182
rect -960 632090 480 632180
rect 2773 632090 2839 632093
rect -960 632088 2839 632090
rect -960 632032 2778 632088
rect 2834 632032 2839 632088
rect -960 632030 2839 632032
rect -960 631940 480 632030
rect 2773 632027 2839 632030
rect 580441 630866 580507 630869
rect 583520 630866 584960 630956
rect 580441 630864 584960 630866
rect 580441 630808 580446 630864
rect 580502 630808 584960 630864
rect 580441 630806 584960 630808
rect 580441 630803 580507 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3509 619170 3575 619173
rect -960 619168 3575 619170
rect -960 619112 3514 619168
rect 3570 619112 3575 619168
rect -960 619110 3575 619112
rect -960 619020 480 619110
rect 3509 619107 3575 619110
rect 579705 617538 579771 617541
rect 583520 617538 584960 617628
rect 579705 617536 584960 617538
rect 579705 617480 579710 617536
rect 579766 617480 584960 617536
rect 579705 617478 584960 617480
rect 579705 617475 579771 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3601 606114 3667 606117
rect -960 606112 3667 606114
rect -960 606056 3606 606112
rect 3662 606056 3667 606112
rect -960 606054 3667 606056
rect -960 605964 480 606054
rect 3601 606051 3667 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580349 591018 580415 591021
rect 583520 591018 584960 591108
rect 580349 591016 584960 591018
rect 580349 590960 580354 591016
rect 580410 590960 584960 591016
rect 580349 590958 584960 590960
rect 580349 590955 580415 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3509 580002 3575 580005
rect -960 580000 3575 580002
rect -960 579944 3514 580000
rect 3570 579944 3575 580000
rect -960 579942 3575 579944
rect -960 579852 480 579942
rect 3509 579939 3575 579942
rect 580625 577690 580691 577693
rect 583520 577690 584960 577780
rect 580625 577688 584960 577690
rect 580625 577632 580630 577688
rect 580686 577632 584960 577688
rect 580625 577630 584960 577632
rect 580625 577627 580691 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3049 566946 3115 566949
rect -960 566944 3115 566946
rect -960 566888 3054 566944
rect 3110 566888 3115 566944
rect -960 566886 3115 566888
rect -960 566796 480 566886
rect 3049 566883 3115 566886
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3509 553890 3575 553893
rect -960 553888 3575 553890
rect -960 553832 3514 553888
rect 3570 553832 3575 553888
rect -960 553830 3575 553832
rect -960 553740 480 553830
rect 3509 553827 3575 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580533 537842 580599 537845
rect 583520 537842 584960 537932
rect 580533 537840 584960 537842
rect 580533 537784 580538 537840
rect 580594 537784 584960 537840
rect 580533 537782 584960 537784
rect 580533 537779 580599 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3877 527914 3943 527917
rect -960 527912 3943 527914
rect -960 527856 3882 527912
rect 3938 527856 3943 527912
rect -960 527854 3943 527856
rect -960 527764 480 527854
rect 3877 527851 3943 527854
rect 580809 524514 580875 524517
rect 583520 524514 584960 524604
rect 580809 524512 584960 524514
rect 580809 524456 580814 524512
rect 580870 524456 584960 524512
rect 580809 524454 584960 524456
rect 580809 524451 580875 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3325 514858 3391 514861
rect -960 514856 3391 514858
rect -960 514800 3330 514856
rect 3386 514800 3391 514856
rect -960 514798 3391 514800
rect -960 514708 480 514798
rect 3325 514795 3391 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3785 501802 3851 501805
rect -960 501800 3851 501802
rect -960 501744 3790 501800
rect 3846 501744 3851 501800
rect -960 501742 3851 501744
rect -960 501652 480 501742
rect 3785 501739 3851 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580717 484666 580783 484669
rect 583520 484666 584960 484756
rect 580717 484664 584960 484666
rect 580717 484608 580722 484664
rect 580778 484608 584960 484664
rect 580717 484606 584960 484608
rect 580717 484603 580783 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 4061 475690 4127 475693
rect -960 475688 4127 475690
rect -960 475632 4066 475688
rect 4122 475632 4127 475688
rect -960 475630 4127 475632
rect -960 475540 480 475630
rect 4061 475627 4127 475630
rect 580901 471474 580967 471477
rect 583520 471474 584960 471564
rect 580901 471472 584960 471474
rect 580901 471416 580906 471472
rect 580962 471416 584960 471472
rect 580901 471414 584960 471416
rect 580901 471411 580967 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 2773 462634 2839 462637
rect -960 462632 2839 462634
rect -960 462576 2778 462632
rect 2834 462576 2839 462632
rect -960 462574 2839 462576
rect -960 462484 480 462574
rect 2773 462571 2839 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3693 449578 3759 449581
rect -960 449576 3759 449578
rect -960 449520 3698 449576
rect 3754 449520 3759 449576
rect -960 449518 3759 449520
rect -960 449428 480 449518
rect 3693 449515 3759 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 579981 431626 580047 431629
rect 583520 431626 584960 431716
rect 579981 431624 584960 431626
rect 579981 431568 579986 431624
rect 580042 431568 584960 431624
rect 579981 431566 584960 431568
rect 579981 431563 580047 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3141 423602 3207 423605
rect -960 423600 3207 423602
rect -960 423544 3146 423600
rect 3202 423544 3207 423600
rect -960 423542 3207 423544
rect -960 423452 480 423542
rect 3141 423539 3207 423542
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3325 410546 3391 410549
rect -960 410544 3391 410546
rect -960 410488 3330 410544
rect 3386 410488 3391 410544
rect -960 410486 3391 410488
rect -960 410396 480 410486
rect 3325 410483 3391 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3969 397490 4035 397493
rect -960 397488 4035 397490
rect -960 397432 3974 397488
rect 4030 397432 4035 397488
rect -960 397430 4035 397432
rect -960 397340 480 397430
rect 3969 397427 4035 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 579797 378450 579863 378453
rect 583520 378450 584960 378540
rect 579797 378448 584960 378450
rect 579797 378392 579802 378448
rect 579858 378392 584960 378448
rect 579797 378390 584960 378392
rect 579797 378387 579863 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3325 371378 3391 371381
rect -960 371376 3391 371378
rect -960 371320 3330 371376
rect 3386 371320 3391 371376
rect -960 371318 3391 371320
rect -960 371228 480 371318
rect 3325 371315 3391 371318
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3325 358458 3391 358461
rect -960 358456 3391 358458
rect -960 358400 3330 358456
rect 3386 358400 3391 358456
rect -960 358398 3391 358400
rect -960 358308 480 358398
rect 3325 358395 3391 358398
rect 580073 351930 580139 351933
rect 583520 351930 584960 352020
rect 580073 351928 584960 351930
rect 580073 351872 580078 351928
rect 580134 351872 584960 351928
rect 580073 351870 584960 351872
rect 580073 351867 580139 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 2773 345402 2839 345405
rect -960 345400 2839 345402
rect -960 345344 2778 345400
rect 2834 345344 2839 345400
rect -960 345342 2839 345344
rect -960 345252 480 345342
rect 2773 345339 2839 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 580073 325274 580139 325277
rect 583520 325274 584960 325364
rect 580073 325272 584960 325274
rect 580073 325216 580078 325272
rect 580134 325216 584960 325272
rect 580073 325214 584960 325216
rect 580073 325211 580139 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3141 319290 3207 319293
rect -960 319288 3207 319290
rect -960 319232 3146 319288
rect 3202 319232 3207 319288
rect -960 319230 3207 319232
rect -960 319140 480 319230
rect 3141 319227 3207 319230
rect 580073 312082 580139 312085
rect 583520 312082 584960 312172
rect 580073 312080 584960 312082
rect 580073 312024 580078 312080
rect 580134 312024 584960 312080
rect 580073 312022 584960 312024
rect 580073 312019 580139 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3233 306234 3299 306237
rect -960 306232 3299 306234
rect -960 306176 3238 306232
rect 3294 306176 3299 306232
rect -960 306174 3299 306176
rect -960 306084 480 306174
rect 3233 306171 3299 306174
rect 580073 298754 580139 298757
rect 583520 298754 584960 298844
rect 580073 298752 584960 298754
rect 580073 298696 580078 298752
rect 580134 298696 584960 298752
rect 580073 298694 584960 298696
rect 580073 298691 580139 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3325 293178 3391 293181
rect -960 293176 3391 293178
rect -960 293120 3330 293176
rect 3386 293120 3391 293176
rect -960 293118 3391 293120
rect -960 293028 480 293118
rect 3325 293115 3391 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 579797 272234 579863 272237
rect 583520 272234 584960 272324
rect 579797 272232 584960 272234
rect 579797 272176 579802 272232
rect 579858 272176 584960 272232
rect 579797 272174 584960 272176
rect 579797 272171 579863 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3141 267202 3207 267205
rect -960 267200 3207 267202
rect -960 267144 3146 267200
rect 3202 267144 3207 267200
rect -960 267142 3207 267144
rect -960 267052 480 267142
rect 3141 267139 3207 267142
rect 579981 258906 580047 258909
rect 583520 258906 584960 258996
rect 579981 258904 584960 258906
rect 579981 258848 579986 258904
rect 580042 258848 584960 258904
rect 579981 258846 584960 258848
rect 579981 258843 580047 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3141 254146 3207 254149
rect -960 254144 3207 254146
rect -960 254088 3146 254144
rect 3202 254088 3207 254144
rect -960 254086 3207 254088
rect -960 253996 480 254086
rect 3141 254083 3207 254086
rect 579981 245578 580047 245581
rect 583520 245578 584960 245668
rect 579981 245576 584960 245578
rect 579981 245520 579986 245576
rect 580042 245520 584960 245576
rect 579981 245518 584960 245520
rect 579981 245515 580047 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 2773 241090 2839 241093
rect -960 241088 2839 241090
rect -960 241032 2778 241088
rect 2834 241032 2839 241088
rect -960 241030 2839 241032
rect -960 240940 480 241030
rect 2773 241027 2839 241030
rect 580073 232386 580139 232389
rect 583520 232386 584960 232476
rect 580073 232384 584960 232386
rect 580073 232328 580078 232384
rect 580134 232328 584960 232384
rect 580073 232326 584960 232328
rect 580073 232323 580139 232326
rect 583520 232236 584960 232326
rect -960 228034 480 228124
rect 3141 228034 3207 228037
rect -960 228032 3207 228034
rect -960 227976 3146 228032
rect 3202 227976 3207 228032
rect -960 227974 3207 227976
rect -960 227884 480 227974
rect 3141 227971 3207 227974
rect 579981 219058 580047 219061
rect 583520 219058 584960 219148
rect 579981 219056 584960 219058
rect 579981 219000 579986 219056
rect 580042 219000 584960 219056
rect 579981 218998 584960 219000
rect 579981 218995 580047 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3141 214978 3207 214981
rect -960 214976 3207 214978
rect -960 214920 3146 214976
rect 3202 214920 3207 214976
rect -960 214918 3207 214920
rect -960 214828 480 214918
rect 3141 214915 3207 214918
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 580165 205667 580231 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3141 201922 3207 201925
rect -960 201920 3207 201922
rect -960 201864 3146 201920
rect 3202 201864 3207 201920
rect -960 201862 3207 201864
rect -960 201772 480 201862
rect 3141 201859 3207 201862
rect 138105 195938 138171 195941
rect 140405 195938 140471 195941
rect 160093 195938 160159 195941
rect 138105 195936 140471 195938
rect 138105 195880 138110 195936
rect 138166 195880 140410 195936
rect 140466 195880 140471 195936
rect 158854 195936 160159 195938
rect 158854 195933 160098 195936
rect 138105 195878 140471 195880
rect 138105 195875 138171 195878
rect 140405 195875 140471 195878
rect 158805 195928 160098 195933
rect 158805 195872 158810 195928
rect 158866 195880 160098 195928
rect 160154 195880 160159 195936
rect 158866 195878 160159 195880
rect 158866 195872 158914 195878
rect 160093 195875 160159 195878
rect 158805 195870 158914 195872
rect 158805 195867 158871 195870
rect 140773 195666 140839 195669
rect 143582 195666 144164 195674
rect 140773 195664 144164 195666
rect 140773 195608 140778 195664
rect 140834 195614 144164 195664
rect 140834 195608 143642 195614
rect 140773 195606 143642 195608
rect 140773 195603 140839 195606
rect 139393 195530 139459 195533
rect 139393 195528 142170 195530
rect 139393 195472 139398 195528
rect 139454 195498 142170 195528
rect 139454 195472 142692 195498
rect 139393 195470 142692 195472
rect 139393 195467 139459 195470
rect 142110 195438 142692 195470
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect 140865 191858 140931 191861
rect 143582 191858 143980 191900
rect 140865 191856 143980 191858
rect 140865 191800 140870 191856
rect 140926 191840 143980 191856
rect 140926 191800 143642 191840
rect 140865 191798 143642 191800
rect 140865 191795 140931 191798
rect 140957 191586 141023 191589
rect 143582 191586 144164 191630
rect 140957 191584 144164 191586
rect 140957 191528 140962 191584
rect 141018 191570 144164 191584
rect 141018 191528 143642 191570
rect 140957 191526 143642 191528
rect 140957 191523 141023 191526
rect 140773 190906 140839 190909
rect 144134 190906 144194 191460
rect 144453 191044 144519 191045
rect 144453 191040 144500 191044
rect 144564 191042 144570 191044
rect 144453 190984 144458 191040
rect 144453 190980 144500 190984
rect 144564 190982 144610 191042
rect 144564 190980 144570 190982
rect 144453 190979 144519 190980
rect 140773 190904 144194 190906
rect 140773 190848 140778 190904
rect 140834 190848 144194 190904
rect 140773 190846 144194 190848
rect 140773 190843 140839 190846
rect 145833 189000 145899 189005
rect -960 188866 480 188956
rect 145833 188944 145838 189000
rect 145894 188944 145899 189000
rect 145833 188939 145899 188944
rect 2773 188866 2839 188869
rect -960 188864 2839 188866
rect -960 188808 2778 188864
rect 2834 188808 2839 188864
rect -960 188806 2839 188808
rect -960 188716 480 188806
rect 2773 188803 2839 188806
rect 145836 188594 145896 188939
rect 146150 188594 146156 188596
rect 145836 188534 146156 188594
rect 146150 188532 146156 188534
rect 146220 188532 146226 188596
rect 144494 185948 144500 186012
rect 144564 186010 144570 186012
rect 146334 186010 146340 186012
rect 144564 185950 146340 186010
rect 144564 185948 144570 185950
rect 146334 185948 146340 185950
rect 146404 185948 146410 186012
rect 140865 184378 140931 184381
rect 142838 184378 142844 184380
rect 140865 184376 142844 184378
rect 140865 184320 140870 184376
rect 140926 184320 142844 184376
rect 140865 184318 142844 184320
rect 140865 184315 140931 184318
rect 142838 184316 142844 184318
rect 142908 184316 142914 184380
rect 140773 184242 140839 184245
rect 140998 184242 141004 184244
rect 140773 184240 141004 184242
rect 140773 184184 140778 184240
rect 140834 184184 141004 184240
rect 140773 184182 141004 184184
rect 140773 184179 140839 184182
rect 140998 184180 141004 184182
rect 141068 184180 141074 184244
rect 140957 184106 141023 184109
rect 143022 184106 143028 184108
rect 140957 184104 143028 184106
rect 140957 184048 140962 184104
rect 141018 184048 143028 184104
rect 140957 184046 143028 184048
rect 140957 184043 141023 184046
rect 143022 184044 143028 184046
rect 143092 184044 143098 184108
rect 142470 181052 142476 181116
rect 142540 181114 142546 181116
rect 144637 181114 144703 181117
rect 142540 181112 144703 181114
rect 142540 181056 144642 181112
rect 144698 181056 144703 181112
rect 142540 181054 144703 181056
rect 142540 181052 142546 181054
rect 144637 181051 144703 181054
rect 144729 180978 144795 180981
rect 144867 180978 144933 180981
rect 144729 180976 144933 180978
rect 144729 180920 144734 180976
rect 144790 180920 144872 180976
rect 144928 180920 144933 180976
rect 144729 180918 144933 180920
rect 144729 180915 144795 180918
rect 144867 180915 144933 180918
rect 157793 180026 157859 180029
rect 159449 180026 159515 180029
rect 157793 180024 159515 180026
rect 157793 179968 157798 180024
rect 157854 179968 159454 180024
rect 159510 179968 159515 180024
rect 157793 179966 159515 179968
rect 157793 179963 157859 179966
rect 159449 179963 159515 179966
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect 143022 178876 143028 178940
rect 143092 178938 143098 178940
rect 144085 178938 144151 178941
rect 143092 178936 144151 178938
rect 143092 178880 144090 178936
rect 144146 178880 144151 178936
rect 143092 178878 144151 178880
rect 143092 178876 143098 178878
rect 144085 178875 144151 178878
rect 140998 178740 141004 178804
rect 141068 178802 141074 178804
rect 141601 178802 141667 178805
rect 141068 178800 141667 178802
rect 141068 178744 141606 178800
rect 141662 178744 141667 178800
rect 141068 178742 141667 178744
rect 141068 178740 141074 178742
rect 141601 178739 141667 178742
rect 142838 178740 142844 178804
rect 142908 178802 142914 178804
rect 143073 178802 143139 178805
rect 142908 178800 143139 178802
rect 142908 178744 143078 178800
rect 143134 178744 143139 178800
rect 142908 178742 143139 178744
rect 142908 178740 142914 178742
rect 143073 178739 143139 178742
rect 158478 176428 158484 176492
rect 158548 176490 158554 176492
rect 158621 176490 158687 176493
rect 158548 176488 158687 176490
rect 158548 176432 158626 176488
rect 158682 176432 158687 176488
rect 158548 176430 158687 176432
rect 158548 176428 158554 176430
rect 158621 176427 158687 176430
rect -960 175796 480 176036
rect 146334 175340 146340 175404
rect 146404 175402 146410 175404
rect 154481 175402 154547 175405
rect 146404 175400 154547 175402
rect 146404 175344 154486 175400
rect 154542 175344 154547 175400
rect 146404 175342 154547 175344
rect 146404 175340 146410 175342
rect 154481 175339 154547 175342
rect 142521 172956 142587 172957
rect 142470 172954 142476 172956
rect 142430 172894 142476 172954
rect 142540 172952 142587 172956
rect 158437 172956 158503 172957
rect 158437 172954 158484 172956
rect 142582 172896 142587 172952
rect 142470 172892 142476 172894
rect 142540 172892 142587 172896
rect 158392 172952 158484 172954
rect 158392 172896 158442 172952
rect 158392 172894 158484 172896
rect 142521 172891 142587 172892
rect 158437 172892 158484 172894
rect 158548 172892 158554 172956
rect 158437 172891 158503 172892
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3141 162890 3207 162893
rect -960 162888 3207 162890
rect -960 162832 3146 162888
rect 3202 162832 3207 162888
rect -960 162830 3207 162832
rect -960 162740 480 162830
rect 3141 162827 3207 162830
rect 580165 152690 580231 152693
rect 583520 152690 584960 152780
rect 580165 152688 584960 152690
rect 580165 152632 580170 152688
rect 580226 152632 584960 152688
rect 580165 152630 584960 152632
rect 580165 152627 580231 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3877 149834 3943 149837
rect -960 149832 3943 149834
rect -960 149776 3882 149832
rect 3938 149776 3943 149832
rect -960 149774 3943 149776
rect -960 149684 480 149774
rect 3877 149771 3943 149774
rect 146150 142700 146156 142764
rect 146220 142762 146226 142764
rect 171501 142762 171567 142765
rect 146220 142760 171567 142762
rect 146220 142704 171506 142760
rect 171562 142704 171567 142760
rect 146220 142702 171567 142704
rect 146220 142700 146226 142702
rect 171501 142699 171567 142702
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect 180977 138682 181043 138685
rect 120582 138680 181043 138682
rect 120582 138624 180982 138680
rect 181038 138624 181043 138680
rect 120582 138622 181043 138624
rect 120582 138380 120642 138622
rect 180977 138619 181043 138622
rect 181253 137594 181319 137597
rect 179860 137592 181319 137594
rect 179860 137536 181258 137592
rect 181314 137536 181319 137592
rect 179860 137534 181319 137536
rect 181253 137531 181319 137534
rect 117313 136914 117379 136917
rect 117313 136912 120060 136914
rect -960 136778 480 136868
rect 117313 136856 117318 136912
rect 117374 136856 120060 136912
rect 117313 136854 120060 136856
rect 117313 136851 117379 136854
rect 3233 136778 3299 136781
rect -960 136776 3299 136778
rect -960 136720 3238 136776
rect 3294 136720 3299 136776
rect -960 136718 3299 136720
rect -960 136628 480 136718
rect 3233 136715 3299 136718
rect 179646 135557 179706 136068
rect 179597 135552 179706 135557
rect 179597 135496 179602 135552
rect 179658 135496 179706 135552
rect 179597 135494 179706 135496
rect 179597 135491 179663 135494
rect 117313 135418 117379 135421
rect 117313 135416 120060 135418
rect 117313 135360 117318 135416
rect 117374 135360 120060 135416
rect 117313 135358 120060 135360
rect 117313 135355 117379 135358
rect 182357 134602 182423 134605
rect 179860 134600 182423 134602
rect 179860 134544 182362 134600
rect 182418 134544 182423 134600
rect 179860 134542 182423 134544
rect 182357 134539 182423 134542
rect 117313 133922 117379 133925
rect 117313 133920 120060 133922
rect 117313 133864 117318 133920
rect 117374 133864 120060 133920
rect 117313 133862 120060 133864
rect 117313 133859 117379 133862
rect 180885 133106 180951 133109
rect 179860 133104 180951 133106
rect 179860 133048 180890 133104
rect 180946 133048 180951 133104
rect 179860 133046 180951 133048
rect 180885 133043 180951 133046
rect 117313 132426 117379 132429
rect 117313 132424 120060 132426
rect 117313 132368 117318 132424
rect 117374 132368 120060 132424
rect 117313 132366 120060 132368
rect 117313 132363 117379 132366
rect 179505 132018 179571 132021
rect 179462 132016 179571 132018
rect 179462 131960 179510 132016
rect 179566 131960 179571 132016
rect 179462 131955 179571 131960
rect 179462 131580 179522 131955
rect 117313 130930 117379 130933
rect 117313 130928 120060 130930
rect 117313 130872 117318 130928
rect 117374 130872 120060 130928
rect 117313 130870 120060 130872
rect 117313 130867 117379 130870
rect 182173 130114 182239 130117
rect 179860 130112 182239 130114
rect 179860 130056 182178 130112
rect 182234 130056 182239 130112
rect 179860 130054 182239 130056
rect 182173 130051 182239 130054
rect 117313 129434 117379 129437
rect 117313 129432 120060 129434
rect 117313 129376 117318 129432
rect 117374 129376 120060 129432
rect 117313 129374 120060 129376
rect 117313 129371 117379 129374
rect 182265 128618 182331 128621
rect 179860 128616 182331 128618
rect 179860 128560 182270 128616
rect 182326 128560 182331 128616
rect 179860 128558 182331 128560
rect 182265 128555 182331 128558
rect 117313 127938 117379 127941
rect 117313 127936 120060 127938
rect 117313 127880 117318 127936
rect 117374 127880 120060 127936
rect 117313 127878 120060 127880
rect 117313 127875 117379 127878
rect 182541 127122 182607 127125
rect 179860 127120 182607 127122
rect 179860 127064 182546 127120
rect 182602 127064 182607 127120
rect 179860 127062 182607 127064
rect 182541 127059 182607 127062
rect 117313 126442 117379 126445
rect 117313 126440 120060 126442
rect 117313 126384 117318 126440
rect 117374 126384 120060 126440
rect 117313 126382 120060 126384
rect 117313 126379 117379 126382
rect 580073 126034 580139 126037
rect 583520 126034 584960 126124
rect 580073 126032 584960 126034
rect 580073 125976 580078 126032
rect 580134 125976 584960 126032
rect 580073 125974 584960 125976
rect 580073 125971 580139 125974
rect 583520 125884 584960 125974
rect 182449 125626 182515 125629
rect 179860 125624 182515 125626
rect 179860 125568 182454 125624
rect 182510 125568 182515 125624
rect 179860 125566 182515 125568
rect 182449 125563 182515 125566
rect 117313 124946 117379 124949
rect 117313 124944 120060 124946
rect 117313 124888 117318 124944
rect 117374 124888 120060 124944
rect 117313 124886 120060 124888
rect 117313 124883 117379 124886
rect 180793 124130 180859 124133
rect 179860 124128 180859 124130
rect 179860 124072 180798 124128
rect 180854 124072 180859 124128
rect 179860 124070 180859 124072
rect 180793 124067 180859 124070
rect -960 123572 480 123812
rect 117313 123450 117379 123453
rect 117313 123448 120060 123450
rect 117313 123392 117318 123448
rect 117374 123392 120060 123448
rect 117313 123390 120060 123392
rect 117313 123387 117379 123390
rect 179413 122906 179479 122909
rect 179413 122904 179522 122906
rect 179413 122848 179418 122904
rect 179474 122848 179522 122904
rect 179413 122843 179522 122848
rect 179462 122604 179522 122843
rect 117313 121954 117379 121957
rect 117313 121952 120060 121954
rect 117313 121896 117318 121952
rect 117374 121896 120060 121952
rect 117313 121894 120060 121896
rect 117313 121891 117379 121894
rect 182633 121138 182699 121141
rect 179860 121136 182699 121138
rect 179860 121080 182638 121136
rect 182694 121080 182699 121136
rect 179860 121078 182699 121080
rect 182633 121075 182699 121078
rect 117313 120458 117379 120461
rect 117313 120456 120060 120458
rect 117313 120400 117318 120456
rect 117374 120400 120060 120456
rect 117313 120398 120060 120400
rect 117313 120395 117379 120398
rect 182725 119642 182791 119645
rect 179860 119640 182791 119642
rect 179860 119584 182730 119640
rect 182786 119584 182791 119640
rect 179860 119582 182791 119584
rect 182725 119579 182791 119582
rect 117313 118962 117379 118965
rect 117313 118960 120060 118962
rect 117313 118904 117318 118960
rect 117374 118904 120060 118960
rect 117313 118902 120060 118904
rect 117313 118899 117379 118902
rect 182357 118146 182423 118149
rect 179860 118144 182423 118146
rect 179860 118088 182362 118144
rect 182418 118088 182423 118144
rect 179860 118086 182423 118088
rect 182357 118083 182423 118086
rect 117313 117466 117379 117469
rect 117313 117464 120060 117466
rect 117313 117408 117318 117464
rect 117374 117408 120060 117464
rect 117313 117406 120060 117408
rect 117313 117403 117379 117406
rect 181161 116650 181227 116653
rect 179860 116648 181227 116650
rect 179860 116592 181166 116648
rect 181222 116592 181227 116648
rect 179860 116590 181227 116592
rect 181161 116587 181227 116590
rect 117313 115970 117379 115973
rect 117313 115968 120060 115970
rect 117313 115912 117318 115968
rect 117374 115912 120060 115968
rect 117313 115910 120060 115912
rect 117313 115907 117379 115910
rect 181069 115154 181135 115157
rect 179860 115152 181135 115154
rect 179860 115096 181074 115152
rect 181130 115096 181135 115152
rect 179860 115094 181135 115096
rect 181069 115091 181135 115094
rect 117313 114474 117379 114477
rect 117313 114472 120060 114474
rect 117313 114416 117318 114472
rect 117374 114416 120060 114472
rect 117313 114414 120060 114416
rect 117313 114411 117379 114414
rect 182265 113658 182331 113661
rect 179860 113656 182331 113658
rect 179860 113600 182270 113656
rect 182326 113600 182331 113656
rect 179860 113598 182331 113600
rect 182265 113595 182331 113598
rect 117313 112978 117379 112981
rect 117313 112976 120060 112978
rect 117313 112920 117318 112976
rect 117374 112920 120060 112976
rect 117313 112918 120060 112920
rect 117313 112915 117379 112918
rect 580165 112842 580231 112845
rect 583520 112842 584960 112932
rect 580165 112840 584960 112842
rect 580165 112784 580170 112840
rect 580226 112784 584960 112840
rect 580165 112782 584960 112784
rect 580165 112779 580231 112782
rect 583520 112692 584960 112782
rect 182173 112162 182239 112165
rect 179860 112160 182239 112162
rect 179860 112104 182178 112160
rect 182234 112104 182239 112160
rect 179860 112102 182239 112104
rect 182173 112099 182239 112102
rect 117313 111482 117379 111485
rect 117313 111480 120060 111482
rect 117313 111424 117318 111480
rect 117374 111424 120060 111480
rect 117313 111422 120060 111424
rect 117313 111419 117379 111422
rect -960 110666 480 110756
rect 3141 110666 3207 110669
rect 183277 110666 183343 110669
rect -960 110664 3207 110666
rect -960 110608 3146 110664
rect 3202 110608 3207 110664
rect -960 110606 3207 110608
rect 179860 110664 183343 110666
rect 179860 110608 183282 110664
rect 183338 110608 183343 110664
rect 179860 110606 183343 110608
rect -960 110516 480 110606
rect 3141 110603 3207 110606
rect 183277 110603 183343 110606
rect 117313 109986 117379 109989
rect 117313 109984 120060 109986
rect 117313 109928 117318 109984
rect 117374 109928 120060 109984
rect 117313 109926 120060 109928
rect 117313 109923 117379 109926
rect 183461 109170 183527 109173
rect 179860 109168 183527 109170
rect 179860 109112 183466 109168
rect 183522 109112 183527 109168
rect 179860 109110 183527 109112
rect 183461 109107 183527 109110
rect 118417 108490 118483 108493
rect 118417 108488 120060 108490
rect 118417 108432 118422 108488
rect 118478 108432 120060 108488
rect 118417 108430 120060 108432
rect 118417 108427 118483 108430
rect 182265 107674 182331 107677
rect 179860 107672 182331 107674
rect 179860 107616 182270 107672
rect 182326 107616 182331 107672
rect 179860 107614 182331 107616
rect 182265 107611 182331 107614
rect 119337 106994 119403 106997
rect 119337 106992 120060 106994
rect 119337 106936 119342 106992
rect 119398 106936 120060 106992
rect 119337 106934 120060 106936
rect 119337 106931 119403 106934
rect 183461 106178 183527 106181
rect 179860 106176 183527 106178
rect 179860 106120 183466 106176
rect 183522 106120 183527 106176
rect 179860 106118 183527 106120
rect 183461 106115 183527 106118
rect 119245 105498 119311 105501
rect 119245 105496 120060 105498
rect 119245 105440 119250 105496
rect 119306 105440 120060 105496
rect 119245 105438 120060 105440
rect 119245 105435 119311 105438
rect 183461 104682 183527 104685
rect 179860 104680 183527 104682
rect 179860 104624 183466 104680
rect 183522 104624 183527 104680
rect 179860 104622 183527 104624
rect 183461 104619 183527 104622
rect 120625 104546 120691 104549
rect 120582 104544 120691 104546
rect 120582 104488 120630 104544
rect 120686 104488 120691 104544
rect 120582 104483 120691 104488
rect 120582 103972 120642 104483
rect 183461 103186 183527 103189
rect 179860 103184 183527 103186
rect 179860 103128 183466 103184
rect 183522 103128 183527 103184
rect 179860 103126 183527 103128
rect 183461 103123 183527 103126
rect 118785 102506 118851 102509
rect 118785 102504 120060 102506
rect 118785 102448 118790 102504
rect 118846 102448 120060 102504
rect 118785 102446 120060 102448
rect 118785 102443 118851 102446
rect 182909 101690 182975 101693
rect 179860 101688 182975 101690
rect 179860 101632 182914 101688
rect 182970 101632 182975 101688
rect 179860 101630 182975 101632
rect 182909 101627 182975 101630
rect 118877 101010 118943 101013
rect 118877 101008 120060 101010
rect 118877 100952 118882 101008
rect 118938 100952 120060 101008
rect 118877 100950 120060 100952
rect 118877 100947 118943 100950
rect 182909 100194 182975 100197
rect 179860 100192 182975 100194
rect 179860 100136 182914 100192
rect 182970 100136 182975 100192
rect 179860 100134 182975 100136
rect 182909 100131 182975 100134
rect 118969 99514 119035 99517
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 118969 99512 120060 99514
rect 118969 99456 118974 99512
rect 119030 99456 120060 99512
rect 118969 99454 120060 99456
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 118969 99451 119035 99454
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect 183093 98698 183159 98701
rect 179860 98696 183159 98698
rect 179860 98640 183098 98696
rect 183154 98640 183159 98696
rect 179860 98638 183159 98640
rect 183093 98635 183159 98638
rect 119153 98018 119219 98021
rect 119153 98016 120060 98018
rect 119153 97960 119158 98016
rect 119214 97960 120060 98016
rect 119153 97958 120060 97960
rect 119153 97955 119219 97958
rect -960 97610 480 97700
rect 3233 97610 3299 97613
rect -960 97608 3299 97610
rect -960 97552 3238 97608
rect 3294 97552 3299 97608
rect -960 97550 3299 97552
rect -960 97460 480 97550
rect 3233 97547 3299 97550
rect 183461 97202 183527 97205
rect 179860 97200 183527 97202
rect 179860 97144 183466 97200
rect 183522 97144 183527 97200
rect 179860 97142 183527 97144
rect 183461 97139 183527 97142
rect 119061 96522 119127 96525
rect 119061 96520 120060 96522
rect 119061 96464 119066 96520
rect 119122 96464 120060 96520
rect 119061 96462 120060 96464
rect 119061 96459 119127 96462
rect 183185 95706 183251 95709
rect 179860 95704 183251 95706
rect 179860 95648 183190 95704
rect 183246 95648 183251 95704
rect 179860 95646 183251 95648
rect 183185 95643 183251 95646
rect 118049 95026 118115 95029
rect 118049 95024 120060 95026
rect 118049 94968 118054 95024
rect 118110 94968 120060 95024
rect 118049 94966 120060 94968
rect 118049 94963 118115 94966
rect 183277 94210 183343 94213
rect 179860 94208 183343 94210
rect 179860 94152 183282 94208
rect 183338 94152 183343 94208
rect 179860 94150 183343 94152
rect 183277 94147 183343 94150
rect 118693 93530 118759 93533
rect 118693 93528 120060 93530
rect 118693 93472 118698 93528
rect 118754 93472 120060 93528
rect 118693 93470 120060 93472
rect 118693 93467 118759 93470
rect 183277 92714 183343 92717
rect 179860 92712 183343 92714
rect 179860 92656 183282 92712
rect 183338 92656 183343 92712
rect 179860 92654 183343 92656
rect 183277 92651 183343 92654
rect 118141 92034 118207 92037
rect 118141 92032 120060 92034
rect 118141 91976 118146 92032
rect 118202 91976 120060 92032
rect 118141 91974 120060 91976
rect 118141 91971 118207 91974
rect 183461 91218 183527 91221
rect 179860 91216 183527 91218
rect 179860 91160 183466 91216
rect 183522 91160 183527 91216
rect 179860 91158 183527 91160
rect 183461 91155 183527 91158
rect 118233 90538 118299 90541
rect 118233 90536 120060 90538
rect 118233 90480 118238 90536
rect 118294 90480 120060 90536
rect 118233 90478 120060 90480
rect 118233 90475 118299 90478
rect 182173 89722 182239 89725
rect 179860 89720 182239 89722
rect 179860 89664 182178 89720
rect 182234 89664 182239 89720
rect 179860 89662 182239 89664
rect 182173 89659 182239 89662
rect 118601 89042 118667 89045
rect 118601 89040 120060 89042
rect 118601 88984 118606 89040
rect 118662 88984 120060 89040
rect 118601 88982 120060 88984
rect 118601 88979 118667 88982
rect 180977 88226 181043 88229
rect 179860 88224 181043 88226
rect 179860 88168 180982 88224
rect 181038 88168 181043 88224
rect 179860 88166 181043 88168
rect 180977 88163 181043 88166
rect 118509 87546 118575 87549
rect 118509 87544 120060 87546
rect 118509 87488 118514 87544
rect 118570 87488 120060 87544
rect 118509 87486 120060 87488
rect 118509 87483 118575 87486
rect 182173 86730 182239 86733
rect 179860 86728 182239 86730
rect 179860 86672 182178 86728
rect 182234 86672 182239 86728
rect 179860 86670 182239 86672
rect 182173 86667 182239 86670
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 118325 86050 118391 86053
rect 118325 86048 120060 86050
rect 118325 85992 118330 86048
rect 118386 85992 120060 86048
rect 583520 86036 584960 86126
rect 118325 85990 120060 85992
rect 118325 85987 118391 85990
rect 182633 85234 182699 85237
rect 179860 85232 182699 85234
rect 179860 85176 182638 85232
rect 182694 85176 182699 85232
rect 179860 85174 182699 85176
rect 182633 85171 182699 85174
rect -960 84690 480 84780
rect 3969 84690 4035 84693
rect -960 84688 4035 84690
rect -960 84632 3974 84688
rect 4030 84632 4035 84688
rect -960 84630 4035 84632
rect -960 84540 480 84630
rect 3969 84627 4035 84630
rect 120582 84285 120642 84524
rect 120582 84280 120691 84285
rect 120582 84224 120630 84280
rect 120686 84224 120691 84280
rect 120582 84222 120691 84224
rect 120625 84219 120691 84222
rect 182817 83738 182883 83741
rect 179860 83736 182883 83738
rect 179860 83680 182822 83736
rect 182878 83680 182883 83736
rect 179860 83678 182883 83680
rect 182817 83675 182883 83678
rect 118509 83058 118575 83061
rect 118509 83056 120060 83058
rect 118509 83000 118514 83056
rect 118570 83000 120060 83056
rect 118509 82998 120060 83000
rect 118509 82995 118575 82998
rect 182449 82242 182515 82245
rect 179860 82240 182515 82242
rect 179860 82184 182454 82240
rect 182510 82184 182515 82240
rect 179860 82182 182515 82184
rect 182449 82179 182515 82182
rect 118417 81562 118483 81565
rect 118417 81560 120060 81562
rect 118417 81504 118422 81560
rect 118478 81504 120060 81560
rect 118417 81502 120060 81504
rect 118417 81499 118483 81502
rect 120625 81426 120691 81429
rect 180333 81426 180399 81429
rect 120625 81424 180399 81426
rect 120625 81368 120630 81424
rect 120686 81368 180338 81424
rect 180394 81368 180399 81424
rect 120625 81366 180399 81368
rect 120625 81363 120691 81366
rect 180333 81363 180399 81366
rect 3693 81290 3759 81293
rect 173566 81290 173572 81292
rect 3693 81288 173572 81290
rect 3693 81232 3698 81288
rect 3754 81232 173572 81288
rect 3693 81230 173572 81232
rect 3693 81227 3759 81230
rect 173566 81228 173572 81230
rect 173636 81228 173642 81292
rect 3509 81154 3575 81157
rect 3509 81152 150450 81154
rect 3509 81096 3514 81152
rect 3570 81096 150450 81152
rect 3509 81094 150450 81096
rect 3509 81091 3575 81094
rect 150390 80474 150450 81094
rect 171542 81092 171548 81156
rect 171612 81154 171618 81156
rect 180149 81154 180215 81157
rect 171612 81152 180215 81154
rect 171612 81096 180154 81152
rect 180210 81096 180215 81152
rect 171612 81094 180215 81096
rect 171612 81092 171618 81094
rect 180149 81091 180215 81094
rect 178493 81018 178559 81021
rect 396717 81018 396783 81021
rect 178493 81016 396783 81018
rect 178493 80960 178498 81016
rect 178554 80960 396722 81016
rect 396778 80960 396783 81016
rect 178493 80958 396783 80960
rect 178493 80955 178559 80958
rect 396717 80955 396783 80958
rect 178585 80882 178651 80885
rect 396901 80882 396967 80885
rect 178585 80880 396967 80882
rect 178585 80824 178590 80880
rect 178646 80824 396906 80880
rect 396962 80824 396967 80880
rect 178585 80822 396967 80824
rect 178585 80819 178651 80822
rect 396901 80819 396967 80822
rect 171174 80684 171180 80748
rect 171244 80746 171250 80748
rect 397085 80746 397151 80749
rect 171244 80744 397151 80746
rect 171244 80688 397090 80744
rect 397146 80688 397151 80744
rect 171244 80686 397151 80688
rect 171244 80684 171250 80686
rect 397085 80683 397151 80686
rect 166206 80548 166212 80612
rect 166276 80610 166282 80612
rect 171358 80610 171364 80612
rect 166276 80550 171364 80610
rect 166276 80548 166282 80550
rect 171358 80548 171364 80550
rect 171428 80548 171434 80612
rect 173198 80474 173204 80476
rect 150390 80414 173204 80474
rect 173198 80412 173204 80414
rect 173268 80412 173274 80476
rect 159038 80278 169770 80338
rect 131798 80140 131804 80204
rect 131868 80202 131874 80204
rect 131868 80142 132970 80202
rect 131868 80140 131874 80142
rect 132910 79967 132970 80142
rect 142838 80140 142844 80204
rect 142908 80202 142914 80204
rect 142908 80142 143458 80202
rect 142908 80140 142914 80142
rect 143398 79967 143458 80142
rect 159038 79967 159098 80278
rect 159214 80140 159220 80204
rect 159284 80202 159290 80204
rect 166206 80202 166212 80204
rect 159284 80142 166212 80202
rect 159284 80140 159290 80142
rect 166206 80140 166212 80142
rect 166276 80140 166282 80204
rect 169710 80202 169770 80278
rect 430573 80202 430639 80205
rect 169710 80200 430639 80202
rect 169710 80144 430578 80200
rect 430634 80144 430639 80200
rect 169710 80142 430639 80144
rect 430573 80139 430639 80142
rect 178493 80066 178559 80069
rect 171734 80064 178559 80066
rect 171734 80008 178498 80064
rect 178554 80008 178559 80064
rect 171734 80006 178559 80008
rect 126651 79962 126717 79967
rect 127663 79964 127729 79967
rect 125731 79932 125797 79933
rect 125726 79930 125732 79932
rect 125640 79870 125732 79930
rect 125726 79868 125732 79870
rect 125796 79868 125802 79932
rect 125910 79868 125916 79932
rect 125980 79930 125986 79932
rect 126191 79930 126257 79933
rect 125980 79928 126257 79930
rect 125980 79872 126196 79928
rect 126252 79872 126257 79928
rect 126651 79906 126656 79962
rect 126712 79906 126717 79962
rect 126651 79901 126717 79906
rect 127528 79962 127729 79964
rect 127528 79906 127668 79962
rect 127724 79906 127729 79962
rect 129963 79962 130029 79967
rect 127528 79904 127729 79906
rect 125980 79870 126257 79872
rect 125980 79868 125986 79870
rect 125731 79867 125797 79868
rect 126191 79867 126257 79870
rect 126513 79658 126579 79661
rect 126654 79658 126714 79901
rect 127203 79894 127269 79899
rect 127203 79838 127208 79894
rect 127264 79838 127269 79894
rect 127203 79833 127269 79838
rect 126513 79656 126714 79658
rect 126513 79600 126518 79656
rect 126574 79600 126714 79656
rect 126513 79598 126714 79600
rect 127065 79658 127131 79661
rect 127206 79658 127266 79833
rect 127528 79794 127588 79904
rect 127663 79901 127729 79904
rect 128123 79928 128189 79933
rect 128123 79872 128128 79928
rect 128184 79872 128189 79928
rect 128123 79867 128189 79872
rect 128486 79868 128492 79932
rect 128556 79930 128562 79932
rect 128767 79930 128833 79933
rect 129043 79932 129109 79933
rect 129038 79930 129044 79932
rect 128556 79928 128833 79930
rect 128556 79872 128772 79928
rect 128828 79872 128833 79928
rect 128556 79870 128833 79872
rect 128952 79870 129044 79930
rect 128556 79868 128562 79870
rect 128767 79867 128833 79870
rect 129038 79868 129044 79870
rect 129108 79868 129114 79932
rect 129411 79928 129477 79933
rect 129963 79932 129968 79962
rect 130024 79932 130029 79962
rect 131619 79962 131685 79967
rect 129411 79872 129416 79928
rect 129472 79872 129477 79928
rect 129043 79867 129109 79868
rect 129411 79867 129477 79872
rect 129779 79894 129845 79899
rect 127801 79794 127867 79797
rect 128126 79794 128186 79867
rect 127528 79792 127867 79794
rect 127528 79736 127806 79792
rect 127862 79736 127867 79792
rect 127528 79734 127867 79736
rect 127801 79731 127867 79734
rect 127942 79734 128186 79794
rect 128307 79792 128373 79797
rect 128307 79736 128312 79792
rect 128368 79736 128373 79792
rect 127065 79656 127266 79658
rect 127065 79600 127070 79656
rect 127126 79600 127266 79656
rect 127065 79598 127266 79600
rect 127341 79660 127407 79661
rect 127341 79656 127388 79660
rect 127452 79658 127458 79660
rect 127709 79658 127775 79661
rect 127942 79658 128002 79734
rect 128307 79731 128373 79736
rect 128997 79794 129063 79797
rect 129414 79794 129474 79867
rect 129779 79838 129784 79894
rect 129840 79838 129845 79894
rect 129958 79868 129964 79932
rect 130028 79930 130034 79932
rect 130028 79870 130086 79930
rect 130515 79928 130581 79933
rect 131619 79932 131624 79962
rect 131680 79932 131685 79962
rect 131895 79964 131961 79967
rect 131895 79962 132004 79964
rect 130515 79872 130520 79928
rect 130576 79872 130581 79928
rect 130028 79868 130034 79870
rect 130515 79867 130581 79872
rect 131614 79868 131620 79932
rect 131684 79930 131690 79932
rect 131684 79870 131742 79930
rect 131895 79906 131900 79962
rect 131956 79906 132004 79962
rect 132539 79962 132605 79967
rect 131895 79901 132004 79906
rect 131684 79868 131690 79870
rect 129779 79833 129845 79838
rect 128997 79792 129474 79794
rect 128997 79736 129002 79792
rect 129058 79736 129474 79792
rect 128997 79734 129474 79736
rect 128997 79731 129063 79734
rect 127341 79600 127346 79656
rect 126513 79595 126579 79598
rect 127065 79595 127131 79598
rect 127341 79596 127388 79600
rect 127452 79598 127498 79658
rect 127709 79656 128002 79658
rect 127709 79600 127714 79656
rect 127770 79600 128002 79656
rect 127709 79598 128002 79600
rect 128169 79658 128235 79661
rect 128310 79658 128370 79731
rect 128169 79656 128370 79658
rect 128169 79600 128174 79656
rect 128230 79600 128370 79656
rect 128169 79598 128370 79600
rect 128721 79658 128787 79661
rect 129782 79660 129842 79833
rect 130518 79797 130578 79867
rect 131343 79826 131409 79831
rect 130518 79792 130627 79797
rect 130518 79736 130566 79792
rect 130622 79736 130627 79792
rect 130518 79734 130627 79736
rect 130561 79731 130627 79734
rect 130878 79732 130884 79796
rect 130948 79794 130954 79796
rect 131343 79794 131348 79826
rect 130948 79770 131348 79794
rect 131404 79770 131409 79826
rect 130948 79765 131409 79770
rect 131573 79794 131639 79797
rect 131944 79794 132004 79901
rect 132355 79928 132421 79933
rect 132355 79872 132360 79928
rect 132416 79872 132421 79928
rect 132539 79906 132544 79962
rect 132600 79906 132605 79962
rect 132907 79962 132973 79967
rect 132539 79901 132605 79906
rect 132723 79930 132789 79933
rect 132723 79928 132832 79930
rect 132355 79867 132421 79872
rect 131573 79792 132004 79794
rect 130948 79734 131406 79765
rect 131573 79736 131578 79792
rect 131634 79736 132004 79792
rect 131573 79734 132004 79736
rect 130948 79732 130954 79734
rect 131573 79731 131639 79734
rect 128854 79658 128860 79660
rect 128721 79656 128860 79658
rect 128721 79600 128726 79656
rect 128782 79600 128860 79656
rect 128721 79598 128860 79600
rect 127452 79596 127458 79598
rect 127341 79595 127407 79596
rect 127709 79595 127775 79598
rect 128169 79595 128235 79598
rect 128721 79595 128787 79598
rect 128854 79596 128860 79598
rect 128924 79596 128930 79660
rect 129774 79596 129780 79660
rect 129844 79596 129850 79660
rect 132217 79658 132283 79661
rect 132358 79658 132418 79867
rect 132542 79661 132602 79901
rect 132723 79872 132728 79928
rect 132784 79872 132832 79928
rect 132907 79906 132912 79962
rect 132968 79906 132973 79962
rect 134471 79964 134537 79967
rect 134471 79962 134580 79964
rect 132907 79901 132973 79906
rect 132723 79867 132832 79872
rect 133454 79868 133460 79932
rect 133524 79930 133530 79932
rect 133735 79930 133801 79933
rect 134011 79932 134077 79933
rect 134006 79930 134012 79932
rect 133524 79928 133801 79930
rect 133524 79872 133740 79928
rect 133796 79872 133801 79928
rect 133524 79870 133801 79872
rect 133920 79870 134012 79930
rect 133524 79868 133530 79870
rect 133735 79867 133801 79870
rect 134006 79868 134012 79870
rect 134076 79868 134082 79932
rect 134287 79930 134353 79933
rect 134152 79928 134353 79930
rect 134152 79872 134292 79928
rect 134348 79872 134353 79928
rect 134471 79906 134476 79962
rect 134532 79932 134580 79962
rect 135851 79962 135917 79967
rect 134532 79906 134564 79932
rect 134471 79901 134564 79906
rect 134152 79870 134353 79872
rect 134520 79870 134564 79901
rect 134011 79867 134077 79868
rect 132772 79794 132832 79867
rect 133086 79794 133092 79796
rect 132772 79734 133092 79794
rect 133086 79732 133092 79734
rect 133156 79732 133162 79796
rect 133270 79732 133276 79796
rect 133340 79794 133346 79796
rect 134152 79794 134212 79870
rect 134287 79867 134353 79870
rect 134558 79868 134564 79870
rect 134628 79868 134634 79932
rect 134931 79928 134997 79933
rect 135483 79932 135549 79933
rect 134931 79872 134936 79928
rect 134992 79872 134997 79928
rect 134931 79867 134997 79872
rect 135478 79868 135484 79932
rect 135548 79930 135554 79932
rect 135548 79870 135640 79930
rect 135851 79906 135856 79962
rect 135912 79906 135917 79962
rect 136403 79962 136469 79967
rect 136403 79932 136408 79962
rect 136464 79932 136469 79962
rect 136587 79962 136653 79967
rect 137047 79964 137113 79967
rect 135851 79901 135917 79906
rect 135548 79868 135554 79870
rect 135483 79867 135549 79868
rect 133340 79734 134212 79794
rect 133340 79732 133346 79734
rect 132217 79656 132418 79658
rect 132217 79600 132222 79656
rect 132278 79600 132418 79656
rect 132217 79598 132418 79600
rect 132493 79656 132602 79661
rect 132493 79600 132498 79656
rect 132554 79600 132602 79656
rect 132493 79598 132602 79600
rect 132769 79658 132835 79661
rect 134934 79658 134994 79867
rect 132769 79656 134994 79658
rect 132769 79600 132774 79656
rect 132830 79600 134994 79656
rect 132769 79598 134994 79600
rect 135621 79658 135687 79661
rect 135854 79658 135914 79901
rect 136398 79868 136404 79932
rect 136468 79930 136474 79932
rect 136468 79870 136526 79930
rect 136587 79906 136592 79962
rect 136648 79906 136653 79962
rect 137004 79962 137113 79964
rect 137004 79932 137052 79962
rect 136587 79901 136653 79906
rect 136468 79868 136474 79870
rect 136590 79797 136650 79901
rect 136950 79868 136956 79932
rect 137020 79906 137052 79932
rect 137108 79906 137113 79962
rect 137020 79901 137113 79906
rect 137691 79962 137757 79967
rect 137691 79906 137696 79962
rect 137752 79930 137757 79962
rect 138243 79962 138309 79967
rect 138054 79930 138060 79932
rect 137752 79906 138060 79930
rect 137691 79901 138060 79906
rect 137020 79870 137064 79901
rect 137694 79870 138060 79901
rect 137020 79868 137026 79870
rect 138054 79868 138060 79870
rect 138124 79868 138130 79932
rect 138243 79906 138248 79962
rect 138304 79906 138309 79962
rect 138243 79901 138309 79906
rect 138611 79962 138677 79967
rect 138611 79906 138616 79962
rect 138672 79906 138677 79962
rect 138611 79901 138677 79906
rect 139347 79962 139413 79967
rect 140543 79964 140609 79967
rect 139347 79906 139352 79962
rect 139408 79906 139413 79962
rect 140500 79962 140609 79964
rect 139531 79930 139597 79933
rect 139347 79901 139413 79906
rect 139488 79928 139597 79930
rect 136541 79792 136650 79797
rect 136541 79736 136546 79792
rect 136602 79736 136650 79792
rect 136541 79734 136650 79736
rect 136541 79731 136607 79734
rect 138246 79661 138306 79901
rect 135621 79656 135914 79658
rect 135621 79600 135626 79656
rect 135682 79600 135914 79656
rect 135621 79598 135914 79600
rect 138197 79656 138306 79661
rect 138197 79600 138202 79656
rect 138258 79600 138306 79656
rect 138197 79598 138306 79600
rect 138614 79658 138674 79901
rect 139350 79797 139410 79901
rect 139488 79872 139536 79928
rect 139592 79872 139597 79928
rect 139488 79867 139597 79872
rect 139715 79928 139781 79933
rect 139715 79872 139720 79928
rect 139776 79872 139781 79928
rect 139715 79867 139781 79872
rect 140262 79868 140268 79932
rect 140332 79930 140338 79932
rect 140500 79930 140548 79962
rect 140332 79906 140548 79930
rect 140604 79906 140609 79962
rect 143395 79962 143461 79967
rect 140332 79901 140609 79906
rect 141279 79930 141345 79933
rect 141831 79930 141897 79933
rect 142751 79930 142817 79933
rect 141279 79928 141480 79930
rect 140332 79870 140560 79901
rect 141279 79872 141284 79928
rect 141340 79872 141480 79928
rect 141279 79870 141480 79872
rect 140332 79868 140338 79870
rect 141279 79867 141345 79870
rect 139488 79797 139548 79867
rect 138790 79732 138796 79796
rect 138860 79794 138866 79796
rect 138979 79794 139045 79797
rect 138860 79792 139045 79794
rect 138860 79736 138984 79792
rect 139040 79736 139045 79792
rect 138860 79734 139045 79736
rect 138860 79732 138866 79734
rect 138979 79731 139045 79734
rect 139117 79796 139183 79797
rect 139117 79792 139164 79796
rect 139228 79794 139234 79796
rect 139117 79736 139122 79792
rect 139117 79732 139164 79736
rect 139228 79734 139274 79794
rect 139347 79792 139413 79797
rect 139347 79736 139352 79792
rect 139408 79736 139413 79792
rect 139228 79732 139234 79734
rect 139117 79731 139183 79732
rect 139347 79731 139413 79736
rect 139485 79792 139551 79797
rect 139485 79736 139490 79792
rect 139546 79736 139551 79792
rect 139485 79731 139551 79736
rect 138933 79658 138999 79661
rect 138614 79656 138999 79658
rect 138614 79600 138938 79656
rect 138994 79600 138999 79656
rect 138614 79598 138999 79600
rect 139718 79658 139778 79867
rect 140078 79732 140084 79796
rect 140148 79794 140154 79796
rect 140451 79794 140517 79797
rect 140148 79792 140517 79794
rect 140148 79736 140456 79792
rect 140512 79736 140517 79792
rect 140148 79734 140517 79736
rect 140148 79732 140154 79734
rect 140451 79731 140517 79734
rect 141233 79794 141299 79797
rect 141420 79794 141480 79870
rect 141831 79928 142032 79930
rect 141831 79872 141836 79928
rect 141892 79872 142032 79928
rect 141831 79870 142032 79872
rect 141831 79867 141897 79870
rect 141233 79792 141480 79794
rect 141233 79736 141238 79792
rect 141294 79736 141480 79792
rect 141233 79734 141480 79736
rect 141233 79731 141299 79734
rect 141972 79661 142032 79870
rect 142751 79928 142860 79930
rect 142751 79872 142756 79928
rect 142812 79872 142860 79928
rect 143395 79906 143400 79962
rect 143456 79906 143461 79962
rect 144867 79962 144933 79967
rect 143855 79930 143921 79933
rect 143395 79901 143461 79906
rect 143582 79928 143921 79930
rect 142751 79867 142860 79872
rect 142800 79797 142860 79867
rect 143582 79872 143860 79928
rect 143916 79872 143921 79928
rect 143582 79870 143921 79872
rect 142751 79792 142860 79797
rect 142751 79736 142756 79792
rect 142812 79736 142860 79792
rect 143119 79828 143185 79831
rect 143119 79826 143228 79828
rect 143119 79770 143124 79826
rect 143180 79770 143228 79826
rect 143119 79765 143228 79770
rect 142751 79734 142860 79736
rect 142751 79731 142817 79734
rect 143168 79661 143228 79765
rect 143582 79797 143642 79870
rect 143855 79867 143921 79870
rect 144494 79868 144500 79932
rect 144564 79930 144570 79932
rect 144867 79930 144872 79962
rect 144564 79906 144872 79930
rect 144928 79906 144933 79962
rect 144564 79901 144933 79906
rect 145051 79962 145117 79967
rect 145051 79906 145056 79962
rect 145112 79906 145117 79962
rect 146707 79962 146773 79967
rect 145051 79901 145117 79906
rect 144564 79870 144930 79901
rect 144564 79868 144570 79870
rect 145054 79797 145114 79901
rect 145598 79868 145604 79932
rect 145668 79930 145674 79932
rect 146155 79930 146221 79933
rect 145668 79928 146221 79930
rect 145668 79872 146160 79928
rect 146216 79872 146221 79928
rect 145668 79870 146221 79872
rect 145668 79868 145674 79870
rect 146155 79867 146221 79870
rect 146339 79928 146405 79933
rect 146707 79932 146712 79962
rect 146768 79932 146773 79962
rect 148915 79962 148981 79967
rect 147075 79932 147141 79933
rect 147811 79932 147877 79933
rect 146339 79872 146344 79928
rect 146400 79872 146405 79928
rect 146339 79867 146405 79872
rect 146702 79868 146708 79932
rect 146772 79930 146778 79932
rect 146772 79870 146830 79930
rect 146772 79868 146778 79870
rect 147070 79868 147076 79932
rect 147140 79930 147146 79932
rect 147806 79930 147812 79932
rect 147140 79870 147232 79930
rect 147720 79870 147812 79930
rect 147140 79868 147146 79870
rect 147806 79868 147812 79870
rect 147876 79868 147882 79932
rect 148639 79928 148705 79933
rect 148915 79932 148920 79962
rect 148976 79932 148981 79962
rect 150295 79962 150361 79967
rect 148639 79872 148644 79928
rect 148700 79872 148705 79928
rect 147075 79867 147141 79868
rect 147811 79867 147877 79868
rect 148639 79867 148705 79872
rect 148910 79868 148916 79932
rect 148980 79930 148986 79932
rect 149191 79930 149257 79933
rect 148980 79870 149038 79930
rect 149191 79928 149530 79930
rect 149191 79872 149196 79928
rect 149252 79872 149530 79928
rect 149191 79870 149530 79872
rect 148980 79868 148986 79870
rect 149191 79867 149257 79870
rect 143582 79792 143691 79797
rect 143582 79736 143630 79792
rect 143686 79736 143691 79792
rect 143582 79734 143691 79736
rect 143625 79731 143691 79734
rect 145005 79792 145114 79797
rect 145005 79736 145010 79792
rect 145066 79736 145114 79792
rect 145005 79734 145114 79736
rect 145005 79731 145071 79734
rect 141141 79658 141207 79661
rect 139718 79656 141207 79658
rect 139718 79600 141146 79656
rect 141202 79600 141207 79656
rect 139718 79598 141207 79600
rect 132217 79595 132283 79598
rect 132493 79595 132559 79598
rect 132769 79595 132835 79598
rect 135621 79595 135687 79598
rect 138197 79595 138263 79598
rect 138933 79595 138999 79598
rect 141141 79595 141207 79598
rect 141969 79656 142035 79661
rect 141969 79600 141974 79656
rect 142030 79600 142035 79656
rect 141969 79595 142035 79600
rect 143165 79656 143231 79661
rect 143165 79600 143170 79656
rect 143226 79600 143231 79656
rect 143165 79595 143231 79600
rect 144310 79596 144316 79660
rect 144380 79658 144386 79660
rect 144453 79658 144519 79661
rect 146201 79660 146267 79661
rect 146150 79658 146156 79660
rect 144380 79656 144519 79658
rect 144380 79600 144458 79656
rect 144514 79600 144519 79656
rect 144380 79598 144519 79600
rect 146110 79598 146156 79658
rect 146220 79656 146267 79660
rect 146262 79600 146267 79656
rect 144380 79596 144386 79598
rect 144453 79595 144519 79598
rect 146150 79596 146156 79598
rect 146220 79596 146267 79600
rect 146342 79658 146402 79867
rect 147765 79658 147831 79661
rect 146342 79656 147831 79658
rect 146342 79600 147770 79656
rect 147826 79600 147831 79656
rect 146342 79598 147831 79600
rect 148642 79658 148702 79867
rect 149145 79794 149211 79797
rect 149470 79794 149530 79870
rect 149646 79868 149652 79932
rect 149716 79930 149722 79932
rect 150295 79930 150300 79962
rect 149716 79906 150300 79930
rect 150356 79906 150361 79962
rect 153147 79962 153213 79967
rect 149716 79901 150361 79906
rect 150755 79928 150821 79933
rect 149716 79870 150358 79901
rect 150755 79872 150760 79928
rect 150816 79872 150821 79928
rect 149716 79868 149722 79870
rect 150755 79867 150821 79872
rect 151399 79930 151465 79933
rect 151670 79930 151676 79932
rect 151399 79928 151676 79930
rect 151399 79872 151404 79928
rect 151460 79872 151676 79928
rect 151399 79870 151676 79872
rect 151399 79867 151465 79870
rect 151670 79868 151676 79870
rect 151740 79868 151746 79932
rect 151951 79930 152017 79933
rect 151951 79928 152290 79930
rect 151951 79872 151956 79928
rect 152012 79872 152290 79928
rect 151951 79870 152290 79872
rect 151951 79867 152017 79870
rect 149145 79792 149530 79794
rect 149145 79736 149150 79792
rect 149206 79736 149530 79792
rect 149145 79734 149530 79736
rect 149145 79731 149211 79734
rect 149830 79732 149836 79796
rect 149900 79794 149906 79796
rect 150111 79794 150177 79797
rect 149900 79792 150177 79794
rect 149900 79736 150116 79792
rect 150172 79736 150177 79792
rect 149900 79734 150177 79736
rect 149900 79732 149906 79734
rect 150111 79731 150177 79734
rect 148869 79658 148935 79661
rect 148642 79656 148935 79658
rect 148642 79600 148874 79656
rect 148930 79600 148935 79656
rect 148642 79598 148935 79600
rect 150758 79658 150818 79867
rect 151486 79732 151492 79796
rect 151556 79794 151562 79796
rect 151767 79794 151833 79797
rect 151556 79792 151833 79794
rect 151556 79736 151772 79792
rect 151828 79736 151833 79792
rect 151556 79734 151833 79736
rect 151556 79732 151562 79734
rect 151767 79731 151833 79734
rect 151997 79794 152063 79797
rect 152230 79794 152290 79870
rect 152595 79928 152661 79933
rect 152779 79932 152845 79933
rect 152595 79872 152600 79928
rect 152656 79872 152661 79928
rect 152595 79867 152661 79872
rect 152774 79868 152780 79932
rect 152844 79930 152850 79932
rect 152844 79870 152936 79930
rect 153147 79906 153152 79962
rect 153208 79930 153213 79962
rect 159035 79962 159101 79967
rect 153208 79906 153394 79930
rect 153147 79901 153394 79906
rect 153150 79870 153394 79901
rect 152844 79868 152850 79870
rect 152779 79867 152845 79868
rect 151997 79792 152290 79794
rect 151997 79736 152002 79792
rect 152058 79736 152290 79792
rect 151997 79734 152290 79736
rect 152598 79794 152658 79867
rect 153101 79794 153167 79797
rect 152598 79792 153167 79794
rect 152598 79736 153106 79792
rect 153162 79736 153167 79792
rect 152598 79734 153167 79736
rect 151997 79731 152063 79734
rect 153101 79731 153167 79734
rect 152457 79658 152523 79661
rect 150758 79656 152523 79658
rect 150758 79600 152462 79656
rect 152518 79600 152523 79656
rect 150758 79598 152523 79600
rect 146201 79595 146267 79596
rect 147765 79595 147831 79598
rect 148869 79595 148935 79598
rect 152457 79595 152523 79598
rect 153193 79658 153259 79661
rect 153334 79658 153394 79870
rect 153699 79928 153765 79933
rect 154067 79932 154133 79933
rect 154062 79930 154068 79932
rect 153699 79872 153704 79928
rect 153760 79872 153765 79928
rect 153699 79867 153765 79872
rect 153976 79870 154068 79930
rect 154062 79868 154068 79870
rect 154132 79868 154138 79932
rect 154246 79868 154252 79932
rect 154316 79930 154322 79932
rect 154435 79930 154501 79933
rect 154316 79928 154501 79930
rect 154316 79872 154440 79928
rect 154496 79872 154501 79928
rect 154316 79870 154501 79872
rect 154316 79868 154322 79870
rect 154067 79867 154133 79868
rect 154435 79867 154501 79870
rect 154711 79930 154777 79933
rect 154982 79930 154988 79932
rect 154711 79928 154988 79930
rect 154711 79872 154716 79928
rect 154772 79872 154988 79928
rect 154711 79870 154988 79872
rect 154711 79867 154777 79870
rect 154982 79868 154988 79870
rect 155052 79868 155058 79932
rect 155447 79930 155513 79933
rect 155723 79932 155789 79933
rect 156091 79932 156157 79933
rect 155718 79930 155724 79932
rect 155174 79928 155513 79930
rect 155174 79872 155452 79928
rect 155508 79872 155513 79928
rect 155174 79870 155513 79872
rect 155632 79870 155724 79930
rect 153193 79656 153394 79658
rect 153193 79600 153198 79656
rect 153254 79600 153394 79656
rect 153193 79598 153394 79600
rect 153702 79658 153762 79867
rect 153878 79732 153884 79796
rect 153948 79794 153954 79796
rect 154159 79794 154225 79797
rect 153948 79792 154225 79794
rect 153948 79736 154164 79792
rect 154220 79736 154225 79792
rect 153948 79734 154225 79736
rect 155174 79794 155234 79870
rect 155447 79867 155513 79870
rect 155718 79868 155724 79870
rect 155788 79868 155794 79932
rect 156086 79930 156092 79932
rect 156000 79870 156092 79930
rect 156086 79868 156092 79870
rect 156156 79868 156162 79932
rect 156551 79930 156617 79933
rect 156278 79928 156617 79930
rect 156278 79872 156556 79928
rect 156612 79872 156617 79928
rect 156278 79870 156617 79872
rect 155723 79867 155789 79868
rect 156091 79867 156157 79868
rect 155401 79794 155467 79797
rect 155174 79792 155467 79794
rect 155174 79736 155406 79792
rect 155462 79736 155467 79792
rect 155174 79734 155467 79736
rect 153948 79732 153954 79734
rect 154159 79731 154225 79734
rect 155401 79731 155467 79734
rect 154573 79658 154639 79661
rect 153702 79656 154639 79658
rect 153702 79600 154578 79656
rect 154634 79600 154639 79656
rect 153702 79598 154639 79600
rect 156278 79658 156338 79870
rect 156551 79867 156617 79870
rect 156822 79868 156828 79932
rect 156892 79930 156898 79932
rect 157103 79930 157169 79933
rect 157747 79932 157813 79933
rect 157742 79930 157748 79932
rect 156892 79928 157169 79930
rect 156892 79872 157108 79928
rect 157164 79872 157169 79928
rect 156892 79870 157169 79872
rect 157656 79870 157748 79930
rect 156892 79868 156898 79870
rect 157103 79867 157169 79870
rect 157742 79868 157748 79870
rect 157812 79868 157818 79932
rect 158110 79868 158116 79932
rect 158180 79930 158186 79932
rect 158483 79930 158549 79933
rect 158180 79928 158549 79930
rect 158180 79872 158488 79928
rect 158544 79872 158549 79928
rect 159035 79906 159040 79962
rect 159096 79906 159101 79962
rect 160691 79962 160757 79967
rect 159035 79901 159101 79906
rect 159955 79928 160021 79933
rect 158180 79870 158549 79872
rect 158180 79868 158186 79870
rect 157747 79867 157813 79868
rect 158483 79867 158549 79870
rect 159955 79872 159960 79928
rect 160016 79872 160021 79928
rect 160691 79906 160696 79962
rect 160752 79906 160757 79962
rect 167499 79962 167565 79967
rect 160691 79901 160757 79906
rect 160875 79928 160941 79933
rect 161243 79932 161309 79933
rect 161238 79930 161244 79932
rect 159955 79867 160021 79872
rect 156505 79794 156571 79797
rect 156505 79792 156890 79794
rect 156505 79736 156510 79792
rect 156566 79736 156890 79792
rect 156505 79734 156890 79736
rect 156505 79731 156571 79734
rect 156413 79658 156479 79661
rect 156278 79656 156479 79658
rect 156278 79600 156418 79656
rect 156474 79600 156479 79656
rect 156278 79598 156479 79600
rect 156830 79658 156890 79734
rect 157006 79732 157012 79796
rect 157076 79794 157082 79796
rect 157195 79794 157261 79797
rect 158299 79796 158365 79797
rect 158294 79794 158300 79796
rect 157076 79792 157261 79794
rect 157076 79736 157200 79792
rect 157256 79736 157261 79792
rect 157076 79734 157261 79736
rect 158208 79734 158300 79794
rect 157076 79732 157082 79734
rect 157195 79731 157261 79734
rect 158294 79732 158300 79734
rect 158364 79732 158370 79796
rect 159030 79732 159036 79796
rect 159100 79794 159106 79796
rect 159958 79794 160018 79867
rect 159100 79734 160018 79794
rect 159100 79732 159106 79734
rect 158299 79731 158365 79732
rect 160694 79661 160754 79901
rect 160875 79872 160880 79928
rect 160936 79872 160941 79928
rect 160875 79867 160941 79872
rect 161152 79870 161244 79930
rect 161238 79868 161244 79870
rect 161308 79868 161314 79932
rect 161611 79928 161677 79933
rect 161611 79872 161616 79928
rect 161672 79872 161677 79928
rect 161243 79867 161309 79868
rect 161611 79867 161677 79872
rect 162439 79930 162505 79933
rect 162710 79930 162716 79932
rect 162439 79928 162716 79930
rect 162439 79872 162444 79928
rect 162500 79872 162716 79928
rect 162439 79870 162716 79872
rect 162439 79867 162505 79870
rect 162710 79868 162716 79870
rect 162780 79868 162786 79932
rect 163267 79928 163333 79933
rect 163267 79872 163272 79928
rect 163328 79872 163333 79928
rect 163267 79867 163333 79872
rect 163446 79868 163452 79932
rect 163516 79930 163522 79932
rect 164003 79930 164069 79933
rect 163516 79928 164069 79930
rect 163516 79872 164008 79928
rect 164064 79872 164069 79928
rect 163516 79870 164069 79872
rect 163516 79868 163522 79870
rect 164003 79867 164069 79870
rect 164555 79928 164621 79933
rect 164923 79932 164989 79933
rect 164918 79930 164924 79932
rect 164555 79872 164560 79928
rect 164616 79872 164621 79928
rect 164555 79867 164621 79872
rect 164832 79870 164924 79930
rect 164918 79868 164924 79870
rect 164988 79868 164994 79932
rect 165102 79868 165108 79932
rect 165172 79930 165178 79932
rect 165567 79930 165633 79933
rect 165172 79928 165633 79930
rect 165172 79872 165572 79928
rect 165628 79872 165633 79928
rect 165172 79870 165633 79872
rect 165172 79868 165178 79870
rect 164923 79867 164989 79868
rect 165567 79867 165633 79870
rect 165935 79930 166001 79933
rect 165935 79928 166274 79930
rect 165935 79872 165940 79928
rect 165996 79872 166274 79928
rect 165935 79870 166274 79872
rect 165935 79867 166001 79870
rect 158253 79658 158319 79661
rect 156830 79656 158319 79658
rect 156830 79600 158258 79656
rect 158314 79600 158319 79656
rect 156830 79598 158319 79600
rect 153193 79595 153259 79598
rect 154573 79595 154639 79598
rect 156413 79595 156479 79598
rect 158253 79595 158319 79598
rect 158989 79658 159055 79661
rect 159909 79658 159975 79661
rect 158989 79656 159975 79658
rect 158989 79600 158994 79656
rect 159050 79600 159914 79656
rect 159970 79600 159975 79656
rect 158989 79598 159975 79600
rect 158989 79595 159055 79598
rect 159909 79595 159975 79598
rect 160134 79596 160140 79660
rect 160204 79658 160210 79660
rect 160369 79658 160435 79661
rect 160204 79656 160435 79658
rect 160204 79600 160374 79656
rect 160430 79600 160435 79656
rect 160204 79598 160435 79600
rect 160694 79656 160803 79661
rect 160694 79600 160742 79656
rect 160798 79600 160803 79656
rect 160694 79598 160803 79600
rect 160878 79658 160938 79867
rect 161614 79794 161674 79867
rect 163270 79797 163330 79867
rect 161933 79794 161999 79797
rect 161614 79792 161999 79794
rect 161614 79736 161938 79792
rect 161994 79736 161999 79792
rect 161614 79734 161999 79736
rect 161933 79731 161999 79734
rect 162342 79732 162348 79796
rect 162412 79794 162418 79796
rect 162623 79794 162689 79797
rect 162412 79792 162689 79794
rect 162412 79736 162628 79792
rect 162684 79736 162689 79792
rect 162412 79734 162689 79736
rect 162412 79732 162418 79734
rect 162623 79731 162689 79734
rect 162899 79792 162965 79797
rect 162899 79736 162904 79792
rect 162960 79736 162965 79792
rect 162899 79731 162965 79736
rect 163270 79792 163379 79797
rect 163270 79736 163318 79792
rect 163374 79736 163379 79792
rect 163270 79734 163379 79736
rect 163313 79731 163379 79734
rect 162209 79658 162275 79661
rect 160878 79656 162275 79658
rect 160878 79600 162214 79656
rect 162270 79600 162275 79656
rect 160878 79598 162275 79600
rect 160204 79596 160210 79598
rect 160369 79595 160435 79598
rect 160737 79595 160803 79598
rect 162209 79595 162275 79598
rect 162526 79596 162532 79660
rect 162596 79658 162602 79660
rect 162669 79658 162735 79661
rect 162596 79656 162735 79658
rect 162596 79600 162674 79656
rect 162730 79600 162735 79656
rect 162596 79598 162735 79600
rect 162902 79658 162962 79731
rect 163957 79658 164023 79661
rect 162902 79656 164023 79658
rect 162902 79600 163962 79656
rect 164018 79600 164023 79656
rect 162902 79598 164023 79600
rect 162596 79596 162602 79598
rect 162669 79595 162735 79598
rect 163957 79595 164023 79598
rect 164141 79658 164207 79661
rect 164366 79658 164372 79660
rect 164141 79656 164372 79658
rect 164141 79600 164146 79656
rect 164202 79600 164372 79656
rect 164141 79598 164372 79600
rect 164141 79595 164207 79598
rect 164366 79596 164372 79598
rect 164436 79596 164442 79660
rect 164558 79658 164618 79867
rect 165291 79796 165357 79797
rect 165286 79794 165292 79796
rect 165200 79734 165292 79794
rect 165286 79732 165292 79734
rect 165356 79732 165362 79796
rect 165889 79794 165955 79797
rect 165889 79792 166090 79794
rect 165889 79736 165894 79792
rect 165950 79736 166090 79792
rect 165889 79734 166090 79736
rect 165291 79731 165357 79732
rect 165889 79731 165955 79734
rect 166030 79661 166090 79734
rect 165245 79658 165311 79661
rect 164558 79656 165311 79658
rect 164558 79600 165250 79656
rect 165306 79600 165311 79656
rect 164558 79598 165311 79600
rect 166030 79656 166139 79661
rect 166030 79600 166078 79656
rect 166134 79600 166139 79656
rect 166030 79598 166139 79600
rect 166214 79658 166274 79870
rect 166390 79868 166396 79932
rect 166460 79930 166466 79932
rect 166763 79930 166829 79933
rect 166460 79928 166829 79930
rect 166460 79872 166768 79928
rect 166824 79872 166829 79928
rect 166460 79870 166829 79872
rect 166460 79868 166466 79870
rect 166763 79867 166829 79870
rect 167131 79928 167197 79933
rect 167131 79872 167136 79928
rect 167192 79872 167197 79928
rect 167131 79867 167197 79872
rect 167315 79928 167381 79933
rect 167499 79932 167504 79962
rect 167560 79932 167565 79962
rect 168419 79962 168485 79967
rect 167315 79872 167320 79928
rect 167376 79872 167381 79928
rect 167315 79867 167381 79872
rect 167494 79868 167500 79932
rect 167564 79930 167570 79932
rect 167564 79870 167622 79930
rect 168419 79906 168424 79962
rect 168480 79930 168485 79962
rect 171734 79933 171794 80006
rect 178493 80003 178559 80006
rect 169339 79932 169405 79933
rect 169150 79930 169156 79932
rect 168480 79906 169156 79930
rect 168419 79901 169156 79906
rect 168422 79870 169156 79901
rect 167564 79868 167570 79870
rect 169150 79868 169156 79870
rect 169220 79868 169226 79932
rect 169334 79868 169340 79932
rect 169404 79930 169410 79932
rect 169983 79930 170049 79933
rect 169404 79870 169496 79930
rect 169710 79928 170049 79930
rect 169710 79872 169988 79928
rect 170044 79872 170049 79928
rect 169710 79870 170049 79872
rect 169404 79868 169410 79870
rect 169339 79867 169405 79868
rect 166574 79732 166580 79796
rect 166644 79794 166650 79796
rect 166947 79794 167013 79797
rect 166644 79792 167013 79794
rect 166644 79736 166952 79792
rect 167008 79736 167013 79792
rect 166644 79734 167013 79736
rect 166644 79732 166650 79734
rect 166947 79731 167013 79734
rect 167134 79661 167194 79867
rect 167318 79794 167378 79867
rect 168557 79794 168623 79797
rect 167318 79792 168623 79794
rect 167318 79736 168562 79792
rect 168618 79736 168623 79792
rect 167318 79734 168623 79736
rect 168557 79731 168623 79734
rect 166625 79658 166691 79661
rect 166214 79656 166691 79658
rect 166214 79600 166630 79656
rect 166686 79600 166691 79656
rect 166214 79598 166691 79600
rect 167134 79656 167243 79661
rect 167134 79600 167182 79656
rect 167238 79600 167243 79656
rect 167134 79598 167243 79600
rect 165245 79595 165311 79598
rect 166073 79595 166139 79598
rect 166625 79595 166691 79598
rect 167177 79595 167243 79598
rect 167862 79596 167868 79660
rect 167932 79658 167938 79660
rect 168281 79658 168347 79661
rect 167932 79656 168347 79658
rect 167932 79600 168286 79656
rect 168342 79600 168347 79656
rect 167932 79598 168347 79600
rect 169710 79658 169770 79870
rect 169983 79867 170049 79870
rect 170438 79868 170444 79932
rect 170508 79930 170514 79932
rect 170811 79930 170877 79933
rect 170508 79928 170877 79930
rect 170508 79872 170816 79928
rect 170872 79872 170877 79928
rect 170508 79870 170877 79872
rect 170508 79868 170514 79870
rect 170811 79867 170877 79870
rect 171174 79868 171180 79932
rect 171244 79930 171250 79932
rect 171547 79930 171613 79933
rect 171244 79928 171613 79930
rect 171244 79872 171552 79928
rect 171608 79872 171613 79928
rect 171244 79870 171613 79872
rect 171244 79868 171250 79870
rect 171547 79867 171613 79870
rect 171731 79928 171797 79933
rect 171915 79932 171981 79933
rect 172375 79932 172441 79933
rect 171731 79872 171736 79928
rect 171792 79872 171797 79928
rect 171731 79867 171797 79872
rect 171910 79868 171916 79932
rect 171980 79930 171986 79932
rect 172375 79930 172422 79932
rect 171980 79870 172072 79930
rect 172330 79928 172422 79930
rect 172330 79872 172380 79928
rect 172330 79870 172422 79872
rect 171980 79868 171986 79870
rect 172375 79868 172422 79870
rect 172486 79868 172492 79932
rect 172559 79930 172625 79933
rect 176653 79930 176719 79933
rect 172559 79928 176719 79930
rect 172559 79872 172564 79928
rect 172620 79872 176658 79928
rect 176714 79872 176719 79928
rect 172559 79870 176719 79872
rect 171915 79867 171981 79868
rect 172375 79867 172441 79868
rect 172559 79867 172625 79870
rect 176653 79867 176719 79870
rect 170259 79794 170325 79797
rect 170581 79794 170647 79797
rect 170259 79792 170647 79794
rect 170259 79736 170264 79792
rect 170320 79736 170586 79792
rect 170642 79736 170647 79792
rect 170259 79734 170647 79736
rect 170259 79731 170325 79734
rect 170581 79731 170647 79734
rect 171358 79732 171364 79796
rect 171428 79794 171434 79796
rect 173203 79794 173269 79797
rect 175089 79794 175155 79797
rect 171428 79792 173269 79794
rect 171428 79736 173208 79792
rect 173264 79736 173269 79792
rect 171428 79734 173269 79736
rect 171428 79732 171434 79734
rect 173203 79731 173269 79734
rect 173344 79792 175155 79794
rect 173344 79736 175094 79792
rect 175150 79736 175155 79792
rect 173344 79734 175155 79736
rect 169937 79658 170003 79661
rect 169710 79656 170003 79658
rect 169710 79600 169942 79656
rect 169998 79600 170003 79656
rect 169710 79598 170003 79600
rect 167932 79596 167938 79598
rect 168281 79595 168347 79598
rect 169937 79595 170003 79598
rect 170397 79658 170463 79661
rect 170622 79658 170628 79660
rect 170397 79656 170628 79658
rect 170397 79600 170402 79656
rect 170458 79600 170628 79656
rect 170397 79598 170628 79600
rect 170397 79595 170463 79598
rect 170622 79596 170628 79598
rect 170692 79596 170698 79660
rect 171041 79658 171107 79661
rect 173344 79658 173404 79734
rect 175089 79731 175155 79734
rect 173617 79660 173683 79661
rect 171041 79656 173404 79658
rect 171041 79600 171046 79656
rect 171102 79600 173404 79656
rect 171041 79598 173404 79600
rect 171041 79595 171107 79598
rect 173566 79596 173572 79660
rect 173636 79658 173683 79660
rect 173636 79656 173728 79658
rect 173678 79600 173728 79656
rect 173636 79598 173728 79600
rect 173636 79596 173683 79598
rect 173617 79595 173683 79596
rect 6913 79522 6979 79525
rect 172973 79522 173039 79525
rect 6913 79520 173039 79522
rect 6913 79464 6918 79520
rect 6974 79464 172978 79520
rect 173034 79464 173039 79520
rect 6913 79462 173039 79464
rect 6913 79459 6979 79462
rect 172973 79459 173039 79462
rect 173198 79460 173204 79524
rect 173268 79522 173274 79524
rect 173341 79522 173407 79525
rect 173268 79520 173407 79522
rect 173268 79464 173346 79520
rect 173402 79464 173407 79520
rect 173268 79462 173407 79464
rect 173268 79460 173274 79462
rect 173341 79459 173407 79462
rect 3785 79386 3851 79389
rect 164417 79386 164483 79389
rect 173249 79386 173315 79389
rect 3785 79384 164483 79386
rect 3785 79328 3790 79384
rect 3846 79328 164422 79384
rect 164478 79328 164483 79384
rect 3785 79326 164483 79328
rect 3785 79323 3851 79326
rect 164417 79323 164483 79326
rect 164558 79384 173315 79386
rect 164558 79328 173254 79384
rect 173310 79328 173315 79384
rect 164558 79326 173315 79328
rect 3601 79250 3667 79253
rect 164558 79250 164618 79326
rect 173249 79323 173315 79326
rect 3601 79248 164618 79250
rect 3601 79192 3606 79248
rect 3662 79192 164618 79248
rect 3601 79190 164618 79192
rect 164785 79250 164851 79253
rect 173985 79250 174051 79253
rect 164785 79248 174051 79250
rect 164785 79192 164790 79248
rect 164846 79192 173990 79248
rect 174046 79192 174051 79248
rect 164785 79190 174051 79192
rect 3601 79187 3667 79190
rect 164785 79187 164851 79190
rect 173985 79187 174051 79190
rect 3417 79114 3483 79117
rect 159214 79114 159220 79116
rect 3417 79112 159220 79114
rect 3417 79056 3422 79112
rect 3478 79056 159220 79112
rect 3417 79054 159220 79056
rect 3417 79051 3483 79054
rect 159214 79052 159220 79054
rect 159284 79052 159290 79116
rect 160369 79114 160435 79117
rect 161238 79114 161244 79116
rect 160369 79112 161244 79114
rect 160369 79056 160374 79112
rect 160430 79056 161244 79112
rect 160369 79054 161244 79056
rect 160369 79051 160435 79054
rect 161238 79052 161244 79054
rect 161308 79052 161314 79116
rect 163630 79052 163636 79116
rect 163700 79114 163706 79116
rect 164049 79114 164115 79117
rect 163700 79112 164115 79114
rect 163700 79056 164054 79112
rect 164110 79056 164115 79112
rect 163700 79054 164115 79056
rect 163700 79052 163706 79054
rect 164049 79051 164115 79054
rect 164417 79114 164483 79117
rect 173433 79114 173499 79117
rect 164417 79112 173499 79114
rect 164417 79056 164422 79112
rect 164478 79056 173438 79112
rect 173494 79056 173499 79112
rect 164417 79054 173499 79056
rect 164417 79051 164483 79054
rect 173433 79051 173499 79054
rect 3233 78978 3299 78981
rect 3233 78976 171748 78978
rect 3233 78920 3238 78976
rect 3294 78920 171748 78976
rect 3233 78918 171748 78920
rect 3233 78915 3299 78918
rect 125777 78842 125843 78845
rect 125910 78842 125916 78844
rect 125777 78840 125916 78842
rect 125777 78784 125782 78840
rect 125838 78784 125916 78840
rect 125777 78782 125916 78784
rect 125777 78779 125843 78782
rect 125910 78780 125916 78782
rect 125980 78780 125986 78844
rect 128537 78842 128603 78845
rect 128670 78842 128676 78844
rect 128537 78840 128676 78842
rect 128537 78784 128542 78840
rect 128598 78784 128676 78840
rect 128537 78782 128676 78784
rect 128537 78779 128603 78782
rect 128670 78780 128676 78782
rect 128740 78780 128746 78844
rect 130009 78842 130075 78845
rect 130326 78842 130332 78844
rect 130009 78840 130332 78842
rect 130009 78784 130014 78840
rect 130070 78784 130332 78840
rect 130009 78782 130332 78784
rect 130009 78779 130075 78782
rect 130326 78780 130332 78782
rect 130396 78780 130402 78844
rect 131614 78780 131620 78844
rect 131684 78842 131690 78844
rect 131757 78842 131823 78845
rect 144361 78844 144427 78845
rect 131684 78840 131823 78842
rect 131684 78784 131762 78840
rect 131818 78784 131823 78840
rect 131684 78782 131823 78784
rect 131684 78780 131690 78782
rect 131757 78779 131823 78782
rect 144310 78780 144316 78844
rect 144380 78842 144427 78844
rect 144380 78840 144472 78842
rect 144422 78784 144472 78840
rect 144380 78782 144472 78784
rect 144380 78780 144427 78782
rect 146150 78780 146156 78844
rect 146220 78842 146226 78844
rect 146753 78842 146819 78845
rect 146220 78840 146819 78842
rect 146220 78784 146758 78840
rect 146814 78784 146819 78840
rect 146220 78782 146819 78784
rect 146220 78780 146226 78782
rect 144361 78779 144427 78780
rect 146753 78779 146819 78782
rect 146937 78842 147003 78845
rect 160093 78842 160159 78845
rect 166349 78842 166415 78845
rect 146937 78840 154590 78842
rect 146937 78784 146942 78840
rect 146998 78784 154590 78840
rect 146937 78782 154590 78784
rect 146937 78779 147003 78782
rect 125869 78708 125935 78709
rect 125869 78704 125916 78708
rect 125980 78706 125986 78708
rect 129825 78706 129891 78709
rect 130142 78706 130148 78708
rect 125869 78648 125874 78704
rect 125869 78644 125916 78648
rect 125980 78646 126026 78706
rect 129825 78704 130148 78706
rect 129825 78648 129830 78704
rect 129886 78648 130148 78704
rect 129825 78646 130148 78648
rect 125980 78644 125986 78646
rect 125869 78643 125935 78644
rect 129825 78643 129891 78646
rect 130142 78644 130148 78646
rect 130212 78644 130218 78708
rect 138974 78644 138980 78708
rect 139044 78706 139050 78708
rect 139117 78706 139183 78709
rect 139044 78704 139183 78706
rect 139044 78648 139122 78704
rect 139178 78648 139183 78704
rect 139044 78646 139183 78648
rect 139044 78644 139050 78646
rect 139117 78643 139183 78646
rect 149973 78708 150039 78709
rect 149973 78704 150020 78708
rect 150084 78706 150090 78708
rect 154530 78706 154590 78782
rect 160093 78840 166415 78842
rect 160093 78784 160098 78840
rect 160154 78784 166354 78840
rect 166410 78784 166415 78840
rect 160093 78782 166415 78784
rect 160093 78779 160159 78782
rect 166349 78779 166415 78782
rect 169385 78842 169451 78845
rect 170673 78842 170739 78845
rect 169385 78840 170739 78842
rect 169385 78784 169390 78840
rect 169446 78784 170678 78840
rect 170734 78784 170739 78840
rect 169385 78782 170739 78784
rect 169385 78779 169451 78782
rect 170673 78779 170739 78782
rect 171133 78842 171199 78845
rect 171542 78842 171548 78844
rect 171133 78840 171548 78842
rect 171133 78784 171138 78840
rect 171194 78784 171548 78840
rect 171133 78782 171548 78784
rect 171133 78779 171199 78782
rect 171542 78780 171548 78782
rect 171612 78780 171618 78844
rect 171688 78842 171748 78918
rect 171910 78916 171916 78980
rect 171980 78978 171986 78980
rect 173065 78978 173131 78981
rect 171980 78976 173131 78978
rect 171980 78920 173070 78976
rect 173126 78920 173131 78976
rect 171980 78918 173131 78920
rect 171980 78916 171986 78918
rect 173065 78915 173131 78918
rect 173157 78842 173223 78845
rect 171688 78840 173223 78842
rect 171688 78784 173162 78840
rect 173218 78784 173223 78840
rect 171688 78782 173223 78784
rect 173157 78779 173223 78782
rect 176561 78842 176627 78845
rect 397453 78842 397519 78845
rect 176561 78840 397519 78842
rect 176561 78784 176566 78840
rect 176622 78784 397458 78840
rect 397514 78784 397519 78840
rect 176561 78782 397519 78784
rect 176561 78779 176627 78782
rect 397453 78779 397519 78782
rect 163405 78706 163471 78709
rect 149973 78648 149978 78704
rect 149973 78644 150020 78648
rect 150084 78646 150130 78706
rect 154530 78704 163471 78706
rect 154530 78648 163410 78704
rect 163466 78648 163471 78704
rect 154530 78646 163471 78648
rect 150084 78644 150090 78646
rect 149973 78643 150039 78644
rect 163405 78643 163471 78646
rect 167678 78644 167684 78708
rect 167748 78706 167754 78708
rect 168097 78706 168163 78709
rect 170121 78708 170187 78709
rect 170070 78706 170076 78708
rect 167748 78704 168163 78706
rect 167748 78648 168102 78704
rect 168158 78648 168163 78704
rect 167748 78646 168163 78648
rect 170030 78646 170076 78706
rect 170140 78704 170187 78708
rect 170182 78648 170187 78704
rect 167748 78644 167754 78646
rect 168097 78643 168163 78646
rect 170070 78644 170076 78646
rect 170140 78644 170187 78648
rect 170121 78643 170187 78644
rect 170949 78708 171015 78709
rect 170949 78704 170996 78708
rect 171060 78706 171066 78708
rect 170949 78648 170954 78704
rect 170949 78644 170996 78648
rect 171060 78646 171106 78706
rect 171060 78644 171066 78646
rect 172462 78644 172468 78708
rect 172532 78706 172538 78708
rect 462313 78706 462379 78709
rect 172532 78704 462379 78706
rect 172532 78648 462318 78704
rect 462374 78648 462379 78704
rect 172532 78646 462379 78648
rect 172532 78644 172538 78646
rect 170949 78643 171015 78644
rect 462313 78643 462379 78646
rect 128813 78570 128879 78573
rect 129038 78570 129044 78572
rect 128813 78568 129044 78570
rect 128813 78512 128818 78568
rect 128874 78512 129044 78568
rect 128813 78510 129044 78512
rect 128813 78507 128879 78510
rect 129038 78508 129044 78510
rect 129108 78508 129114 78572
rect 129365 78570 129431 78573
rect 130878 78570 130884 78572
rect 129365 78568 130884 78570
rect 129365 78512 129370 78568
rect 129426 78512 130884 78568
rect 129365 78510 130884 78512
rect 129365 78507 129431 78510
rect 130878 78508 130884 78510
rect 130948 78508 130954 78572
rect 139301 78570 139367 78573
rect 141969 78570 142035 78573
rect 139301 78568 142035 78570
rect 139301 78512 139306 78568
rect 139362 78512 141974 78568
rect 142030 78512 142035 78568
rect 139301 78510 142035 78512
rect 139301 78507 139367 78510
rect 141969 78507 142035 78510
rect 145230 78508 145236 78572
rect 145300 78570 145306 78572
rect 146293 78570 146359 78573
rect 145300 78568 146359 78570
rect 145300 78512 146298 78568
rect 146354 78512 146359 78568
rect 145300 78510 146359 78512
rect 145300 78508 145306 78510
rect 146293 78507 146359 78510
rect 149462 78508 149468 78572
rect 149532 78570 149538 78572
rect 150249 78570 150315 78573
rect 149532 78568 150315 78570
rect 149532 78512 150254 78568
rect 150310 78512 150315 78568
rect 149532 78510 150315 78512
rect 149532 78508 149538 78510
rect 150249 78507 150315 78510
rect 152733 78570 152799 78573
rect 160134 78570 160140 78572
rect 152733 78568 160140 78570
rect 152733 78512 152738 78568
rect 152794 78512 160140 78568
rect 152733 78510 160140 78512
rect 152733 78507 152799 78510
rect 160134 78508 160140 78510
rect 160204 78508 160210 78572
rect 162761 78570 162827 78573
rect 162761 78568 171794 78570
rect 162761 78512 162766 78568
rect 162822 78512 171794 78568
rect 162761 78510 171794 78512
rect 162761 78507 162827 78510
rect 131430 78372 131436 78436
rect 131500 78434 131506 78436
rect 131757 78434 131823 78437
rect 131500 78432 131823 78434
rect 131500 78376 131762 78432
rect 131818 78376 131823 78432
rect 131500 78374 131823 78376
rect 131500 78372 131506 78374
rect 131757 78371 131823 78374
rect 148542 78372 148548 78436
rect 148612 78434 148618 78436
rect 149053 78434 149119 78437
rect 148612 78432 149119 78434
rect 148612 78376 149058 78432
rect 149114 78376 149119 78432
rect 148612 78374 149119 78376
rect 148612 78372 148618 78374
rect 149053 78371 149119 78374
rect 155033 78298 155099 78301
rect 164785 78298 164851 78301
rect 155033 78296 164851 78298
rect 155033 78240 155038 78296
rect 155094 78240 164790 78296
rect 164846 78240 164851 78296
rect 155033 78238 164851 78240
rect 155033 78235 155099 78238
rect 164785 78235 164851 78238
rect 165153 78298 165219 78301
rect 171317 78298 171383 78301
rect 165153 78296 171383 78298
rect 165153 78240 165158 78296
rect 165214 78240 171322 78296
rect 171378 78240 171383 78296
rect 165153 78238 171383 78240
rect 165153 78235 165219 78238
rect 171317 78235 171383 78238
rect 136909 78164 136975 78165
rect 155033 78164 155099 78165
rect 136909 78162 136956 78164
rect 136864 78160 136956 78162
rect 136864 78104 136914 78160
rect 136864 78102 136956 78104
rect 136909 78100 136956 78102
rect 137020 78100 137026 78164
rect 154982 78100 154988 78164
rect 155052 78162 155099 78164
rect 157057 78162 157123 78165
rect 171133 78162 171199 78165
rect 155052 78160 155144 78162
rect 155094 78104 155144 78160
rect 155052 78102 155144 78104
rect 157057 78160 171199 78162
rect 157057 78104 157062 78160
rect 157118 78104 171138 78160
rect 171194 78104 171199 78160
rect 157057 78102 171199 78104
rect 155052 78100 155099 78102
rect 136909 78099 136975 78100
rect 155033 78099 155099 78100
rect 157057 78099 157123 78102
rect 171133 78099 171199 78102
rect 146661 78028 146727 78029
rect 146661 78026 146708 78028
rect 146616 78024 146708 78026
rect 146616 77968 146666 78024
rect 146616 77966 146708 77968
rect 146661 77964 146708 77966
rect 146772 77964 146778 78028
rect 146937 78026 147003 78029
rect 147305 78028 147371 78029
rect 147070 78026 147076 78028
rect 146937 78024 147076 78026
rect 146937 77968 146942 78024
rect 146998 77968 147076 78024
rect 146937 77966 147076 77968
rect 146661 77963 146727 77964
rect 146937 77963 147003 77966
rect 147070 77964 147076 77966
rect 147140 77964 147146 78028
rect 147254 78026 147260 78028
rect 147214 77966 147260 78026
rect 147324 78024 147371 78028
rect 147366 77968 147371 78024
rect 147254 77964 147260 77966
rect 147324 77964 147371 77968
rect 147305 77963 147371 77964
rect 159725 78026 159791 78029
rect 171734 78026 171794 78510
rect 172053 78434 172119 78437
rect 396758 78434 396764 78436
rect 172053 78432 396764 78434
rect 172053 78376 172058 78432
rect 172114 78376 396764 78432
rect 172053 78374 396764 78376
rect 172053 78371 172119 78374
rect 396758 78372 396764 78374
rect 396828 78372 396834 78436
rect 172237 78162 172303 78165
rect 396574 78162 396580 78164
rect 172237 78160 396580 78162
rect 172237 78104 172242 78160
rect 172298 78104 396580 78160
rect 172237 78102 396580 78104
rect 172237 78099 172303 78102
rect 396574 78100 396580 78102
rect 396644 78100 396650 78164
rect 478873 78026 478939 78029
rect 159725 78024 171426 78026
rect 159725 77968 159730 78024
rect 159786 77968 171426 78024
rect 159725 77966 171426 77968
rect 171734 78024 478939 78026
rect 171734 77968 478878 78024
rect 478934 77968 478939 78024
rect 171734 77966 478939 77968
rect 159725 77963 159791 77966
rect 148358 77828 148364 77892
rect 148428 77890 148434 77892
rect 148777 77890 148843 77893
rect 148428 77888 148843 77890
rect 148428 77832 148782 77888
rect 148838 77832 148843 77888
rect 148428 77830 148843 77832
rect 148428 77828 148434 77830
rect 148777 77827 148843 77830
rect 156965 77890 157031 77893
rect 165153 77890 165219 77893
rect 156965 77888 165219 77890
rect 156965 77832 156970 77888
rect 157026 77832 165158 77888
rect 165214 77832 165219 77888
rect 156965 77830 165219 77832
rect 156965 77827 157031 77830
rect 165153 77827 165219 77830
rect 131982 77692 131988 77756
rect 132052 77754 132058 77756
rect 171366 77754 171426 77966
rect 478873 77963 478939 77966
rect 171501 77890 171567 77893
rect 483013 77890 483079 77893
rect 171501 77888 483079 77890
rect 171501 77832 171506 77888
rect 171562 77832 483018 77888
rect 483074 77832 483079 77888
rect 171501 77830 483079 77832
rect 171501 77827 171567 77830
rect 483013 77827 483079 77830
rect 171961 77754 172027 77757
rect 132052 77694 138030 77754
rect 171366 77752 172027 77754
rect 171366 77696 171966 77752
rect 172022 77696 172027 77752
rect 171366 77694 172027 77696
rect 132052 77692 132058 77694
rect 125869 77618 125935 77621
rect 127382 77618 127388 77620
rect 125869 77616 127388 77618
rect 125869 77560 125874 77616
rect 125930 77560 127388 77616
rect 125869 77558 127388 77560
rect 125869 77555 125935 77558
rect 127382 77556 127388 77558
rect 127452 77556 127458 77620
rect 137970 77618 138030 77694
rect 171961 77691 172027 77694
rect 147673 77618 147739 77621
rect 137970 77616 147739 77618
rect 137970 77560 147678 77616
rect 147734 77560 147739 77616
rect 137970 77558 147739 77560
rect 147673 77555 147739 77558
rect 155953 77618 156019 77621
rect 162669 77618 162735 77621
rect 155953 77616 162735 77618
rect 155953 77560 155958 77616
rect 156014 77560 162674 77616
rect 162730 77560 162735 77616
rect 155953 77558 162735 77560
rect 155953 77555 156019 77558
rect 162669 77555 162735 77558
rect 171317 77618 171383 77621
rect 172145 77618 172211 77621
rect 171317 77616 172211 77618
rect 171317 77560 171322 77616
rect 171378 77560 172150 77616
rect 172206 77560 172211 77616
rect 171317 77558 172211 77560
rect 171317 77555 171383 77558
rect 172145 77555 172211 77558
rect 127157 77482 127223 77485
rect 127382 77482 127388 77484
rect 127157 77480 127388 77482
rect 127157 77424 127162 77480
rect 127218 77424 127388 77480
rect 127157 77422 127388 77424
rect 127157 77419 127223 77422
rect 127382 77420 127388 77422
rect 127452 77420 127458 77484
rect 171133 77482 171199 77485
rect 172329 77482 172395 77485
rect 171133 77480 172395 77482
rect 171133 77424 171138 77480
rect 171194 77424 172334 77480
rect 172390 77424 172395 77480
rect 171133 77422 172395 77424
rect 171133 77419 171199 77422
rect 172329 77419 172395 77422
rect 127249 77348 127315 77349
rect 127198 77284 127204 77348
rect 127268 77346 127315 77348
rect 127268 77344 127360 77346
rect 127310 77288 127360 77344
rect 127268 77286 127360 77288
rect 127268 77284 127315 77286
rect 147070 77284 147076 77348
rect 147140 77346 147146 77348
rect 147397 77346 147463 77349
rect 147140 77344 147463 77346
rect 147140 77288 147402 77344
rect 147458 77288 147463 77344
rect 147140 77286 147463 77288
rect 147140 77284 147146 77286
rect 127249 77283 127315 77284
rect 147397 77283 147463 77286
rect 160277 77346 160343 77349
rect 161238 77346 161244 77348
rect 160277 77344 161244 77346
rect 160277 77288 160282 77344
rect 160338 77288 161244 77344
rect 160277 77286 161244 77288
rect 160277 77283 160343 77286
rect 161238 77284 161244 77286
rect 161308 77284 161314 77348
rect 169150 77284 169156 77348
rect 169220 77346 169226 77348
rect 171174 77346 171180 77348
rect 169220 77286 171180 77346
rect 169220 77284 169226 77286
rect 171174 77284 171180 77286
rect 171244 77284 171250 77348
rect 173249 77210 173315 77213
rect 150390 77208 173315 77210
rect 150390 77152 173254 77208
rect 173310 77152 173315 77208
rect 150390 77150 173315 77152
rect 131297 77076 131363 77077
rect 131246 77074 131252 77076
rect 131206 77014 131252 77074
rect 131316 77072 131363 77076
rect 131358 77016 131363 77072
rect 131246 77012 131252 77014
rect 131316 77012 131363 77016
rect 133822 77012 133828 77076
rect 133892 77074 133898 77076
rect 134241 77074 134307 77077
rect 133892 77072 134307 77074
rect 133892 77016 134246 77072
rect 134302 77016 134307 77072
rect 133892 77014 134307 77016
rect 133892 77012 133898 77014
rect 131297 77011 131363 77012
rect 134241 77011 134307 77014
rect 142153 77074 142219 77077
rect 150390 77074 150450 77150
rect 173249 77147 173315 77150
rect 142153 77072 150450 77074
rect 142153 77016 142158 77072
rect 142214 77016 150450 77072
rect 142153 77014 150450 77016
rect 142153 77011 142219 77014
rect 152590 77012 152596 77076
rect 152660 77074 152666 77076
rect 153377 77074 153443 77077
rect 152660 77072 153443 77074
rect 152660 77016 153382 77072
rect 153438 77016 153443 77072
rect 152660 77014 153443 77016
rect 152660 77012 152666 77014
rect 153377 77011 153443 77014
rect 111793 76938 111859 76941
rect 133270 76938 133276 76940
rect 111793 76936 133276 76938
rect 111793 76880 111798 76936
rect 111854 76880 133276 76936
rect 111793 76878 133276 76880
rect 111793 76875 111859 76878
rect 133270 76876 133276 76878
rect 133340 76876 133346 76940
rect 144821 76938 144887 76941
rect 247033 76938 247099 76941
rect 144821 76936 247099 76938
rect 144821 76880 144826 76936
rect 144882 76880 247038 76936
rect 247094 76880 247099 76936
rect 144821 76878 247099 76880
rect 144821 76875 144887 76878
rect 247033 76875 247099 76878
rect 93853 76802 93919 76805
rect 131798 76802 131804 76804
rect 93853 76800 131804 76802
rect 93853 76744 93858 76800
rect 93914 76744 131804 76800
rect 93853 76742 131804 76744
rect 93853 76739 93919 76742
rect 131798 76740 131804 76742
rect 131868 76740 131874 76804
rect 137686 76740 137692 76804
rect 137756 76802 137762 76804
rect 137829 76802 137895 76805
rect 137756 76800 137895 76802
rect 137756 76744 137834 76800
rect 137890 76744 137895 76800
rect 137756 76742 137895 76744
rect 137756 76740 137762 76742
rect 137829 76739 137895 76742
rect 147489 76802 147555 76805
rect 282913 76802 282979 76805
rect 147489 76800 282979 76802
rect 147489 76744 147494 76800
rect 147550 76744 282918 76800
rect 282974 76744 282979 76800
rect 147489 76742 282979 76744
rect 147489 76739 147555 76742
rect 282913 76739 282979 76742
rect 20713 76666 20779 76669
rect 127065 76666 127131 76669
rect 20713 76664 127131 76666
rect 20713 76608 20718 76664
rect 20774 76608 127070 76664
rect 127126 76608 127131 76664
rect 20713 76606 127131 76608
rect 20713 76603 20779 76606
rect 127065 76603 127131 76606
rect 132769 76666 132835 76669
rect 133454 76666 133460 76668
rect 132769 76664 133460 76666
rect 132769 76608 132774 76664
rect 132830 76608 133460 76664
rect 132769 76606 133460 76608
rect 132769 76603 132835 76606
rect 133454 76604 133460 76606
rect 133524 76604 133530 76668
rect 133965 76666 134031 76669
rect 134609 76668 134675 76669
rect 134190 76666 134196 76668
rect 133965 76664 134196 76666
rect 133965 76608 133970 76664
rect 134026 76608 134196 76664
rect 133965 76606 134196 76608
rect 133965 76603 134031 76606
rect 134190 76604 134196 76606
rect 134260 76604 134266 76668
rect 134558 76604 134564 76668
rect 134628 76666 134675 76668
rect 135529 76666 135595 76669
rect 137921 76668 137987 76669
rect 136398 76666 136404 76668
rect 134628 76664 134720 76666
rect 134670 76608 134720 76664
rect 134628 76606 134720 76608
rect 135529 76664 136404 76666
rect 135529 76608 135534 76664
rect 135590 76608 136404 76664
rect 135529 76606 136404 76608
rect 134628 76604 134675 76606
rect 134609 76603 134675 76604
rect 135529 76603 135595 76606
rect 136398 76604 136404 76606
rect 136468 76604 136474 76668
rect 137870 76666 137876 76668
rect 137830 76606 137876 76666
rect 137940 76664 137987 76668
rect 137982 76608 137987 76664
rect 137870 76604 137876 76606
rect 137940 76604 137987 76608
rect 138054 76604 138060 76668
rect 138124 76666 138130 76668
rect 140405 76666 140471 76669
rect 138124 76664 140471 76666
rect 138124 76608 140410 76664
rect 140466 76608 140471 76664
rect 138124 76606 140471 76608
rect 138124 76604 138130 76606
rect 137921 76603 137987 76604
rect 140405 76603 140471 76606
rect 151629 76668 151695 76669
rect 153009 76668 153075 76669
rect 151629 76664 151676 76668
rect 151740 76666 151746 76668
rect 152958 76666 152964 76668
rect 151629 76608 151634 76664
rect 151629 76604 151676 76608
rect 151740 76606 151786 76666
rect 152918 76606 152964 76666
rect 153028 76664 153075 76668
rect 153070 76608 153075 76664
rect 151740 76604 151746 76606
rect 152958 76604 152964 76606
rect 153028 76604 153075 76608
rect 151629 76603 151695 76604
rect 153009 76603 153075 76604
rect 153377 76666 153443 76669
rect 154389 76668 154455 76669
rect 155585 76668 155651 76669
rect 154062 76666 154068 76668
rect 153377 76664 154068 76666
rect 153377 76608 153382 76664
rect 153438 76608 154068 76664
rect 153377 76606 154068 76608
rect 153377 76603 153443 76606
rect 154062 76604 154068 76606
rect 154132 76604 154138 76668
rect 154389 76664 154436 76668
rect 154500 76666 154506 76668
rect 155534 76666 155540 76668
rect 154389 76608 154394 76664
rect 154389 76604 154436 76608
rect 154500 76606 154546 76666
rect 155494 76606 155540 76666
rect 155604 76664 155651 76668
rect 155646 76608 155651 76664
rect 154500 76604 154506 76606
rect 155534 76604 155540 76606
rect 155604 76604 155651 76608
rect 156086 76604 156092 76668
rect 156156 76666 156162 76668
rect 156413 76666 156479 76669
rect 156156 76664 156479 76666
rect 156156 76608 156418 76664
rect 156474 76608 156479 76664
rect 156156 76606 156479 76608
rect 156156 76604 156162 76606
rect 154389 76603 154455 76604
rect 155585 76603 155651 76604
rect 156413 76603 156479 76606
rect 156638 76604 156644 76668
rect 156708 76666 156714 76668
rect 157241 76666 157307 76669
rect 156708 76664 157307 76666
rect 156708 76608 157246 76664
rect 157302 76608 157307 76664
rect 156708 76606 157307 76608
rect 156708 76604 156714 76606
rect 157241 76603 157307 76606
rect 157517 76666 157583 76669
rect 158529 76668 158595 76669
rect 157742 76666 157748 76668
rect 157517 76664 157748 76666
rect 157517 76608 157522 76664
rect 157578 76608 157748 76664
rect 157517 76606 157748 76608
rect 157517 76603 157583 76606
rect 157742 76604 157748 76606
rect 157812 76604 157818 76668
rect 158478 76666 158484 76668
rect 158438 76606 158484 76666
rect 158548 76664 158595 76668
rect 158590 76608 158595 76664
rect 158478 76604 158484 76606
rect 158548 76604 158595 76608
rect 160870 76604 160876 76668
rect 160940 76666 160946 76668
rect 161381 76666 161447 76669
rect 160940 76664 161447 76666
rect 160940 76608 161386 76664
rect 161442 76608 161447 76664
rect 160940 76606 161447 76608
rect 160940 76604 160946 76606
rect 158529 76603 158595 76604
rect 161381 76603 161447 76606
rect 164417 76666 164483 76669
rect 165429 76668 165495 76669
rect 166809 76668 166875 76669
rect 164918 76666 164924 76668
rect 164417 76664 164924 76666
rect 164417 76608 164422 76664
rect 164478 76608 164924 76664
rect 164417 76606 164924 76608
rect 164417 76603 164483 76606
rect 164918 76604 164924 76606
rect 164988 76604 164994 76668
rect 165429 76664 165476 76668
rect 165540 76666 165546 76668
rect 166758 76666 166764 76668
rect 165429 76608 165434 76664
rect 165429 76604 165476 76608
rect 165540 76606 165586 76666
rect 166718 76606 166764 76666
rect 166828 76664 166875 76668
rect 166870 76608 166875 76664
rect 165540 76604 165546 76606
rect 166758 76604 166764 76606
rect 166828 76604 166875 76608
rect 168046 76604 168052 76668
rect 168116 76666 168122 76668
rect 168189 76666 168255 76669
rect 168116 76664 168255 76666
rect 168116 76608 168194 76664
rect 168250 76608 168255 76664
rect 168116 76606 168255 76608
rect 168116 76604 168122 76606
rect 165429 76603 165495 76604
rect 166809 76603 166875 76604
rect 168189 76603 168255 76606
rect 169385 76666 169451 76669
rect 549253 76666 549319 76669
rect 169385 76664 549319 76666
rect 169385 76608 169390 76664
rect 169446 76608 549258 76664
rect 549314 76608 549319 76664
rect 169385 76606 549319 76608
rect 169385 76603 169451 76606
rect 549253 76603 549319 76606
rect 1393 76530 1459 76533
rect 125593 76530 125659 76533
rect 1393 76528 125659 76530
rect 1393 76472 1398 76528
rect 1454 76472 125598 76528
rect 125654 76472 125659 76528
rect 1393 76470 125659 76472
rect 1393 76467 1459 76470
rect 125593 76467 125659 76470
rect 136398 76468 136404 76532
rect 136468 76530 136474 76532
rect 138013 76530 138079 76533
rect 136468 76528 138079 76530
rect 136468 76472 138018 76528
rect 138074 76472 138079 76528
rect 136468 76470 138079 76472
rect 136468 76468 136474 76470
rect 138013 76467 138079 76470
rect 151302 76468 151308 76532
rect 151372 76530 151378 76532
rect 151721 76530 151787 76533
rect 152825 76532 152891 76533
rect 152774 76530 152780 76532
rect 151372 76528 151787 76530
rect 151372 76472 151726 76528
rect 151782 76472 151787 76528
rect 151372 76470 151787 76472
rect 152734 76470 152780 76530
rect 152844 76528 152891 76532
rect 152886 76472 152891 76528
rect 151372 76468 151378 76470
rect 151721 76467 151787 76470
rect 152774 76468 152780 76470
rect 152844 76468 152891 76472
rect 154062 76468 154068 76532
rect 154132 76530 154138 76532
rect 154481 76530 154547 76533
rect 154132 76528 154547 76530
rect 154132 76472 154486 76528
rect 154542 76472 154547 76528
rect 154132 76470 154547 76472
rect 154132 76468 154138 76470
rect 152825 76467 152891 76468
rect 154481 76467 154547 76470
rect 157926 76468 157932 76532
rect 157996 76530 158002 76532
rect 158437 76530 158503 76533
rect 157996 76528 158503 76530
rect 157996 76472 158442 76528
rect 158498 76472 158503 76528
rect 157996 76470 158503 76472
rect 157996 76468 158002 76470
rect 158437 76467 158503 76470
rect 160686 76468 160692 76532
rect 160756 76530 160762 76532
rect 161105 76530 161171 76533
rect 160756 76528 161171 76530
rect 160756 76472 161110 76528
rect 161166 76472 161171 76528
rect 160756 76470 161171 76472
rect 160756 76468 160762 76470
rect 161105 76467 161171 76470
rect 164918 76468 164924 76532
rect 164988 76530 164994 76532
rect 165521 76530 165587 76533
rect 164988 76528 165587 76530
rect 164988 76472 165526 76528
rect 165582 76472 165587 76528
rect 164988 76470 165587 76472
rect 164988 76468 164994 76470
rect 165521 76467 165587 76470
rect 168833 76530 168899 76533
rect 169334 76530 169340 76532
rect 168833 76528 169340 76530
rect 168833 76472 168838 76528
rect 168894 76472 169340 76528
rect 168833 76470 169340 76472
rect 168833 76467 168899 76470
rect 169334 76468 169340 76470
rect 169404 76468 169410 76532
rect 169569 76530 169635 76533
rect 565813 76530 565879 76533
rect 169569 76528 565879 76530
rect 169569 76472 169574 76528
rect 169630 76472 565818 76528
rect 565874 76472 565879 76528
rect 169569 76470 565879 76472
rect 169569 76467 169635 76470
rect 565813 76467 565879 76470
rect 140129 76394 140195 76397
rect 140446 76394 140452 76396
rect 140129 76392 140452 76394
rect 140129 76336 140134 76392
rect 140190 76336 140452 76392
rect 140129 76334 140452 76336
rect 140129 76331 140195 76334
rect 140446 76332 140452 76334
rect 140516 76332 140522 76396
rect 151854 76332 151860 76396
rect 151924 76394 151930 76396
rect 154205 76394 154271 76397
rect 151924 76392 154271 76394
rect 151924 76336 154210 76392
rect 154266 76336 154271 76392
rect 151924 76334 154271 76336
rect 151924 76332 151930 76334
rect 154205 76331 154271 76334
rect 160369 76394 160435 76397
rect 167545 76396 167611 76397
rect 161054 76394 161060 76396
rect 160369 76392 161060 76394
rect 160369 76336 160374 76392
rect 160430 76336 161060 76392
rect 160369 76334 161060 76336
rect 160369 76331 160435 76334
rect 161054 76332 161060 76334
rect 161124 76332 161130 76396
rect 167494 76332 167500 76396
rect 167564 76394 167611 76396
rect 167564 76392 167656 76394
rect 167606 76336 167656 76392
rect 167564 76334 167656 76336
rect 167564 76332 167611 76334
rect 167545 76331 167611 76332
rect 158846 76196 158852 76260
rect 158916 76258 158922 76260
rect 160001 76258 160067 76261
rect 158916 76256 160067 76258
rect 158916 76200 160006 76256
rect 160062 76200 160067 76256
rect 158916 76198 160067 76200
rect 158916 76196 158922 76198
rect 160001 76195 160067 76198
rect 170305 76258 170371 76261
rect 170806 76258 170812 76260
rect 170305 76256 170812 76258
rect 170305 76200 170310 76256
rect 170366 76200 170812 76256
rect 170305 76198 170812 76200
rect 170305 76195 170371 76198
rect 170806 76196 170812 76198
rect 170876 76196 170882 76260
rect 144126 76060 144132 76124
rect 144196 76122 144202 76124
rect 144637 76122 144703 76125
rect 144196 76120 144703 76122
rect 144196 76064 144642 76120
rect 144698 76064 144703 76120
rect 144196 76062 144703 76064
rect 144196 76060 144202 76062
rect 144637 76059 144703 76062
rect 169334 76060 169340 76124
rect 169404 76122 169410 76124
rect 169753 76122 169819 76125
rect 169404 76120 169819 76122
rect 169404 76064 169758 76120
rect 169814 76064 169819 76120
rect 169404 76062 169819 76064
rect 169404 76060 169410 76062
rect 169753 76059 169819 76062
rect 170990 76060 170996 76124
rect 171060 76122 171066 76124
rect 177297 76122 177363 76125
rect 171060 76120 177363 76122
rect 171060 76064 177302 76120
rect 177358 76064 177363 76120
rect 171060 76062 177363 76064
rect 171060 76060 171066 76062
rect 177297 76059 177363 76062
rect 140998 75924 141004 75988
rect 141068 75986 141074 75988
rect 142061 75986 142127 75989
rect 143257 75988 143323 75989
rect 143206 75986 143212 75988
rect 141068 75984 142127 75986
rect 141068 75928 142066 75984
rect 142122 75928 142127 75984
rect 141068 75926 142127 75928
rect 143166 75926 143212 75986
rect 143276 75984 143323 75988
rect 143318 75928 143323 75984
rect 141068 75924 141074 75926
rect 142061 75923 142127 75926
rect 143206 75924 143212 75926
rect 143276 75924 143323 75928
rect 145414 75924 145420 75988
rect 145484 75986 145490 75988
rect 146109 75986 146175 75989
rect 147857 75988 147923 75989
rect 145484 75984 146175 75986
rect 145484 75928 146114 75984
rect 146170 75928 146175 75984
rect 145484 75926 146175 75928
rect 145484 75924 145490 75926
rect 143257 75923 143323 75924
rect 146109 75923 146175 75926
rect 147806 75924 147812 75988
rect 147876 75986 147923 75988
rect 147876 75984 147968 75986
rect 147918 75928 147968 75984
rect 147876 75926 147968 75928
rect 147876 75924 147923 75926
rect 148726 75924 148732 75988
rect 148796 75986 148802 75988
rect 148961 75986 149027 75989
rect 148796 75984 149027 75986
rect 148796 75928 148966 75984
rect 149022 75928 149027 75984
rect 148796 75926 149027 75928
rect 148796 75924 148802 75926
rect 147857 75923 147923 75924
rect 148961 75923 149027 75926
rect 169845 75986 169911 75989
rect 171726 75986 171732 75988
rect 169845 75984 171732 75986
rect 169845 75928 169850 75984
rect 169906 75928 171732 75984
rect 169845 75926 171732 75928
rect 169845 75923 169911 75926
rect 171726 75924 171732 75926
rect 171796 75924 171802 75988
rect 132677 75850 132743 75853
rect 133270 75850 133276 75852
rect 132677 75848 133276 75850
rect 132677 75792 132682 75848
rect 132738 75792 133276 75848
rect 132677 75790 133276 75792
rect 132677 75787 132743 75790
rect 133270 75788 133276 75790
rect 133340 75788 133346 75852
rect 143022 75788 143028 75852
rect 143092 75850 143098 75852
rect 143349 75850 143415 75853
rect 143092 75848 143415 75850
rect 143092 75792 143354 75848
rect 143410 75792 143415 75848
rect 143092 75790 143415 75792
rect 143092 75788 143098 75790
rect 143349 75787 143415 75790
rect 169753 75850 169819 75853
rect 170070 75850 170076 75852
rect 169753 75848 170076 75850
rect 169753 75792 169758 75848
rect 169814 75792 170076 75848
rect 169753 75790 170076 75792
rect 169753 75787 169819 75790
rect 170070 75788 170076 75790
rect 170140 75788 170146 75852
rect 170857 75850 170923 75853
rect 171910 75850 171916 75852
rect 170857 75848 171916 75850
rect 170857 75792 170862 75848
rect 170918 75792 171916 75848
rect 170857 75790 171916 75792
rect 170857 75787 170923 75790
rect 171910 75788 171916 75790
rect 171980 75788 171986 75852
rect 139158 75652 139164 75716
rect 139228 75714 139234 75716
rect 173893 75714 173959 75717
rect 139228 75712 173959 75714
rect 139228 75656 173898 75712
rect 173954 75656 173959 75712
rect 139228 75654 173959 75656
rect 139228 75652 139234 75654
rect 173893 75651 173959 75654
rect 57973 75578 58039 75581
rect 130326 75578 130332 75580
rect 57973 75576 130332 75578
rect 57973 75520 57978 75576
rect 58034 75520 130332 75576
rect 57973 75518 130332 75520
rect 57973 75515 58039 75518
rect 130326 75516 130332 75518
rect 130396 75516 130402 75580
rect 141969 75578 142035 75581
rect 176653 75578 176719 75581
rect 141969 75576 176719 75578
rect 141969 75520 141974 75576
rect 142030 75520 176658 75576
rect 176714 75520 176719 75576
rect 141969 75518 176719 75520
rect 141969 75515 142035 75518
rect 176653 75515 176719 75518
rect 53833 75442 53899 75445
rect 129774 75442 129780 75444
rect 53833 75440 129780 75442
rect 53833 75384 53838 75440
rect 53894 75384 129780 75440
rect 53833 75382 129780 75384
rect 53833 75379 53899 75382
rect 129774 75380 129780 75382
rect 129844 75380 129850 75444
rect 157977 75442 158043 75445
rect 402973 75442 403039 75445
rect 157977 75440 403039 75442
rect 157977 75384 157982 75440
rect 158038 75384 402978 75440
rect 403034 75384 403039 75440
rect 157977 75382 403039 75384
rect 157977 75379 158043 75382
rect 402973 75379 403039 75382
rect 35893 75306 35959 75309
rect 128353 75306 128419 75309
rect 35893 75304 128419 75306
rect 35893 75248 35898 75304
rect 35954 75248 128358 75304
rect 128414 75248 128419 75304
rect 35893 75246 128419 75248
rect 35893 75243 35959 75246
rect 128353 75243 128419 75246
rect 164550 75244 164556 75308
rect 164620 75306 164626 75308
rect 496813 75306 496879 75309
rect 164620 75304 496879 75306
rect 164620 75248 496818 75304
rect 496874 75248 496879 75304
rect 164620 75246 496879 75248
rect 164620 75244 164626 75246
rect 496813 75243 496879 75246
rect 2773 75170 2839 75173
rect 125726 75170 125732 75172
rect 2773 75168 125732 75170
rect 2773 75112 2778 75168
rect 2834 75112 125732 75168
rect 2773 75110 125732 75112
rect 2773 75107 2839 75110
rect 125726 75108 125732 75110
rect 125796 75108 125802 75172
rect 166901 75170 166967 75173
rect 528553 75170 528619 75173
rect 166901 75168 528619 75170
rect 166901 75112 166906 75168
rect 166962 75112 528558 75168
rect 528614 75112 528619 75168
rect 166901 75110 528619 75112
rect 166901 75107 166967 75110
rect 528553 75107 528619 75110
rect 130377 74490 130443 74493
rect 135253 74490 135319 74493
rect 130377 74488 135319 74490
rect 130377 74432 130382 74488
rect 130438 74432 135258 74488
rect 135314 74432 135319 74488
rect 130377 74430 135319 74432
rect 130377 74427 130443 74430
rect 135253 74427 135319 74430
rect 140589 74082 140655 74085
rect 194593 74082 194659 74085
rect 140589 74080 194659 74082
rect 140589 74024 140594 74080
rect 140650 74024 194598 74080
rect 194654 74024 194659 74080
rect 140589 74022 194659 74024
rect 140589 74019 140655 74022
rect 194593 74019 194659 74022
rect 143533 73946 143599 73949
rect 230473 73946 230539 73949
rect 143533 73944 230539 73946
rect 143533 73888 143538 73944
rect 143594 73888 230478 73944
rect 230534 73888 230539 73944
rect 143533 73886 230539 73888
rect 143533 73883 143599 73886
rect 230473 73883 230539 73886
rect 40033 73810 40099 73813
rect 128854 73810 128860 73812
rect 40033 73808 128860 73810
rect 40033 73752 40038 73808
rect 40094 73752 128860 73808
rect 40033 73750 128860 73752
rect 40033 73747 40099 73750
rect 128854 73748 128860 73750
rect 128924 73748 128930 73812
rect 146201 73810 146267 73813
rect 244273 73810 244339 73813
rect 146201 73808 244339 73810
rect 146201 73752 146206 73808
rect 146262 73752 244278 73808
rect 244334 73752 244339 73808
rect 146201 73750 244339 73752
rect 146201 73747 146267 73750
rect 244273 73747 244339 73750
rect 131062 73204 131068 73268
rect 131132 73266 131138 73268
rect 131205 73266 131271 73269
rect 131132 73264 131271 73266
rect 131132 73208 131210 73264
rect 131266 73208 131271 73264
rect 131132 73206 131271 73208
rect 131132 73204 131138 73206
rect 131205 73203 131271 73206
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect 162853 72722 162919 72725
rect 178677 72722 178743 72725
rect 162853 72720 178743 72722
rect 162853 72664 162858 72720
rect 162914 72664 178682 72720
rect 178738 72664 178743 72720
rect 162853 72662 178743 72664
rect 162853 72659 162919 72662
rect 178677 72659 178743 72662
rect 147581 72586 147647 72589
rect 284293 72586 284359 72589
rect 147581 72584 284359 72586
rect 147581 72528 147586 72584
rect 147642 72528 284298 72584
rect 284354 72528 284359 72584
rect 147581 72526 284359 72528
rect 147581 72523 147647 72526
rect 284293 72523 284359 72526
rect 148358 72388 148364 72452
rect 148428 72450 148434 72452
rect 298093 72450 298159 72453
rect 148428 72448 298159 72450
rect 148428 72392 298098 72448
rect 298154 72392 298159 72448
rect 148428 72390 298159 72392
rect 148428 72388 148434 72390
rect 298093 72387 298159 72390
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 152958 71164 152964 71228
rect 153028 71226 153034 71228
rect 353293 71226 353359 71229
rect 153028 71224 353359 71226
rect 153028 71168 353298 71224
rect 353354 71168 353359 71224
rect 153028 71166 353359 71168
rect 153028 71164 153034 71166
rect 353293 71163 353359 71166
rect 163446 71028 163452 71092
rect 163516 71090 163522 71092
rect 494053 71090 494119 71093
rect 163516 71088 494119 71090
rect 163516 71032 494058 71088
rect 494114 71032 494119 71088
rect 163516 71030 494119 71032
rect 163516 71028 163522 71030
rect 494053 71027 494119 71030
rect 138974 69532 138980 69596
rect 139044 69594 139050 69596
rect 175273 69594 175339 69597
rect 139044 69592 175339 69594
rect 139044 69536 175278 69592
rect 175334 69536 175339 69592
rect 139044 69534 175339 69536
rect 139044 69532 139050 69534
rect 175273 69531 175339 69534
rect 165470 68172 165476 68236
rect 165540 68234 165546 68236
rect 511993 68234 512059 68237
rect 165540 68232 512059 68234
rect 165540 68176 511998 68232
rect 512054 68176 512059 68232
rect 165540 68174 512059 68176
rect 165540 68172 165546 68174
rect 511993 68171 512059 68174
rect 140262 65452 140268 65516
rect 140332 65514 140338 65516
rect 193213 65514 193279 65517
rect 140332 65512 193279 65514
rect 140332 65456 193218 65512
rect 193274 65456 193279 65512
rect 140332 65454 193279 65456
rect 140332 65452 140338 65454
rect 193213 65451 193279 65454
rect 166390 62868 166396 62932
rect 166460 62930 166466 62932
rect 529933 62930 529999 62933
rect 166460 62928 529999 62930
rect 166460 62872 529938 62928
rect 529994 62872 529999 62928
rect 166460 62870 529999 62872
rect 166460 62868 166466 62870
rect 529933 62867 529999 62870
rect 171174 62732 171180 62796
rect 171244 62794 171250 62796
rect 550633 62794 550699 62797
rect 171244 62792 550699 62794
rect 171244 62736 550638 62792
rect 550694 62736 550699 62792
rect 171244 62734 550699 62736
rect 171244 62732 171250 62734
rect 550633 62731 550699 62734
rect 160686 61372 160692 61436
rect 160756 61434 160762 61436
rect 459553 61434 459619 61437
rect 160756 61432 459619 61434
rect 160756 61376 459558 61432
rect 459614 61376 459619 61432
rect 160756 61374 459619 61376
rect 160756 61372 160762 61374
rect 459553 61371 459619 61374
rect 138790 60012 138796 60076
rect 138860 60074 138866 60076
rect 172513 60074 172579 60077
rect 138860 60072 172579 60074
rect 138860 60016 172518 60072
rect 172574 60016 172579 60072
rect 138860 60014 172579 60016
rect 138860 60012 138866 60014
rect 172513 60011 172579 60014
rect 143022 59876 143028 59940
rect 143092 59938 143098 59940
rect 227713 59938 227779 59941
rect 143092 59936 227779 59938
rect 143092 59880 227718 59936
rect 227774 59880 227779 59936
rect 143092 59878 227779 59880
rect 143092 59876 143098 59878
rect 227713 59875 227779 59878
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 4061 58578 4127 58581
rect -960 58576 4127 58578
rect -960 58520 4066 58576
rect 4122 58520 4127 58576
rect -960 58518 4127 58520
rect -960 58428 480 58518
rect 4061 58515 4127 58518
rect 149462 53076 149468 53140
rect 149532 53138 149538 53140
rect 316033 53138 316099 53141
rect 149532 53136 316099 53138
rect 149532 53080 316038 53136
rect 316094 53080 316099 53136
rect 149532 53078 316099 53080
rect 149532 53076 149538 53078
rect 316033 53075 316099 53078
rect 152590 47500 152596 47564
rect 152660 47562 152666 47564
rect 351913 47562 351979 47565
rect 152660 47560 351979 47562
rect 152660 47504 351918 47560
rect 351974 47504 351979 47560
rect 152660 47502 351979 47504
rect 152660 47500 152666 47502
rect 351913 47499 351979 47502
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 127065 44978 127131 44981
rect 135294 44978 135300 44980
rect 127065 44976 135300 44978
rect 127065 44920 127070 44976
rect 127126 44920 135300 44976
rect 127065 44918 135300 44920
rect 127065 44915 127131 44918
rect 135294 44916 135300 44918
rect 135364 44916 135370 44980
rect 91093 44842 91159 44845
rect 133270 44842 133276 44844
rect 91093 44840 133276 44842
rect 91093 44784 91098 44840
rect 91154 44784 133276 44840
rect 91093 44782 133276 44784
rect 91093 44779 91159 44782
rect 133270 44780 133276 44782
rect 133340 44780 133346 44844
rect 147254 44780 147260 44844
rect 147324 44842 147330 44844
rect 280153 44842 280219 44845
rect 147324 44840 280219 44842
rect 147324 44784 280158 44840
rect 280214 44784 280219 44840
rect 147324 44782 280219 44784
rect 147324 44780 147330 44782
rect 280153 44779 280219 44782
rect 22093 43482 22159 43485
rect 127198 43482 127204 43484
rect 22093 43480 127204 43482
rect 22093 43424 22098 43480
rect 22154 43424 127204 43480
rect 22093 43422 127204 43424
rect 22093 43419 22159 43422
rect 127198 43420 127204 43422
rect 127268 43420 127274 43484
rect 153878 40564 153884 40628
rect 153948 40626 153954 40628
rect 367093 40626 367159 40629
rect 153948 40624 367159 40626
rect 153948 40568 367098 40624
rect 367154 40568 367159 40624
rect 153948 40566 367159 40568
rect 153948 40564 153954 40566
rect 367093 40563 367159 40566
rect 154062 35124 154068 35188
rect 154132 35186 154138 35188
rect 372613 35186 372679 35189
rect 154132 35184 372679 35186
rect 154132 35128 372618 35184
rect 372674 35128 372679 35184
rect 154132 35126 372679 35128
rect 154132 35124 154138 35126
rect 372613 35123 372679 35126
rect 143206 34036 143212 34100
rect 143276 34098 143282 34100
rect 226425 34098 226491 34101
rect 143276 34096 226491 34098
rect 143276 34040 226430 34096
rect 226486 34040 226491 34096
rect 143276 34038 226491 34040
rect 143276 34036 143282 34038
rect 226425 34035 226491 34038
rect 145230 33900 145236 33964
rect 145300 33962 145306 33964
rect 266353 33962 266419 33965
rect 145300 33960 266419 33962
rect 145300 33904 266358 33960
rect 266414 33904 266419 33960
rect 145300 33902 266419 33904
rect 145300 33900 145306 33902
rect 266353 33899 266419 33902
rect 170622 33764 170628 33828
rect 170692 33826 170698 33828
rect 578233 33826 578299 33829
rect 170692 33824 578299 33826
rect 170692 33768 578238 33824
rect 578294 33768 578299 33824
rect 170692 33766 578299 33768
rect 170692 33764 170698 33766
rect 578233 33763 578299 33766
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 166574 32540 166580 32604
rect 166644 32602 166650 32604
rect 531313 32602 531379 32605
rect 166644 32600 531379 32602
rect 166644 32544 531318 32600
rect 531374 32544 531379 32600
rect 166644 32542 531379 32544
rect 166644 32540 166650 32542
rect 531313 32539 531379 32542
rect 3417 32466 3483 32469
rect -960 32464 3483 32466
rect -960 32408 3422 32464
rect 3478 32408 3483 32464
rect -960 32406 3483 32408
rect -960 32316 480 32406
rect 3417 32403 3483 32406
rect 169334 32404 169340 32468
rect 169404 32466 169410 32468
rect 567193 32466 567259 32469
rect 169404 32464 567259 32466
rect 169404 32408 567198 32464
rect 567254 32408 567259 32464
rect 169404 32406 567259 32408
rect 169404 32404 169410 32406
rect 567193 32403 567259 32406
rect 167678 30908 167684 30972
rect 167748 30970 167754 30972
rect 546493 30970 546559 30973
rect 167748 30968 546559 30970
rect 167748 30912 546498 30968
rect 546554 30912 546559 30968
rect 167748 30910 546559 30912
rect 167748 30908 167754 30910
rect 546493 30907 546559 30910
rect 149646 29548 149652 29612
rect 149716 29610 149722 29612
rect 317413 29610 317479 29613
rect 149716 29608 317479 29610
rect 149716 29552 317418 29608
rect 317474 29552 317479 29608
rect 149716 29550 317479 29552
rect 149716 29548 149722 29550
rect 317413 29547 317479 29550
rect 140446 28460 140452 28524
rect 140516 28522 140522 28524
rect 193305 28522 193371 28525
rect 140516 28520 193371 28522
rect 140516 28464 193310 28520
rect 193366 28464 193371 28520
rect 140516 28462 193371 28464
rect 140516 28460 140522 28462
rect 193305 28459 193371 28462
rect 142838 28324 142844 28388
rect 142908 28386 142914 28388
rect 229093 28386 229159 28389
rect 142908 28384 229159 28386
rect 142908 28328 229098 28384
rect 229154 28328 229159 28384
rect 142908 28326 229159 28328
rect 142908 28324 142914 28326
rect 229093 28323 229159 28326
rect 165102 28188 165108 28252
rect 165172 28250 165178 28252
rect 514845 28250 514911 28253
rect 165172 28248 514911 28250
rect 165172 28192 514850 28248
rect 514906 28192 514911 28248
rect 165172 28190 514911 28192
rect 165172 28188 165178 28190
rect 514845 28187 514911 28190
rect 165286 26964 165292 27028
rect 165356 27026 165362 27028
rect 510613 27026 510679 27029
rect 165356 27024 510679 27026
rect 165356 26968 510618 27024
rect 510674 26968 510679 27024
rect 165356 26966 510679 26968
rect 165356 26964 165362 26966
rect 510613 26963 510679 26966
rect 170806 26828 170812 26892
rect 170876 26890 170882 26892
rect 576853 26890 576919 26893
rect 170876 26888 576919 26890
rect 170876 26832 576858 26888
rect 576914 26832 576919 26888
rect 170876 26830 576919 26832
rect 170876 26828 170882 26830
rect 576853 26827 576919 26830
rect 155534 25468 155540 25532
rect 155604 25530 155610 25532
rect 386413 25530 386479 25533
rect 155604 25528 386479 25530
rect 155604 25472 386418 25528
rect 386474 25472 386479 25528
rect 155604 25470 386479 25472
rect 155604 25468 155610 25470
rect 386413 25467 386479 25470
rect 157926 24108 157932 24172
rect 157996 24170 158002 24172
rect 422293 24170 422359 24173
rect 157996 24168 422359 24170
rect 157996 24112 422298 24168
rect 422354 24112 422359 24168
rect 157996 24110 422359 24112
rect 157996 24108 158002 24110
rect 422293 24107 422359 24110
rect 170438 21660 170444 21724
rect 170508 21722 170514 21724
rect 319437 21722 319503 21725
rect 170508 21720 319503 21722
rect 170508 21664 319442 21720
rect 319498 21664 319503 21720
rect 170508 21662 319503 21664
rect 170508 21660 170514 21662
rect 319437 21659 319503 21662
rect 158846 21524 158852 21588
rect 158916 21586 158922 21588
rect 442993 21586 443059 21589
rect 158916 21584 443059 21586
rect 158916 21528 442998 21584
rect 443054 21528 443059 21584
rect 158916 21526 443059 21528
rect 158916 21524 158922 21526
rect 442993 21523 443059 21526
rect 160870 21388 160876 21452
rect 160940 21450 160946 21452
rect 460933 21450 460999 21453
rect 160940 21448 460999 21450
rect 160940 21392 460938 21448
rect 460994 21392 460999 21448
rect 160940 21390 460999 21392
rect 160940 21388 160946 21390
rect 460933 21387 460999 21390
rect 162342 21252 162348 21316
rect 162412 21314 162418 21316
rect 476113 21314 476179 21317
rect 162412 21312 476179 21314
rect 162412 21256 476118 21312
rect 476174 21256 476179 21312
rect 162412 21254 476179 21256
rect 162412 21252 162418 21254
rect 476113 21251 476179 21254
rect 144494 20164 144500 20228
rect 144564 20226 144570 20228
rect 248413 20226 248479 20229
rect 144564 20224 248479 20226
rect 144564 20168 248418 20224
rect 248474 20168 248479 20224
rect 144564 20166 248479 20168
rect 144564 20164 144570 20166
rect 248413 20163 248479 20166
rect 161054 20028 161060 20092
rect 161124 20090 161130 20092
rect 458173 20090 458239 20093
rect 161124 20088 458239 20090
rect 161124 20032 458178 20088
rect 458234 20032 458239 20088
rect 161124 20030 458239 20032
rect 161124 20028 161130 20030
rect 458173 20027 458239 20030
rect 137686 19892 137692 19956
rect 137756 19954 137762 19956
rect 160553 19954 160619 19957
rect 137756 19952 160619 19954
rect 137756 19896 160558 19952
rect 160614 19896 160619 19952
rect 137756 19894 160619 19896
rect 137756 19892 137762 19894
rect 160553 19891 160619 19894
rect 163630 19892 163636 19956
rect 163700 19954 163706 19956
rect 495433 19954 495499 19957
rect 163700 19952 495499 19954
rect 163700 19896 495438 19952
rect 495494 19896 495499 19952
rect 163700 19894 495499 19896
rect 163700 19892 163706 19894
rect 495433 19891 495499 19894
rect 580165 19818 580231 19821
rect 583520 19818 584960 19908
rect 580165 19816 584960 19818
rect 580165 19760 580170 19816
rect 580226 19760 584960 19816
rect 580165 19758 584960 19760
rect 580165 19755 580231 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3877 19410 3943 19413
rect -960 19408 3943 19410
rect -960 19352 3882 19408
rect 3938 19352 3943 19408
rect -960 19350 3943 19352
rect -960 19260 480 19350
rect 3877 19347 3943 19350
rect 140078 18940 140084 19004
rect 140148 19002 140154 19004
rect 191833 19002 191899 19005
rect 140148 19000 191899 19002
rect 140148 18944 191838 19000
rect 191894 18944 191899 19000
rect 140148 18942 191899 18944
rect 140148 18940 140154 18942
rect 191833 18939 191899 18942
rect 152774 18804 152780 18868
rect 152844 18866 152850 18868
rect 350533 18866 350599 18869
rect 152844 18864 350599 18866
rect 152844 18808 350538 18864
rect 350594 18808 350599 18864
rect 152844 18806 350599 18808
rect 152844 18804 152850 18806
rect 350533 18803 350599 18806
rect 158110 18668 158116 18732
rect 158180 18730 158186 18732
rect 423673 18730 423739 18733
rect 158180 18728 423739 18730
rect 158180 18672 423678 18728
rect 423734 18672 423739 18728
rect 158180 18670 423739 18672
rect 158180 18668 158186 18670
rect 423673 18667 423739 18670
rect 167862 18532 167868 18596
rect 167932 18594 167938 18596
rect 547873 18594 547939 18597
rect 167932 18592 547939 18594
rect 167932 18536 547878 18592
rect 547934 18536 547939 18592
rect 167932 18534 547939 18536
rect 167932 18532 167938 18534
rect 547873 18531 547939 18534
rect 156822 17308 156828 17372
rect 156892 17370 156898 17372
rect 405733 17370 405799 17373
rect 156892 17368 405799 17370
rect 156892 17312 405738 17368
rect 405794 17312 405799 17368
rect 156892 17310 405799 17312
rect 156892 17308 156898 17310
rect 405733 17307 405799 17310
rect 161238 17172 161244 17236
rect 161308 17234 161314 17236
rect 456885 17234 456951 17237
rect 161308 17232 456951 17234
rect 161308 17176 456890 17232
rect 456946 17176 456951 17232
rect 161308 17174 456951 17176
rect 161308 17172 161314 17174
rect 456885 17171 456951 17174
rect 149830 16220 149836 16284
rect 149900 16282 149906 16284
rect 316217 16282 316283 16285
rect 149900 16280 316283 16282
rect 149900 16224 316222 16280
rect 316278 16224 316283 16280
rect 149900 16222 316283 16224
rect 149900 16220 149906 16222
rect 316217 16219 316283 16222
rect 154246 16084 154252 16148
rect 154316 16146 154322 16148
rect 371233 16146 371299 16149
rect 154316 16144 371299 16146
rect 154316 16088 371238 16144
rect 371294 16088 371299 16144
rect 154316 16086 371299 16088
rect 154316 16084 154322 16086
rect 371233 16083 371299 16086
rect 155718 15948 155724 16012
rect 155788 16010 155794 16012
rect 387793 16010 387859 16013
rect 155788 16008 387859 16010
rect 155788 15952 387798 16008
rect 387854 15952 387859 16008
rect 155788 15950 387859 15952
rect 155788 15948 155794 15950
rect 387793 15947 387859 15950
rect 158294 15812 158300 15876
rect 158364 15874 158370 15876
rect 420913 15874 420979 15877
rect 158364 15872 420979 15874
rect 158364 15816 420918 15872
rect 420974 15816 420979 15872
rect 158364 15814 420979 15816
rect 158364 15812 158370 15814
rect 420913 15811 420979 15814
rect 154430 14724 154436 14788
rect 154500 14786 154506 14788
rect 370129 14786 370195 14789
rect 154500 14784 370195 14786
rect 154500 14728 370134 14784
rect 370190 14728 370195 14784
rect 154500 14726 370195 14728
rect 154500 14724 154506 14726
rect 370129 14723 370195 14726
rect 157006 14588 157012 14652
rect 157076 14650 157082 14652
rect 407205 14650 407271 14653
rect 157076 14648 407271 14650
rect 157076 14592 407210 14648
rect 407266 14592 407271 14648
rect 157076 14590 407271 14592
rect 157076 14588 157082 14590
rect 407205 14587 407271 14590
rect 162526 14452 162532 14516
rect 162596 14514 162602 14516
rect 478137 14514 478203 14517
rect 162596 14512 478203 14514
rect 162596 14456 478142 14512
rect 478198 14456 478203 14512
rect 162596 14454 478203 14456
rect 162596 14452 162602 14454
rect 478137 14451 478203 14454
rect 148542 13228 148548 13292
rect 148612 13290 148618 13292
rect 301497 13290 301563 13293
rect 148612 13288 301563 13290
rect 148612 13232 301502 13288
rect 301558 13232 301563 13288
rect 148612 13230 301563 13232
rect 148612 13228 148618 13230
rect 301497 13227 301563 13230
rect 152406 13092 152412 13156
rect 152476 13154 152482 13156
rect 349245 13154 349311 13157
rect 152476 13152 349311 13154
rect 152476 13096 349250 13152
rect 349306 13096 349311 13152
rect 152476 13094 349311 13096
rect 152476 13092 152482 13094
rect 349245 13091 349311 13094
rect 166758 12956 166764 13020
rect 166828 13018 166834 13020
rect 531405 13018 531471 13021
rect 166828 13016 531471 13018
rect 166828 12960 531410 13016
rect 531466 12960 531471 13016
rect 166828 12958 531471 12960
rect 166828 12956 166834 12958
rect 531405 12955 531471 12958
rect 158478 11732 158484 11796
rect 158548 11794 158554 11796
rect 423765 11794 423831 11797
rect 158548 11792 423831 11794
rect 158548 11736 423770 11792
rect 423826 11736 423831 11792
rect 158548 11734 423831 11736
rect 158548 11732 158554 11734
rect 423765 11731 423831 11734
rect 162710 11596 162716 11660
rect 162780 11658 162786 11660
rect 474089 11658 474155 11661
rect 162780 11656 474155 11658
rect 162780 11600 474094 11656
rect 474150 11600 474155 11656
rect 162780 11598 474155 11600
rect 162780 11596 162786 11598
rect 474089 11595 474155 11598
rect 140998 10644 141004 10708
rect 141068 10706 141074 10708
rect 213361 10706 213427 10709
rect 141068 10704 213427 10706
rect 141068 10648 213366 10704
rect 213422 10648 213427 10704
rect 141068 10646 213427 10648
rect 141068 10644 141074 10646
rect 213361 10643 213427 10646
rect 147070 10508 147076 10572
rect 147140 10570 147146 10572
rect 281533 10570 281599 10573
rect 147140 10568 281599 10570
rect 147140 10512 281538 10568
rect 281594 10512 281599 10568
rect 147140 10510 281599 10512
rect 147140 10508 147146 10510
rect 281533 10507 281599 10510
rect 110505 10434 110571 10437
rect 134190 10434 134196 10436
rect 110505 10432 134196 10434
rect 110505 10376 110510 10432
rect 110566 10376 134196 10432
rect 110505 10374 134196 10376
rect 110505 10371 110571 10374
rect 134190 10372 134196 10374
rect 134260 10372 134266 10436
rect 148726 10372 148732 10436
rect 148796 10434 148802 10436
rect 299657 10434 299723 10437
rect 148796 10432 299723 10434
rect 148796 10376 299662 10432
rect 299718 10376 299723 10432
rect 148796 10374 299723 10376
rect 148796 10372 148802 10374
rect 299657 10371 299723 10374
rect 92473 10298 92539 10301
rect 133086 10298 133092 10300
rect 92473 10296 133092 10298
rect 92473 10240 92478 10296
rect 92534 10240 133092 10296
rect 92473 10238 133092 10240
rect 92473 10235 92539 10238
rect 133086 10236 133092 10238
rect 133156 10236 133162 10300
rect 164918 10236 164924 10300
rect 164988 10298 164994 10300
rect 513373 10298 513439 10301
rect 164988 10296 513439 10298
rect 164988 10240 513378 10296
rect 513434 10240 513439 10296
rect 164988 10238 513439 10240
rect 164988 10236 164994 10238
rect 513373 10235 513439 10238
rect 145414 9148 145420 9212
rect 145484 9210 145490 9212
rect 264145 9210 264211 9213
rect 145484 9208 264211 9210
rect 145484 9152 264150 9208
rect 264206 9152 264211 9208
rect 145484 9150 264211 9152
rect 145484 9148 145490 9150
rect 264145 9147 264211 9150
rect 78581 9074 78647 9077
rect 131430 9074 131436 9076
rect 78581 9072 131436 9074
rect 78581 9016 78586 9072
rect 78642 9016 131436 9072
rect 78581 9014 131436 9016
rect 78581 9011 78647 9014
rect 131430 9012 131436 9014
rect 131500 9012 131506 9076
rect 148910 9012 148916 9076
rect 148980 9074 148986 9076
rect 300761 9074 300827 9077
rect 148980 9072 300827 9074
rect 148980 9016 300766 9072
rect 300822 9016 300827 9072
rect 148980 9014 300827 9016
rect 148980 9012 148986 9014
rect 300761 9011 300827 9014
rect 57145 8938 57211 8941
rect 129958 8938 129964 8940
rect 57145 8936 129964 8938
rect 57145 8880 57150 8936
rect 57206 8880 129964 8936
rect 57145 8878 129964 8880
rect 57145 8875 57211 8878
rect 129958 8876 129964 8878
rect 130028 8876 130034 8940
rect 156638 8876 156644 8940
rect 156708 8938 156714 8940
rect 408401 8938 408467 8941
rect 156708 8936 408467 8938
rect 156708 8880 408406 8936
rect 408462 8880 408467 8936
rect 156708 8878 408467 8880
rect 156708 8876 156714 8878
rect 408401 8875 408467 8878
rect 109309 7986 109375 7989
rect 134006 7986 134012 7988
rect 109309 7984 134012 7986
rect 109309 7928 109314 7984
rect 109370 7928 134012 7984
rect 109309 7926 134012 7928
rect 109309 7923 109375 7926
rect 134006 7924 134012 7926
rect 134076 7924 134082 7988
rect 56041 7850 56107 7853
rect 130142 7850 130148 7852
rect 56041 7848 130148 7850
rect 56041 7792 56046 7848
rect 56102 7792 130148 7848
rect 56041 7790 130148 7792
rect 56041 7787 56107 7790
rect 130142 7788 130148 7790
rect 130212 7788 130218 7852
rect 41873 7714 41939 7717
rect 128670 7714 128676 7716
rect 41873 7712 128676 7714
rect 41873 7656 41878 7712
rect 41934 7656 128676 7712
rect 41873 7654 128676 7656
rect 41873 7651 41939 7654
rect 128670 7652 128676 7654
rect 128740 7652 128746 7716
rect 144126 7652 144132 7716
rect 144196 7714 144202 7716
rect 246389 7714 246455 7717
rect 144196 7712 246455 7714
rect 144196 7656 246394 7712
rect 246450 7656 246455 7712
rect 144196 7654 246455 7656
rect 144196 7652 144202 7654
rect 246389 7651 246455 7654
rect 38377 7578 38443 7581
rect 128854 7578 128860 7580
rect 38377 7576 128860 7578
rect 38377 7520 38382 7576
rect 38438 7520 128860 7576
rect 38377 7518 128860 7520
rect 38377 7515 38443 7518
rect 128854 7516 128860 7518
rect 128924 7516 128930 7580
rect 145598 7516 145604 7580
rect 145668 7578 145674 7580
rect 265341 7578 265407 7581
rect 145668 7576 265407 7578
rect 145668 7520 265346 7576
rect 265402 7520 265407 7576
rect 145668 7518 265407 7520
rect 145668 7516 145674 7518
rect 265341 7515 265407 7518
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 151302 6428 151308 6492
rect 151372 6490 151378 6492
rect 336273 6490 336339 6493
rect 151372 6488 336339 6490
rect 151372 6432 336278 6488
rect 336334 6432 336339 6488
rect 583520 6476 584960 6566
rect 151372 6430 336339 6432
rect 151372 6428 151378 6430
rect 336273 6427 336339 6430
rect 111609 6354 111675 6357
rect 133822 6354 133828 6356
rect 111609 6352 133828 6354
rect 111609 6296 111614 6352
rect 111670 6296 133828 6352
rect 111609 6294 133828 6296
rect 111609 6291 111675 6294
rect 133822 6292 133828 6294
rect 133892 6292 133898 6356
rect 151486 6292 151492 6356
rect 151556 6354 151562 6356
rect 337469 6354 337535 6357
rect 151556 6352 337535 6354
rect 151556 6296 337474 6352
rect 337530 6296 337535 6352
rect 151556 6294 337535 6296
rect 151556 6292 151562 6294
rect 337469 6291 337535 6294
rect 73797 6218 73863 6221
rect 131246 6218 131252 6220
rect 73797 6216 131252 6218
rect 73797 6160 73802 6216
rect 73858 6160 131252 6216
rect 73797 6158 131252 6160
rect 73797 6155 73863 6158
rect 131246 6156 131252 6158
rect 131316 6156 131322 6220
rect 131982 6156 131988 6220
rect 132052 6218 132058 6220
rect 333881 6218 333947 6221
rect 132052 6216 333947 6218
rect 132052 6160 333886 6216
rect 333942 6160 333947 6216
rect 132052 6158 333947 6160
rect 132052 6156 132058 6158
rect 333881 6155 333947 6158
rect 150014 5068 150020 5132
rect 150084 5130 150090 5132
rect 315021 5130 315087 5133
rect 150084 5128 315087 5130
rect 150084 5072 315026 5128
rect 315082 5072 315087 5128
rect 150084 5070 315087 5072
rect 150084 5068 150090 5070
rect 315021 5067 315087 5070
rect 159030 4932 159036 4996
rect 159100 4994 159106 4996
rect 442625 4994 442691 4997
rect 159100 4992 442691 4994
rect 159100 4936 442630 4992
rect 442686 4936 442691 4992
rect 159100 4934 442691 4936
rect 159100 4932 159106 4934
rect 442625 4931 442691 4934
rect 4061 4858 4127 4861
rect 125910 4858 125916 4860
rect 4061 4856 125916 4858
rect 4061 4800 4066 4856
rect 4122 4800 125916 4856
rect 4061 4798 125916 4800
rect 4061 4795 4127 4798
rect 125910 4796 125916 4798
rect 125980 4796 125986 4860
rect 137870 4796 137876 4860
rect 137940 4858 137946 4860
rect 158897 4858 158963 4861
rect 137940 4856 158963 4858
rect 137940 4800 158902 4856
rect 158958 4800 158963 4856
rect 137940 4798 158963 4800
rect 137940 4796 137946 4798
rect 158897 4795 158963 4798
rect 168046 4796 168052 4860
rect 168116 4858 168122 4860
rect 547873 4858 547939 4861
rect 168116 4856 547939 4858
rect 168116 4800 547878 4856
rect 547934 4800 547939 4856
rect 168116 4798 547939 4800
rect 168116 4796 168122 4798
rect 547873 4795 547939 4798
rect 151670 3572 151676 3636
rect 151740 3634 151746 3636
rect 335077 3634 335143 3637
rect 151740 3632 335143 3634
rect 151740 3576 335082 3632
rect 335138 3576 335143 3632
rect 151740 3574 335143 3576
rect 151740 3572 151746 3574
rect 335077 3571 335143 3574
rect 72601 3498 72667 3501
rect 131062 3498 131068 3500
rect 72601 3496 131068 3498
rect 72601 3440 72606 3496
rect 72662 3440 131068 3496
rect 72601 3438 131068 3440
rect 72601 3435 72667 3438
rect 131062 3436 131068 3438
rect 131132 3436 131138 3500
rect 171726 3436 171732 3500
rect 171796 3498 171802 3500
rect 570321 3498 570387 3501
rect 171796 3496 570387 3498
rect 171796 3440 570326 3496
rect 570382 3440 570387 3496
rect 171796 3438 570387 3440
rect 171796 3436 171802 3438
rect 570321 3435 570387 3438
rect 20621 3362 20687 3365
rect 127382 3362 127388 3364
rect 20621 3360 127388 3362
rect 20621 3304 20626 3360
rect 20682 3304 127388 3360
rect 20621 3302 127388 3304
rect 20621 3299 20687 3302
rect 127382 3300 127388 3302
rect 127452 3300 127458 3364
rect 136398 3300 136404 3364
rect 136468 3362 136474 3364
rect 161289 3362 161355 3365
rect 136468 3360 161355 3362
rect 136468 3304 161294 3360
rect 161350 3304 161355 3360
rect 136468 3302 161355 3304
rect 136468 3300 136474 3302
rect 161289 3299 161355 3302
rect 171910 3300 171916 3364
rect 171980 3362 171986 3364
rect 580993 3362 581059 3365
rect 171980 3360 581059 3362
rect 171980 3304 580998 3360
rect 581054 3304 581059 3360
rect 171980 3302 581059 3304
rect 171980 3300 171986 3302
rect 580993 3299 581059 3302
<< via3 >>
rect 396580 696900 396644 696964
rect 396764 643180 396828 643244
rect 144500 191040 144564 191044
rect 144500 190984 144514 191040
rect 144514 190984 144564 191040
rect 144500 190980 144564 190984
rect 146156 188532 146220 188596
rect 144500 185948 144564 186012
rect 146340 185948 146404 186012
rect 142844 184316 142908 184380
rect 141004 184180 141068 184244
rect 143028 184044 143092 184108
rect 142476 181052 142540 181116
rect 143028 178876 143092 178940
rect 141004 178740 141068 178804
rect 142844 178740 142908 178804
rect 158484 176428 158548 176492
rect 146340 175340 146404 175404
rect 142476 172952 142540 172956
rect 142476 172896 142526 172952
rect 142526 172896 142540 172952
rect 142476 172892 142540 172896
rect 158484 172952 158548 172956
rect 158484 172896 158498 172952
rect 158498 172896 158548 172952
rect 158484 172892 158548 172896
rect 146156 142700 146220 142764
rect 173572 81228 173636 81292
rect 171548 81092 171612 81156
rect 171180 80684 171244 80748
rect 166212 80548 166276 80612
rect 171364 80548 171428 80612
rect 173204 80412 173268 80476
rect 131804 80140 131868 80204
rect 142844 80140 142908 80204
rect 159220 80140 159284 80204
rect 166212 80140 166276 80204
rect 125732 79928 125796 79932
rect 125732 79872 125736 79928
rect 125736 79872 125792 79928
rect 125792 79872 125796 79928
rect 125732 79868 125796 79872
rect 125916 79868 125980 79932
rect 128492 79868 128556 79932
rect 129044 79928 129108 79932
rect 129044 79872 129048 79928
rect 129048 79872 129104 79928
rect 129104 79872 129108 79928
rect 129044 79868 129108 79872
rect 127388 79656 127452 79660
rect 129964 79906 129968 79932
rect 129968 79906 130024 79932
rect 130024 79906 130028 79932
rect 129964 79868 130028 79906
rect 131620 79906 131624 79932
rect 131624 79906 131680 79932
rect 131680 79906 131684 79932
rect 131620 79868 131684 79906
rect 127388 79600 127402 79656
rect 127402 79600 127452 79656
rect 127388 79596 127452 79600
rect 130884 79732 130948 79796
rect 128860 79596 128924 79660
rect 129780 79596 129844 79660
rect 133460 79868 133524 79932
rect 134012 79928 134076 79932
rect 134012 79872 134016 79928
rect 134016 79872 134072 79928
rect 134072 79872 134076 79928
rect 134012 79868 134076 79872
rect 133092 79732 133156 79796
rect 133276 79732 133340 79796
rect 134564 79868 134628 79932
rect 135484 79928 135548 79932
rect 135484 79872 135488 79928
rect 135488 79872 135544 79928
rect 135544 79872 135548 79928
rect 135484 79868 135548 79872
rect 136404 79906 136408 79932
rect 136408 79906 136464 79932
rect 136464 79906 136468 79932
rect 136404 79868 136468 79906
rect 136956 79868 137020 79932
rect 138060 79868 138124 79932
rect 140268 79868 140332 79932
rect 138796 79732 138860 79796
rect 139164 79792 139228 79796
rect 139164 79736 139178 79792
rect 139178 79736 139228 79792
rect 139164 79732 139228 79736
rect 140084 79732 140148 79796
rect 144500 79868 144564 79932
rect 145604 79868 145668 79932
rect 146708 79906 146712 79932
rect 146712 79906 146768 79932
rect 146768 79906 146772 79932
rect 146708 79868 146772 79906
rect 147076 79928 147140 79932
rect 147076 79872 147080 79928
rect 147080 79872 147136 79928
rect 147136 79872 147140 79928
rect 147076 79868 147140 79872
rect 147812 79928 147876 79932
rect 147812 79872 147816 79928
rect 147816 79872 147872 79928
rect 147872 79872 147876 79928
rect 147812 79868 147876 79872
rect 148916 79906 148920 79932
rect 148920 79906 148976 79932
rect 148976 79906 148980 79932
rect 148916 79868 148980 79906
rect 144316 79596 144380 79660
rect 146156 79656 146220 79660
rect 146156 79600 146206 79656
rect 146206 79600 146220 79656
rect 146156 79596 146220 79600
rect 149652 79868 149716 79932
rect 151676 79868 151740 79932
rect 149836 79732 149900 79796
rect 151492 79732 151556 79796
rect 152780 79928 152844 79932
rect 152780 79872 152784 79928
rect 152784 79872 152840 79928
rect 152840 79872 152844 79928
rect 152780 79868 152844 79872
rect 154068 79928 154132 79932
rect 154068 79872 154072 79928
rect 154072 79872 154128 79928
rect 154128 79872 154132 79928
rect 154068 79868 154132 79872
rect 154252 79868 154316 79932
rect 154988 79868 155052 79932
rect 155724 79928 155788 79932
rect 155724 79872 155728 79928
rect 155728 79872 155784 79928
rect 155784 79872 155788 79928
rect 153884 79732 153948 79796
rect 155724 79868 155788 79872
rect 156092 79928 156156 79932
rect 156092 79872 156096 79928
rect 156096 79872 156152 79928
rect 156152 79872 156156 79928
rect 156092 79868 156156 79872
rect 156828 79868 156892 79932
rect 157748 79928 157812 79932
rect 157748 79872 157752 79928
rect 157752 79872 157808 79928
rect 157808 79872 157812 79928
rect 157748 79868 157812 79872
rect 158116 79868 158180 79932
rect 157012 79732 157076 79796
rect 158300 79792 158364 79796
rect 158300 79736 158304 79792
rect 158304 79736 158360 79792
rect 158360 79736 158364 79792
rect 158300 79732 158364 79736
rect 159036 79732 159100 79796
rect 161244 79928 161308 79932
rect 161244 79872 161248 79928
rect 161248 79872 161304 79928
rect 161304 79872 161308 79928
rect 161244 79868 161308 79872
rect 162716 79868 162780 79932
rect 163452 79868 163516 79932
rect 164924 79928 164988 79932
rect 164924 79872 164928 79928
rect 164928 79872 164984 79928
rect 164984 79872 164988 79928
rect 164924 79868 164988 79872
rect 165108 79868 165172 79932
rect 160140 79596 160204 79660
rect 162348 79732 162412 79796
rect 162532 79596 162596 79660
rect 164372 79596 164436 79660
rect 165292 79792 165356 79796
rect 165292 79736 165296 79792
rect 165296 79736 165352 79792
rect 165352 79736 165356 79792
rect 165292 79732 165356 79736
rect 166396 79868 166460 79932
rect 167500 79906 167504 79932
rect 167504 79906 167560 79932
rect 167560 79906 167564 79932
rect 167500 79868 167564 79906
rect 169156 79868 169220 79932
rect 169340 79928 169404 79932
rect 169340 79872 169344 79928
rect 169344 79872 169400 79928
rect 169400 79872 169404 79928
rect 169340 79868 169404 79872
rect 166580 79732 166644 79796
rect 167868 79596 167932 79660
rect 170444 79868 170508 79932
rect 171180 79868 171244 79932
rect 171916 79928 171980 79932
rect 171916 79872 171920 79928
rect 171920 79872 171976 79928
rect 171976 79872 171980 79928
rect 171916 79868 171980 79872
rect 172422 79928 172486 79932
rect 172422 79872 172436 79928
rect 172436 79872 172486 79928
rect 172422 79868 172486 79872
rect 171364 79732 171428 79796
rect 170628 79596 170692 79660
rect 173572 79656 173636 79660
rect 173572 79600 173622 79656
rect 173622 79600 173636 79656
rect 173572 79596 173636 79600
rect 173204 79460 173268 79524
rect 159220 79052 159284 79116
rect 161244 79052 161308 79116
rect 163636 79052 163700 79116
rect 125916 78780 125980 78844
rect 128676 78780 128740 78844
rect 130332 78780 130396 78844
rect 131620 78780 131684 78844
rect 144316 78840 144380 78844
rect 144316 78784 144366 78840
rect 144366 78784 144380 78840
rect 144316 78780 144380 78784
rect 146156 78780 146220 78844
rect 125916 78704 125980 78708
rect 125916 78648 125930 78704
rect 125930 78648 125980 78704
rect 125916 78644 125980 78648
rect 130148 78644 130212 78708
rect 138980 78644 139044 78708
rect 150020 78704 150084 78708
rect 171548 78780 171612 78844
rect 171916 78916 171980 78980
rect 150020 78648 150034 78704
rect 150034 78648 150084 78704
rect 150020 78644 150084 78648
rect 167684 78644 167748 78708
rect 170076 78704 170140 78708
rect 170076 78648 170126 78704
rect 170126 78648 170140 78704
rect 170076 78644 170140 78648
rect 170996 78704 171060 78708
rect 170996 78648 171010 78704
rect 171010 78648 171060 78704
rect 170996 78644 171060 78648
rect 172468 78644 172532 78708
rect 129044 78508 129108 78572
rect 130884 78508 130948 78572
rect 145236 78508 145300 78572
rect 149468 78508 149532 78572
rect 160140 78508 160204 78572
rect 131436 78372 131500 78436
rect 148548 78372 148612 78436
rect 136956 78160 137020 78164
rect 136956 78104 136970 78160
rect 136970 78104 137020 78160
rect 136956 78100 137020 78104
rect 154988 78160 155052 78164
rect 154988 78104 155038 78160
rect 155038 78104 155052 78160
rect 154988 78100 155052 78104
rect 146708 78024 146772 78028
rect 146708 77968 146722 78024
rect 146722 77968 146772 78024
rect 146708 77964 146772 77968
rect 147076 77964 147140 78028
rect 147260 78024 147324 78028
rect 147260 77968 147310 78024
rect 147310 77968 147324 78024
rect 147260 77964 147324 77968
rect 396764 78372 396828 78436
rect 396580 78100 396644 78164
rect 148364 77828 148428 77892
rect 131988 77692 132052 77756
rect 127388 77556 127452 77620
rect 127388 77420 127452 77484
rect 127204 77344 127268 77348
rect 127204 77288 127254 77344
rect 127254 77288 127268 77344
rect 127204 77284 127268 77288
rect 147076 77284 147140 77348
rect 161244 77284 161308 77348
rect 169156 77284 169220 77348
rect 171180 77284 171244 77348
rect 131252 77072 131316 77076
rect 131252 77016 131302 77072
rect 131302 77016 131316 77072
rect 131252 77012 131316 77016
rect 133828 77012 133892 77076
rect 152596 77012 152660 77076
rect 133276 76876 133340 76940
rect 131804 76740 131868 76804
rect 137692 76740 137756 76804
rect 133460 76604 133524 76668
rect 134196 76604 134260 76668
rect 134564 76664 134628 76668
rect 134564 76608 134614 76664
rect 134614 76608 134628 76664
rect 134564 76604 134628 76608
rect 136404 76604 136468 76668
rect 137876 76664 137940 76668
rect 137876 76608 137926 76664
rect 137926 76608 137940 76664
rect 137876 76604 137940 76608
rect 138060 76604 138124 76668
rect 151676 76664 151740 76668
rect 151676 76608 151690 76664
rect 151690 76608 151740 76664
rect 151676 76604 151740 76608
rect 152964 76664 153028 76668
rect 152964 76608 153014 76664
rect 153014 76608 153028 76664
rect 152964 76604 153028 76608
rect 154068 76604 154132 76668
rect 154436 76664 154500 76668
rect 154436 76608 154450 76664
rect 154450 76608 154500 76664
rect 154436 76604 154500 76608
rect 155540 76664 155604 76668
rect 155540 76608 155590 76664
rect 155590 76608 155604 76664
rect 155540 76604 155604 76608
rect 156092 76604 156156 76668
rect 156644 76604 156708 76668
rect 157748 76604 157812 76668
rect 158484 76664 158548 76668
rect 158484 76608 158534 76664
rect 158534 76608 158548 76664
rect 158484 76604 158548 76608
rect 160876 76604 160940 76668
rect 164924 76604 164988 76668
rect 165476 76664 165540 76668
rect 165476 76608 165490 76664
rect 165490 76608 165540 76664
rect 165476 76604 165540 76608
rect 166764 76664 166828 76668
rect 166764 76608 166814 76664
rect 166814 76608 166828 76664
rect 166764 76604 166828 76608
rect 168052 76604 168116 76668
rect 136404 76468 136468 76532
rect 151308 76468 151372 76532
rect 152780 76528 152844 76532
rect 152780 76472 152830 76528
rect 152830 76472 152844 76528
rect 152780 76468 152844 76472
rect 154068 76468 154132 76532
rect 157932 76468 157996 76532
rect 160692 76468 160756 76532
rect 164924 76468 164988 76532
rect 169340 76468 169404 76532
rect 140452 76332 140516 76396
rect 151860 76332 151924 76396
rect 161060 76332 161124 76396
rect 167500 76392 167564 76396
rect 167500 76336 167550 76392
rect 167550 76336 167564 76392
rect 167500 76332 167564 76336
rect 158852 76196 158916 76260
rect 170812 76196 170876 76260
rect 144132 76060 144196 76124
rect 169340 76060 169404 76124
rect 170996 76060 171060 76124
rect 141004 75924 141068 75988
rect 143212 75984 143276 75988
rect 143212 75928 143262 75984
rect 143262 75928 143276 75984
rect 143212 75924 143276 75928
rect 145420 75924 145484 75988
rect 147812 75984 147876 75988
rect 147812 75928 147862 75984
rect 147862 75928 147876 75984
rect 147812 75924 147876 75928
rect 148732 75924 148796 75988
rect 171732 75924 171796 75988
rect 133276 75788 133340 75852
rect 143028 75788 143092 75852
rect 170076 75788 170140 75852
rect 171916 75788 171980 75852
rect 139164 75652 139228 75716
rect 130332 75516 130396 75580
rect 129780 75380 129844 75444
rect 164556 75244 164620 75308
rect 125732 75108 125796 75172
rect 128860 73748 128924 73812
rect 131068 73204 131132 73268
rect 148364 72388 148428 72452
rect 152964 71164 153028 71228
rect 163452 71028 163516 71092
rect 138980 69532 139044 69596
rect 165476 68172 165540 68236
rect 140268 65452 140332 65516
rect 166396 62868 166460 62932
rect 171180 62732 171244 62796
rect 160692 61372 160756 61436
rect 138796 60012 138860 60076
rect 143028 59876 143092 59940
rect 149468 53076 149532 53140
rect 152596 47500 152660 47564
rect 135300 44916 135364 44980
rect 133276 44780 133340 44844
rect 147260 44780 147324 44844
rect 127204 43420 127268 43484
rect 153884 40564 153948 40628
rect 154068 35124 154132 35188
rect 143212 34036 143276 34100
rect 145236 33900 145300 33964
rect 170628 33764 170692 33828
rect 166580 32540 166644 32604
rect 169340 32404 169404 32468
rect 167684 30908 167748 30972
rect 149652 29548 149716 29612
rect 140452 28460 140516 28524
rect 142844 28324 142908 28388
rect 165108 28188 165172 28252
rect 165292 26964 165356 27028
rect 170812 26828 170876 26892
rect 155540 25468 155604 25532
rect 157932 24108 157996 24172
rect 170444 21660 170508 21724
rect 158852 21524 158916 21588
rect 160876 21388 160940 21452
rect 162348 21252 162412 21316
rect 144500 20164 144564 20228
rect 161060 20028 161124 20092
rect 137692 19892 137756 19956
rect 163636 19892 163700 19956
rect 140084 18940 140148 19004
rect 152780 18804 152844 18868
rect 158116 18668 158180 18732
rect 167868 18532 167932 18596
rect 156828 17308 156892 17372
rect 161244 17172 161308 17236
rect 149836 16220 149900 16284
rect 154252 16084 154316 16148
rect 155724 15948 155788 16012
rect 158300 15812 158364 15876
rect 154436 14724 154500 14788
rect 157012 14588 157076 14652
rect 162532 14452 162596 14516
rect 148548 13228 148612 13292
rect 152412 13092 152476 13156
rect 166764 12956 166828 13020
rect 158484 11732 158548 11796
rect 162716 11596 162780 11660
rect 141004 10644 141068 10708
rect 147076 10508 147140 10572
rect 134196 10372 134260 10436
rect 148732 10372 148796 10436
rect 133092 10236 133156 10300
rect 164924 10236 164988 10300
rect 145420 9148 145484 9212
rect 131436 9012 131500 9076
rect 148916 9012 148980 9076
rect 129964 8876 130028 8940
rect 156644 8876 156708 8940
rect 134012 7924 134076 7988
rect 130148 7788 130212 7852
rect 128676 7652 128740 7716
rect 144132 7652 144196 7716
rect 128860 7516 128924 7580
rect 145604 7516 145668 7580
rect 151308 6428 151372 6492
rect 133828 6292 133892 6356
rect 151492 6292 151556 6356
rect 131252 6156 131316 6220
rect 131988 6156 132052 6220
rect 150020 5068 150084 5132
rect 159036 4932 159100 4996
rect 125916 4796 125980 4860
rect 137876 4796 137940 4860
rect 168052 4796 168116 4860
rect 151676 3572 151740 3636
rect 131068 3436 131132 3500
rect 171732 3436 171796 3500
rect 127388 3300 127452 3364
rect 136404 3300 136468 3364
rect 171916 3300 171980 3364
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 682954 -8106 711002
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 -8106 682954
rect -8726 682634 -8106 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 -8106 682634
rect -8726 646954 -8106 682398
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 -8106 646954
rect -8726 646634 -8106 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 -8106 646634
rect -8726 610954 -8106 646398
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 -8106 610954
rect -8726 610634 -8106 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 -8106 610634
rect -8726 574954 -8106 610398
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 -8106 574954
rect -8726 574634 -8106 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 -8106 574634
rect -8726 538954 -8106 574398
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 -8106 538954
rect -8726 538634 -8106 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 -8106 538634
rect -8726 502954 -8106 538398
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 -8106 502954
rect -8726 502634 -8106 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 -8106 502634
rect -8726 466954 -8106 502398
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 -8106 466954
rect -8726 466634 -8106 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 -8106 466634
rect -8726 430954 -8106 466398
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 -8106 430954
rect -8726 430634 -8106 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 -8106 430634
rect -8726 394954 -8106 430398
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 -8106 394954
rect -8726 394634 -8106 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 -8106 394634
rect -8726 358954 -8106 394398
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 -8106 358954
rect -8726 358634 -8106 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 -8106 358634
rect -8726 322954 -8106 358398
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 -8106 322954
rect -8726 322634 -8106 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 -8106 322634
rect -8726 286954 -8106 322398
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 -8106 286954
rect -8726 286634 -8106 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 -8106 286634
rect -8726 250954 -8106 286398
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 -8106 250954
rect -8726 250634 -8106 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 -8106 250634
rect -8726 214954 -8106 250398
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 -8106 214954
rect -8726 214634 -8106 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 -8106 214634
rect -8726 178954 -8106 214398
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 -8106 178954
rect -8726 178634 -8106 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 -8106 178634
rect -8726 142954 -8106 178398
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 -8106 142954
rect -8726 142634 -8106 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 -8106 142634
rect -8726 106954 -8106 142398
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 -8106 106954
rect -8726 106634 -8106 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 -8106 106634
rect -8726 70954 -8106 106398
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 -8106 70954
rect -8726 70634 -8106 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 -8106 70634
rect -8726 34954 -8106 70398
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 -8106 34954
rect -8726 34634 -8106 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 -8106 34634
rect -8726 -7066 -8106 34398
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 678454 -7146 710042
rect -7766 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 -7146 678454
rect -7766 678134 -7146 678218
rect -7766 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 -7146 678134
rect -7766 642454 -7146 677898
rect -7766 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 -7146 642454
rect -7766 642134 -7146 642218
rect -7766 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 -7146 642134
rect -7766 606454 -7146 641898
rect -7766 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 -7146 606454
rect -7766 606134 -7146 606218
rect -7766 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 -7146 606134
rect -7766 570454 -7146 605898
rect -7766 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 -7146 570454
rect -7766 570134 -7146 570218
rect -7766 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 -7146 570134
rect -7766 534454 -7146 569898
rect -7766 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 -7146 534454
rect -7766 534134 -7146 534218
rect -7766 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 -7146 534134
rect -7766 498454 -7146 533898
rect -7766 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 -7146 498454
rect -7766 498134 -7146 498218
rect -7766 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 -7146 498134
rect -7766 462454 -7146 497898
rect -7766 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 -7146 462454
rect -7766 462134 -7146 462218
rect -7766 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 -7146 462134
rect -7766 426454 -7146 461898
rect -7766 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 -7146 426454
rect -7766 426134 -7146 426218
rect -7766 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 -7146 426134
rect -7766 390454 -7146 425898
rect -7766 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 -7146 390454
rect -7766 390134 -7146 390218
rect -7766 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 -7146 390134
rect -7766 354454 -7146 389898
rect -7766 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 -7146 354454
rect -7766 354134 -7146 354218
rect -7766 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 -7146 354134
rect -7766 318454 -7146 353898
rect -7766 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 -7146 318454
rect -7766 318134 -7146 318218
rect -7766 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 -7146 318134
rect -7766 282454 -7146 317898
rect -7766 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 -7146 282454
rect -7766 282134 -7146 282218
rect -7766 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 -7146 282134
rect -7766 246454 -7146 281898
rect -7766 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 -7146 246454
rect -7766 246134 -7146 246218
rect -7766 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 -7146 246134
rect -7766 210454 -7146 245898
rect -7766 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 -7146 210454
rect -7766 210134 -7146 210218
rect -7766 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 -7146 210134
rect -7766 174454 -7146 209898
rect -7766 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 -7146 174454
rect -7766 174134 -7146 174218
rect -7766 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 -7146 174134
rect -7766 138454 -7146 173898
rect -7766 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 -7146 138454
rect -7766 138134 -7146 138218
rect -7766 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 -7146 138134
rect -7766 102454 -7146 137898
rect -7766 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 -7146 102454
rect -7766 102134 -7146 102218
rect -7766 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 -7146 102134
rect -7766 66454 -7146 101898
rect -7766 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 -7146 66454
rect -7766 66134 -7146 66218
rect -7766 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 -7146 66134
rect -7766 30454 -7146 65898
rect -7766 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 -7146 30454
rect -7766 30134 -7146 30218
rect -7766 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 -7146 30134
rect -7766 -6106 -7146 29898
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 673954 -6186 709082
rect -6806 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 -6186 673954
rect -6806 673634 -6186 673718
rect -6806 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 -6186 673634
rect -6806 637954 -6186 673398
rect -6806 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 -6186 637954
rect -6806 637634 -6186 637718
rect -6806 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 -6186 637634
rect -6806 601954 -6186 637398
rect -6806 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 -6186 601954
rect -6806 601634 -6186 601718
rect -6806 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 -6186 601634
rect -6806 565954 -6186 601398
rect -6806 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 -6186 565954
rect -6806 565634 -6186 565718
rect -6806 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 -6186 565634
rect -6806 529954 -6186 565398
rect -6806 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 -6186 529954
rect -6806 529634 -6186 529718
rect -6806 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 -6186 529634
rect -6806 493954 -6186 529398
rect -6806 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 -6186 493954
rect -6806 493634 -6186 493718
rect -6806 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 -6186 493634
rect -6806 457954 -6186 493398
rect -6806 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 -6186 457954
rect -6806 457634 -6186 457718
rect -6806 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 -6186 457634
rect -6806 421954 -6186 457398
rect -6806 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 -6186 421954
rect -6806 421634 -6186 421718
rect -6806 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 -6186 421634
rect -6806 385954 -6186 421398
rect -6806 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 -6186 385954
rect -6806 385634 -6186 385718
rect -6806 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 -6186 385634
rect -6806 349954 -6186 385398
rect -6806 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 -6186 349954
rect -6806 349634 -6186 349718
rect -6806 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 -6186 349634
rect -6806 313954 -6186 349398
rect -6806 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 -6186 313954
rect -6806 313634 -6186 313718
rect -6806 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 -6186 313634
rect -6806 277954 -6186 313398
rect -6806 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 -6186 277954
rect -6806 277634 -6186 277718
rect -6806 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 -6186 277634
rect -6806 241954 -6186 277398
rect -6806 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 -6186 241954
rect -6806 241634 -6186 241718
rect -6806 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 -6186 241634
rect -6806 205954 -6186 241398
rect -6806 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 -6186 205954
rect -6806 205634 -6186 205718
rect -6806 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 -6186 205634
rect -6806 169954 -6186 205398
rect -6806 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 -6186 169954
rect -6806 169634 -6186 169718
rect -6806 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 -6186 169634
rect -6806 133954 -6186 169398
rect -6806 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 -6186 133954
rect -6806 133634 -6186 133718
rect -6806 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 -6186 133634
rect -6806 97954 -6186 133398
rect -6806 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 -6186 97954
rect -6806 97634 -6186 97718
rect -6806 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 -6186 97634
rect -6806 61954 -6186 97398
rect -6806 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 -6186 61954
rect -6806 61634 -6186 61718
rect -6806 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 -6186 61634
rect -6806 25954 -6186 61398
rect -6806 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 -6186 25954
rect -6806 25634 -6186 25718
rect -6806 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 -6186 25634
rect -6806 -5146 -6186 25398
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 669454 -5226 708122
rect -5846 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 -5226 669454
rect -5846 669134 -5226 669218
rect -5846 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 -5226 669134
rect -5846 633454 -5226 668898
rect -5846 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 -5226 633454
rect -5846 633134 -5226 633218
rect -5846 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 -5226 633134
rect -5846 597454 -5226 632898
rect -5846 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 -5226 597454
rect -5846 597134 -5226 597218
rect -5846 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 -5226 597134
rect -5846 561454 -5226 596898
rect -5846 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 -5226 561454
rect -5846 561134 -5226 561218
rect -5846 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 -5226 561134
rect -5846 525454 -5226 560898
rect -5846 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 -5226 525454
rect -5846 525134 -5226 525218
rect -5846 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 -5226 525134
rect -5846 489454 -5226 524898
rect -5846 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 -5226 489454
rect -5846 489134 -5226 489218
rect -5846 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 -5226 489134
rect -5846 453454 -5226 488898
rect -5846 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 -5226 453454
rect -5846 453134 -5226 453218
rect -5846 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 -5226 453134
rect -5846 417454 -5226 452898
rect -5846 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 -5226 417454
rect -5846 417134 -5226 417218
rect -5846 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 -5226 417134
rect -5846 381454 -5226 416898
rect -5846 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 -5226 381454
rect -5846 381134 -5226 381218
rect -5846 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 -5226 381134
rect -5846 345454 -5226 380898
rect -5846 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 -5226 345454
rect -5846 345134 -5226 345218
rect -5846 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 -5226 345134
rect -5846 309454 -5226 344898
rect -5846 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 -5226 309454
rect -5846 309134 -5226 309218
rect -5846 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 -5226 309134
rect -5846 273454 -5226 308898
rect -5846 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 -5226 273454
rect -5846 273134 -5226 273218
rect -5846 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 -5226 273134
rect -5846 237454 -5226 272898
rect -5846 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 -5226 237454
rect -5846 237134 -5226 237218
rect -5846 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 -5226 237134
rect -5846 201454 -5226 236898
rect -5846 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 -5226 201454
rect -5846 201134 -5226 201218
rect -5846 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 -5226 201134
rect -5846 165454 -5226 200898
rect -5846 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 -5226 165454
rect -5846 165134 -5226 165218
rect -5846 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 -5226 165134
rect -5846 129454 -5226 164898
rect -5846 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 -5226 129454
rect -5846 129134 -5226 129218
rect -5846 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 -5226 129134
rect -5846 93454 -5226 128898
rect -5846 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 -5226 93454
rect -5846 93134 -5226 93218
rect -5846 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 -5226 93134
rect -5846 57454 -5226 92898
rect -5846 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 -5226 57454
rect -5846 57134 -5226 57218
rect -5846 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 -5226 57134
rect -5846 21454 -5226 56898
rect -5846 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 -5226 21454
rect -5846 21134 -5226 21218
rect -5846 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 -5226 21134
rect -5846 -4186 -5226 20898
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 700954 -4266 707162
rect -4886 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 -4266 700954
rect -4886 700634 -4266 700718
rect -4886 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 -4266 700634
rect -4886 664954 -4266 700398
rect -4886 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 -4266 664954
rect -4886 664634 -4266 664718
rect -4886 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 -4266 664634
rect -4886 628954 -4266 664398
rect -4886 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 -4266 628954
rect -4886 628634 -4266 628718
rect -4886 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 -4266 628634
rect -4886 592954 -4266 628398
rect -4886 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 -4266 592954
rect -4886 592634 -4266 592718
rect -4886 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 -4266 592634
rect -4886 556954 -4266 592398
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 -4266 556954
rect -4886 556634 -4266 556718
rect -4886 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 -4266 556634
rect -4886 520954 -4266 556398
rect -4886 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 -4266 520954
rect -4886 520634 -4266 520718
rect -4886 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 -4266 520634
rect -4886 484954 -4266 520398
rect -4886 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 -4266 484954
rect -4886 484634 -4266 484718
rect -4886 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 -4266 484634
rect -4886 448954 -4266 484398
rect -4886 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 -4266 448954
rect -4886 448634 -4266 448718
rect -4886 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 -4266 448634
rect -4886 412954 -4266 448398
rect -4886 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 -4266 412954
rect -4886 412634 -4266 412718
rect -4886 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 -4266 412634
rect -4886 376954 -4266 412398
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 -4266 376954
rect -4886 376634 -4266 376718
rect -4886 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 -4266 376634
rect -4886 340954 -4266 376398
rect -4886 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 -4266 340954
rect -4886 340634 -4266 340718
rect -4886 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 -4266 340634
rect -4886 304954 -4266 340398
rect -4886 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 -4266 304954
rect -4886 304634 -4266 304718
rect -4886 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 -4266 304634
rect -4886 268954 -4266 304398
rect -4886 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 -4266 268954
rect -4886 268634 -4266 268718
rect -4886 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 -4266 268634
rect -4886 232954 -4266 268398
rect -4886 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 -4266 232954
rect -4886 232634 -4266 232718
rect -4886 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 -4266 232634
rect -4886 196954 -4266 232398
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 -4266 196954
rect -4886 196634 -4266 196718
rect -4886 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 -4266 196634
rect -4886 160954 -4266 196398
rect -4886 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 -4266 160954
rect -4886 160634 -4266 160718
rect -4886 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 -4266 160634
rect -4886 124954 -4266 160398
rect -4886 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 -4266 124954
rect -4886 124634 -4266 124718
rect -4886 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 -4266 124634
rect -4886 88954 -4266 124398
rect -4886 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 -4266 88954
rect -4886 88634 -4266 88718
rect -4886 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 -4266 88634
rect -4886 52954 -4266 88398
rect -4886 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 -4266 52954
rect -4886 52634 -4266 52718
rect -4886 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 -4266 52634
rect -4886 16954 -4266 52398
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 -4266 16954
rect -4886 16634 -4266 16718
rect -4886 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 -4266 16634
rect -4886 -3226 -4266 16398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 696454 -3306 706202
rect -3926 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 -3306 696454
rect -3926 696134 -3306 696218
rect -3926 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 -3306 696134
rect -3926 660454 -3306 695898
rect -3926 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 -3306 660454
rect -3926 660134 -3306 660218
rect -3926 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 -3306 660134
rect -3926 624454 -3306 659898
rect -3926 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 -3306 624454
rect -3926 624134 -3306 624218
rect -3926 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 -3306 624134
rect -3926 588454 -3306 623898
rect -3926 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 -3306 588454
rect -3926 588134 -3306 588218
rect -3926 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 -3306 588134
rect -3926 552454 -3306 587898
rect -3926 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 -3306 552454
rect -3926 552134 -3306 552218
rect -3926 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 -3306 552134
rect -3926 516454 -3306 551898
rect -3926 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 -3306 516454
rect -3926 516134 -3306 516218
rect -3926 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 -3306 516134
rect -3926 480454 -3306 515898
rect -3926 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 -3306 480454
rect -3926 480134 -3306 480218
rect -3926 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 -3306 480134
rect -3926 444454 -3306 479898
rect -3926 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 -3306 444454
rect -3926 444134 -3306 444218
rect -3926 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 -3306 444134
rect -3926 408454 -3306 443898
rect -3926 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 -3306 408454
rect -3926 408134 -3306 408218
rect -3926 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 -3306 408134
rect -3926 372454 -3306 407898
rect -3926 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 -3306 372454
rect -3926 372134 -3306 372218
rect -3926 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 -3306 372134
rect -3926 336454 -3306 371898
rect -3926 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 -3306 336454
rect -3926 336134 -3306 336218
rect -3926 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 -3306 336134
rect -3926 300454 -3306 335898
rect -3926 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 -3306 300454
rect -3926 300134 -3306 300218
rect -3926 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 -3306 300134
rect -3926 264454 -3306 299898
rect -3926 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 -3306 264454
rect -3926 264134 -3306 264218
rect -3926 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 -3306 264134
rect -3926 228454 -3306 263898
rect -3926 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 -3306 228454
rect -3926 228134 -3306 228218
rect -3926 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 -3306 228134
rect -3926 192454 -3306 227898
rect -3926 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 -3306 192454
rect -3926 192134 -3306 192218
rect -3926 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 -3306 192134
rect -3926 156454 -3306 191898
rect -3926 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 -3306 156454
rect -3926 156134 -3306 156218
rect -3926 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 -3306 156134
rect -3926 120454 -3306 155898
rect -3926 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 -3306 120454
rect -3926 120134 -3306 120218
rect -3926 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 -3306 120134
rect -3926 84454 -3306 119898
rect -3926 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 -3306 84454
rect -3926 84134 -3306 84218
rect -3926 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 -3306 84134
rect -3926 48454 -3306 83898
rect -3926 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 -3306 48454
rect -3926 48134 -3306 48218
rect -3926 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 -3306 48134
rect -3926 12454 -3306 47898
rect -3926 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 -3306 12454
rect -3926 12134 -3306 12218
rect -3926 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 -3306 12134
rect -3926 -2266 -3306 11898
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691954 -2346 705242
rect -2966 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 -2346 691954
rect -2966 691634 -2346 691718
rect -2966 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 -2346 691634
rect -2966 655954 -2346 691398
rect -2966 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 -2346 655954
rect -2966 655634 -2346 655718
rect -2966 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 -2346 655634
rect -2966 619954 -2346 655398
rect -2966 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 -2346 619954
rect -2966 619634 -2346 619718
rect -2966 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 -2346 619634
rect -2966 583954 -2346 619398
rect -2966 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 -2346 583954
rect -2966 583634 -2346 583718
rect -2966 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 -2346 583634
rect -2966 547954 -2346 583398
rect -2966 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 -2346 547954
rect -2966 547634 -2346 547718
rect -2966 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 -2346 547634
rect -2966 511954 -2346 547398
rect -2966 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 -2346 511954
rect -2966 511634 -2346 511718
rect -2966 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 -2346 511634
rect -2966 475954 -2346 511398
rect -2966 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 -2346 475954
rect -2966 475634 -2346 475718
rect -2966 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 -2346 475634
rect -2966 439954 -2346 475398
rect -2966 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 -2346 439954
rect -2966 439634 -2346 439718
rect -2966 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 -2346 439634
rect -2966 403954 -2346 439398
rect -2966 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 -2346 403954
rect -2966 403634 -2346 403718
rect -2966 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 -2346 403634
rect -2966 367954 -2346 403398
rect -2966 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 -2346 367954
rect -2966 367634 -2346 367718
rect -2966 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 -2346 367634
rect -2966 331954 -2346 367398
rect -2966 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 -2346 331954
rect -2966 331634 -2346 331718
rect -2966 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 -2346 331634
rect -2966 295954 -2346 331398
rect -2966 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 -2346 295954
rect -2966 295634 -2346 295718
rect -2966 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 -2346 295634
rect -2966 259954 -2346 295398
rect -2966 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 -2346 259954
rect -2966 259634 -2346 259718
rect -2966 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 -2346 259634
rect -2966 223954 -2346 259398
rect -2966 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 -2346 223954
rect -2966 223634 -2346 223718
rect -2966 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 -2346 223634
rect -2966 187954 -2346 223398
rect -2966 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 -2346 187954
rect -2966 187634 -2346 187718
rect -2966 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 -2346 187634
rect -2966 151954 -2346 187398
rect -2966 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 -2346 151954
rect -2966 151634 -2346 151718
rect -2966 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 -2346 151634
rect -2966 115954 -2346 151398
rect -2966 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 -2346 115954
rect -2966 115634 -2346 115718
rect -2966 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 -2346 115634
rect -2966 79954 -2346 115398
rect -2966 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 -2346 79954
rect -2966 79634 -2346 79718
rect -2966 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 -2346 79634
rect -2966 43954 -2346 79398
rect -2966 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 -2346 43954
rect -2966 43634 -2346 43718
rect -2966 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 -2346 43634
rect -2966 7954 -2346 43398
rect -2966 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 -2346 7954
rect -2966 7634 -2346 7718
rect -2966 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 -2346 7634
rect -2966 -1306 -2346 7398
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 6294 705798 6914 711590
rect 6294 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 6914 705798
rect 6294 705478 6914 705562
rect 6294 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 6914 705478
rect 6294 691954 6914 705242
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1306 6914 7398
rect 6294 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 6914 -1306
rect 6294 -1626 6914 -1542
rect 6294 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 6914 -1626
rect 6294 -7654 6914 -1862
rect 10794 706758 11414 711590
rect 10794 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 11414 706758
rect 10794 706438 11414 706522
rect 10794 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 11414 706438
rect 10794 696454 11414 706202
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2266 11414 11898
rect 10794 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 11414 -2266
rect 10794 -2586 11414 -2502
rect 10794 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 11414 -2586
rect 10794 -7654 11414 -2822
rect 15294 707718 15914 711590
rect 15294 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 15914 707718
rect 15294 707398 15914 707482
rect 15294 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 15914 707398
rect 15294 700954 15914 707162
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3226 15914 16398
rect 15294 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 15914 -3226
rect 15294 -3546 15914 -3462
rect 15294 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 15914 -3546
rect 15294 -7654 15914 -3782
rect 19794 708678 20414 711590
rect 19794 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 20414 708678
rect 19794 708358 20414 708442
rect 19794 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 20414 708358
rect 19794 669454 20414 708122
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4186 20414 20898
rect 19794 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 20414 -4186
rect 19794 -4506 20414 -4422
rect 19794 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 20414 -4506
rect 19794 -7654 20414 -4742
rect 24294 709638 24914 711590
rect 24294 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 24914 709638
rect 24294 709318 24914 709402
rect 24294 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 24914 709318
rect 24294 673954 24914 709082
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 133954 24914 169398
rect 24294 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 24914 133954
rect 24294 133634 24914 133718
rect 24294 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 24914 133634
rect 24294 97954 24914 133398
rect 24294 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 24914 97954
rect 24294 97634 24914 97718
rect 24294 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 24914 97634
rect 24294 61954 24914 97398
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5146 24914 25398
rect 24294 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 24914 -5146
rect 24294 -5466 24914 -5382
rect 24294 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 24914 -5466
rect 24294 -7654 24914 -5702
rect 28794 710598 29414 711590
rect 28794 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 29414 710598
rect 28794 710278 29414 710362
rect 28794 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 29414 710278
rect 28794 678454 29414 710042
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 138454 29414 173898
rect 28794 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 29414 138454
rect 28794 138134 29414 138218
rect 28794 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 29414 138134
rect 28794 102454 29414 137898
rect 28794 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 29414 102454
rect 28794 102134 29414 102218
rect 28794 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 29414 102134
rect 28794 66454 29414 101898
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6106 29414 29898
rect 28794 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 29414 -6106
rect 28794 -6426 29414 -6342
rect 28794 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 29414 -6426
rect 28794 -7654 29414 -6662
rect 33294 711558 33914 711590
rect 33294 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 33914 711558
rect 33294 711238 33914 711322
rect 33294 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 33914 711238
rect 33294 682954 33914 711002
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 646954 33914 682398
rect 33294 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 33914 646954
rect 33294 646634 33914 646718
rect 33294 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 33914 646634
rect 33294 610954 33914 646398
rect 33294 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 33914 610954
rect 33294 610634 33914 610718
rect 33294 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 33914 610634
rect 33294 574954 33914 610398
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 33294 502954 33914 538398
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 33294 466954 33914 502398
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 33294 394954 33914 430398
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 142954 33914 178398
rect 33294 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 33914 142954
rect 33294 142634 33914 142718
rect 33294 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 33914 142634
rect 33294 106954 33914 142398
rect 33294 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 33914 106954
rect 33294 106634 33914 106718
rect 33294 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 33914 106634
rect 33294 70954 33914 106398
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7066 33914 34398
rect 33294 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 33914 -7066
rect 33294 -7386 33914 -7302
rect 33294 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 33914 -7386
rect 33294 -7654 33914 -7622
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 42294 705798 42914 711590
rect 42294 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 42914 705798
rect 42294 705478 42914 705562
rect 42294 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 42914 705478
rect 42294 691954 42914 705242
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 655954 42914 691398
rect 42294 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 42914 655954
rect 42294 655634 42914 655718
rect 42294 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 42914 655634
rect 42294 619954 42914 655398
rect 42294 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 42914 619954
rect 42294 619634 42914 619718
rect 42294 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 42914 619634
rect 42294 583954 42914 619398
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 511954 42914 547398
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 42294 475954 42914 511398
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42294 439954 42914 475398
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 46794 706758 47414 711590
rect 46794 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 47414 706758
rect 46794 706438 47414 706522
rect 46794 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 47414 706438
rect 46794 696454 47414 706202
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 660454 47414 695898
rect 46794 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 47414 660454
rect 46794 660134 47414 660218
rect 46794 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 47414 660134
rect 46794 624454 47414 659898
rect 46794 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 47414 624454
rect 46794 624134 47414 624218
rect 46794 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 47414 624134
rect 46794 588454 47414 623898
rect 46794 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 47414 588454
rect 46794 588134 47414 588218
rect 46794 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 47414 588134
rect 46794 552454 47414 587898
rect 46794 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 47414 552454
rect 46794 552134 47414 552218
rect 46794 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 47414 552134
rect 46794 516454 47414 551898
rect 46794 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 47414 516454
rect 46794 516134 47414 516218
rect 46794 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 47414 516134
rect 46794 480454 47414 515898
rect 46794 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 47414 480454
rect 46794 480134 47414 480218
rect 46794 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 47414 480134
rect 46794 444454 47414 479898
rect 46794 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 47414 444454
rect 46794 444134 47414 444218
rect 46794 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 47414 444134
rect 46794 408454 47414 443898
rect 46794 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 47414 408454
rect 46794 408134 47414 408218
rect 46794 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 47414 408134
rect 46794 372454 47414 407898
rect 46794 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 47414 372454
rect 46794 372134 47414 372218
rect 46794 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 47414 372134
rect 46794 336454 47414 371898
rect 46794 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 47414 336454
rect 46794 336134 47414 336218
rect 46794 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 47414 336134
rect 46794 300454 47414 335898
rect 46794 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 47414 300454
rect 46794 300134 47414 300218
rect 46794 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 47414 300134
rect 46794 264454 47414 299898
rect 46794 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 47414 264454
rect 46794 264134 47414 264218
rect 46794 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 47414 264134
rect 46794 248684 47414 263898
rect 51294 707718 51914 711590
rect 51294 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 51914 707718
rect 51294 707398 51914 707482
rect 51294 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 51914 707398
rect 51294 700954 51914 707162
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 664954 51914 700398
rect 51294 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 51914 664954
rect 51294 664634 51914 664718
rect 51294 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 51914 664634
rect 51294 628954 51914 664398
rect 51294 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 51914 628954
rect 51294 628634 51914 628718
rect 51294 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 51914 628634
rect 51294 592954 51914 628398
rect 51294 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 51914 592954
rect 51294 592634 51914 592718
rect 51294 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 51914 592634
rect 51294 556954 51914 592398
rect 51294 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 51914 556954
rect 51294 556634 51914 556718
rect 51294 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 51914 556634
rect 51294 520954 51914 556398
rect 51294 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 51914 520954
rect 51294 520634 51914 520718
rect 51294 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 51914 520634
rect 51294 484954 51914 520398
rect 51294 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 51914 484954
rect 51294 484634 51914 484718
rect 51294 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 51914 484634
rect 51294 448954 51914 484398
rect 51294 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 51914 448954
rect 51294 448634 51914 448718
rect 51294 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 51914 448634
rect 51294 412954 51914 448398
rect 51294 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 51914 412954
rect 51294 412634 51914 412718
rect 51294 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 51914 412634
rect 51294 376954 51914 412398
rect 51294 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 51914 376954
rect 51294 376634 51914 376718
rect 51294 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 51914 376634
rect 51294 340954 51914 376398
rect 51294 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 51914 340954
rect 51294 340634 51914 340718
rect 51294 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 51914 340634
rect 51294 304954 51914 340398
rect 51294 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 51914 304954
rect 51294 304634 51914 304718
rect 51294 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 51914 304634
rect 51294 268954 51914 304398
rect 51294 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 51914 268954
rect 51294 268634 51914 268718
rect 51294 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 51914 268634
rect 51294 248684 51914 268398
rect 55794 708678 56414 711590
rect 55794 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 56414 708678
rect 55794 708358 56414 708442
rect 55794 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 56414 708358
rect 55794 669454 56414 708122
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 248684 56414 272898
rect 60294 709638 60914 711590
rect 60294 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 60914 709638
rect 60294 709318 60914 709402
rect 60294 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 60914 709318
rect 60294 673954 60914 709082
rect 60294 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 60914 673954
rect 60294 673634 60914 673718
rect 60294 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 60914 673634
rect 60294 637954 60914 673398
rect 60294 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 60914 637954
rect 60294 637634 60914 637718
rect 60294 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 60914 637634
rect 60294 601954 60914 637398
rect 60294 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 60914 601954
rect 60294 601634 60914 601718
rect 60294 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 60914 601634
rect 60294 565954 60914 601398
rect 60294 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 60914 565954
rect 60294 565634 60914 565718
rect 60294 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 60914 565634
rect 60294 529954 60914 565398
rect 60294 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 60914 529954
rect 60294 529634 60914 529718
rect 60294 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 60914 529634
rect 60294 493954 60914 529398
rect 60294 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 60914 493954
rect 60294 493634 60914 493718
rect 60294 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 60914 493634
rect 60294 457954 60914 493398
rect 60294 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 60914 457954
rect 60294 457634 60914 457718
rect 60294 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 60914 457634
rect 60294 421954 60914 457398
rect 60294 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 60914 421954
rect 60294 421634 60914 421718
rect 60294 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 60914 421634
rect 60294 385954 60914 421398
rect 60294 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 60914 385954
rect 60294 385634 60914 385718
rect 60294 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 60914 385634
rect 60294 349954 60914 385398
rect 60294 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 60914 349954
rect 60294 349634 60914 349718
rect 60294 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 60914 349634
rect 60294 313954 60914 349398
rect 60294 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 60914 313954
rect 60294 313634 60914 313718
rect 60294 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 60914 313634
rect 60294 277954 60914 313398
rect 60294 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 60914 277954
rect 60294 277634 60914 277718
rect 60294 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 60914 277634
rect 60294 248684 60914 277398
rect 64794 710598 65414 711590
rect 64794 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 65414 710598
rect 64794 710278 65414 710362
rect 64794 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 65414 710278
rect 64794 678454 65414 710042
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 642454 65414 677898
rect 64794 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 65414 642454
rect 64794 642134 65414 642218
rect 64794 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 65414 642134
rect 64794 606454 65414 641898
rect 64794 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 65414 606454
rect 64794 606134 65414 606218
rect 64794 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 65414 606134
rect 64794 570454 65414 605898
rect 64794 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 65414 570454
rect 64794 570134 65414 570218
rect 64794 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 65414 570134
rect 64794 534454 65414 569898
rect 64794 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 65414 534454
rect 64794 534134 65414 534218
rect 64794 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 65414 534134
rect 64794 498454 65414 533898
rect 64794 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 65414 498454
rect 64794 498134 65414 498218
rect 64794 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 65414 498134
rect 64794 462454 65414 497898
rect 64794 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 65414 462454
rect 64794 462134 65414 462218
rect 64794 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 65414 462134
rect 64794 426454 65414 461898
rect 64794 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 65414 426454
rect 64794 426134 65414 426218
rect 64794 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 65414 426134
rect 64794 390454 65414 425898
rect 64794 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 65414 390454
rect 64794 390134 65414 390218
rect 64794 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 65414 390134
rect 64794 354454 65414 389898
rect 64794 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 65414 354454
rect 64794 354134 65414 354218
rect 64794 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 65414 354134
rect 64794 318454 65414 353898
rect 64794 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 65414 318454
rect 64794 318134 65414 318218
rect 64794 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 65414 318134
rect 64794 282454 65414 317898
rect 64794 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 65414 282454
rect 64794 282134 65414 282218
rect 64794 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 65414 282134
rect 64794 248684 65414 281898
rect 69294 711558 69914 711590
rect 69294 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 69914 711558
rect 69294 711238 69914 711322
rect 69294 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 69914 711238
rect 69294 682954 69914 711002
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 646954 69914 682398
rect 69294 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 69914 646954
rect 69294 646634 69914 646718
rect 69294 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 69914 646634
rect 69294 610954 69914 646398
rect 69294 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 69914 610954
rect 69294 610634 69914 610718
rect 69294 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 69914 610634
rect 69294 574954 69914 610398
rect 69294 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 69914 574954
rect 69294 574634 69914 574718
rect 69294 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 69914 574634
rect 69294 538954 69914 574398
rect 69294 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 69914 538954
rect 69294 538634 69914 538718
rect 69294 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 69914 538634
rect 69294 502954 69914 538398
rect 69294 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 69914 502954
rect 69294 502634 69914 502718
rect 69294 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 69914 502634
rect 69294 466954 69914 502398
rect 69294 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 69914 466954
rect 69294 466634 69914 466718
rect 69294 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 69914 466634
rect 69294 430954 69914 466398
rect 69294 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 69914 430954
rect 69294 430634 69914 430718
rect 69294 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 69914 430634
rect 69294 394954 69914 430398
rect 69294 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 69914 394954
rect 69294 394634 69914 394718
rect 69294 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 69914 394634
rect 69294 358954 69914 394398
rect 69294 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 69914 358954
rect 69294 358634 69914 358718
rect 69294 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 69914 358634
rect 69294 322954 69914 358398
rect 69294 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 69914 322954
rect 69294 322634 69914 322718
rect 69294 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 69914 322634
rect 69294 286954 69914 322398
rect 69294 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 69914 286954
rect 69294 286634 69914 286718
rect 69294 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 69914 286634
rect 69294 250954 69914 286398
rect 69294 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 69914 250954
rect 69294 250634 69914 250718
rect 69294 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 69914 250634
rect 69294 248684 69914 250398
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 248684 74414 254898
rect 78294 705798 78914 711590
rect 78294 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 78914 705798
rect 78294 705478 78914 705562
rect 78294 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 78914 705478
rect 78294 691954 78914 705242
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 655954 78914 691398
rect 78294 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 78914 655954
rect 78294 655634 78914 655718
rect 78294 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 78914 655634
rect 78294 619954 78914 655398
rect 78294 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 78914 619954
rect 78294 619634 78914 619718
rect 78294 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 78914 619634
rect 78294 583954 78914 619398
rect 78294 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 78914 583954
rect 78294 583634 78914 583718
rect 78294 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 78914 583634
rect 78294 547954 78914 583398
rect 78294 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 78914 547954
rect 78294 547634 78914 547718
rect 78294 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 78914 547634
rect 78294 511954 78914 547398
rect 78294 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 78914 511954
rect 78294 511634 78914 511718
rect 78294 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 78914 511634
rect 78294 475954 78914 511398
rect 78294 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 78914 475954
rect 78294 475634 78914 475718
rect 78294 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 78914 475634
rect 78294 439954 78914 475398
rect 78294 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 78914 439954
rect 78294 439634 78914 439718
rect 78294 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 78914 439634
rect 78294 403954 78914 439398
rect 78294 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 78914 403954
rect 78294 403634 78914 403718
rect 78294 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 78914 403634
rect 78294 367954 78914 403398
rect 78294 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 78914 367954
rect 78294 367634 78914 367718
rect 78294 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 78914 367634
rect 78294 331954 78914 367398
rect 78294 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 78914 331954
rect 78294 331634 78914 331718
rect 78294 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 78914 331634
rect 78294 295954 78914 331398
rect 78294 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 78914 295954
rect 78294 295634 78914 295718
rect 78294 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 78914 295634
rect 78294 259954 78914 295398
rect 78294 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 78914 259954
rect 78294 259634 78914 259718
rect 78294 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 78914 259634
rect 78294 248684 78914 259398
rect 82794 706758 83414 711590
rect 82794 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 83414 706758
rect 82794 706438 83414 706522
rect 82794 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 83414 706438
rect 82794 696454 83414 706202
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 660454 83414 695898
rect 82794 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 83414 660454
rect 82794 660134 83414 660218
rect 82794 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 83414 660134
rect 82794 624454 83414 659898
rect 82794 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 83414 624454
rect 82794 624134 83414 624218
rect 82794 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 83414 624134
rect 82794 588454 83414 623898
rect 82794 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 83414 588454
rect 82794 588134 83414 588218
rect 82794 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 83414 588134
rect 82794 552454 83414 587898
rect 82794 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 83414 552454
rect 82794 552134 83414 552218
rect 82794 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 83414 552134
rect 82794 516454 83414 551898
rect 82794 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 83414 516454
rect 82794 516134 83414 516218
rect 82794 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 83414 516134
rect 82794 480454 83414 515898
rect 82794 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 83414 480454
rect 82794 480134 83414 480218
rect 82794 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 83414 480134
rect 82794 444454 83414 479898
rect 82794 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 83414 444454
rect 82794 444134 83414 444218
rect 82794 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 83414 444134
rect 82794 408454 83414 443898
rect 82794 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 83414 408454
rect 82794 408134 83414 408218
rect 82794 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 83414 408134
rect 82794 372454 83414 407898
rect 82794 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 83414 372454
rect 82794 372134 83414 372218
rect 82794 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 83414 372134
rect 82794 336454 83414 371898
rect 82794 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 83414 336454
rect 82794 336134 83414 336218
rect 82794 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 83414 336134
rect 82794 300454 83414 335898
rect 82794 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 83414 300454
rect 82794 300134 83414 300218
rect 82794 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 83414 300134
rect 82794 264454 83414 299898
rect 82794 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 83414 264454
rect 82794 264134 83414 264218
rect 82794 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 83414 264134
rect 82794 248684 83414 263898
rect 87294 707718 87914 711590
rect 87294 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 87914 707718
rect 87294 707398 87914 707482
rect 87294 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 87914 707398
rect 87294 700954 87914 707162
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 664954 87914 700398
rect 87294 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 87914 664954
rect 87294 664634 87914 664718
rect 87294 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 87914 664634
rect 87294 628954 87914 664398
rect 87294 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 87914 628954
rect 87294 628634 87914 628718
rect 87294 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 87914 628634
rect 87294 592954 87914 628398
rect 87294 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 87914 592954
rect 87294 592634 87914 592718
rect 87294 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 87914 592634
rect 87294 556954 87914 592398
rect 87294 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 87914 556954
rect 87294 556634 87914 556718
rect 87294 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 87914 556634
rect 87294 520954 87914 556398
rect 87294 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 87914 520954
rect 87294 520634 87914 520718
rect 87294 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 87914 520634
rect 87294 484954 87914 520398
rect 87294 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 87914 484954
rect 87294 484634 87914 484718
rect 87294 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 87914 484634
rect 87294 448954 87914 484398
rect 87294 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 87914 448954
rect 87294 448634 87914 448718
rect 87294 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 87914 448634
rect 87294 412954 87914 448398
rect 87294 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 87914 412954
rect 87294 412634 87914 412718
rect 87294 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 87914 412634
rect 87294 376954 87914 412398
rect 87294 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 87914 376954
rect 87294 376634 87914 376718
rect 87294 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 87914 376634
rect 87294 340954 87914 376398
rect 87294 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 87914 340954
rect 87294 340634 87914 340718
rect 87294 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 87914 340634
rect 87294 304954 87914 340398
rect 87294 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 87914 304954
rect 87294 304634 87914 304718
rect 87294 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 87914 304634
rect 87294 268954 87914 304398
rect 87294 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 87914 268954
rect 87294 268634 87914 268718
rect 87294 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 87914 268634
rect 87294 248684 87914 268398
rect 91794 708678 92414 711590
rect 91794 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 92414 708678
rect 91794 708358 92414 708442
rect 91794 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 92414 708358
rect 91794 669454 92414 708122
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 248684 92414 272898
rect 96294 709638 96914 711590
rect 96294 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 96914 709638
rect 96294 709318 96914 709402
rect 96294 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 96914 709318
rect 96294 673954 96914 709082
rect 96294 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 96914 673954
rect 96294 673634 96914 673718
rect 96294 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 96914 673634
rect 96294 637954 96914 673398
rect 96294 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 96914 637954
rect 96294 637634 96914 637718
rect 96294 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 96914 637634
rect 96294 601954 96914 637398
rect 96294 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 96914 601954
rect 96294 601634 96914 601718
rect 96294 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 96914 601634
rect 96294 565954 96914 601398
rect 96294 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 96914 565954
rect 96294 565634 96914 565718
rect 96294 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 96914 565634
rect 96294 529954 96914 565398
rect 96294 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 96914 529954
rect 96294 529634 96914 529718
rect 96294 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 96914 529634
rect 96294 493954 96914 529398
rect 96294 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 96914 493954
rect 96294 493634 96914 493718
rect 96294 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 96914 493634
rect 96294 457954 96914 493398
rect 96294 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 96914 457954
rect 96294 457634 96914 457718
rect 96294 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 96914 457634
rect 96294 421954 96914 457398
rect 96294 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 96914 421954
rect 96294 421634 96914 421718
rect 96294 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 96914 421634
rect 96294 385954 96914 421398
rect 96294 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 96914 385954
rect 96294 385634 96914 385718
rect 96294 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 96914 385634
rect 96294 349954 96914 385398
rect 96294 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 96914 349954
rect 96294 349634 96914 349718
rect 96294 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 96914 349634
rect 96294 313954 96914 349398
rect 96294 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 96914 313954
rect 96294 313634 96914 313718
rect 96294 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 96914 313634
rect 96294 277954 96914 313398
rect 96294 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 96914 277954
rect 96294 277634 96914 277718
rect 96294 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 96914 277634
rect 96294 248684 96914 277398
rect 100794 710598 101414 711590
rect 100794 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 101414 710598
rect 100794 710278 101414 710362
rect 100794 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 101414 710278
rect 100794 678454 101414 710042
rect 100794 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 101414 678454
rect 100794 678134 101414 678218
rect 100794 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 101414 678134
rect 100794 642454 101414 677898
rect 100794 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 101414 642454
rect 100794 642134 101414 642218
rect 100794 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 101414 642134
rect 100794 606454 101414 641898
rect 100794 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 101414 606454
rect 100794 606134 101414 606218
rect 100794 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 101414 606134
rect 100794 570454 101414 605898
rect 100794 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 101414 570454
rect 100794 570134 101414 570218
rect 100794 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 101414 570134
rect 100794 534454 101414 569898
rect 100794 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 101414 534454
rect 100794 534134 101414 534218
rect 100794 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 101414 534134
rect 100794 498454 101414 533898
rect 100794 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 101414 498454
rect 100794 498134 101414 498218
rect 100794 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 101414 498134
rect 100794 462454 101414 497898
rect 100794 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 101414 462454
rect 100794 462134 101414 462218
rect 100794 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 101414 462134
rect 100794 426454 101414 461898
rect 100794 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 101414 426454
rect 100794 426134 101414 426218
rect 100794 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 101414 426134
rect 100794 390454 101414 425898
rect 100794 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 101414 390454
rect 100794 390134 101414 390218
rect 100794 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 101414 390134
rect 100794 354454 101414 389898
rect 100794 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 101414 354454
rect 100794 354134 101414 354218
rect 100794 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 101414 354134
rect 100794 318454 101414 353898
rect 100794 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 101414 318454
rect 100794 318134 101414 318218
rect 100794 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 101414 318134
rect 100794 282454 101414 317898
rect 100794 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 101414 282454
rect 100794 282134 101414 282218
rect 100794 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 101414 282134
rect 100794 248684 101414 281898
rect 105294 711558 105914 711590
rect 105294 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 105914 711558
rect 105294 711238 105914 711322
rect 105294 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 105914 711238
rect 105294 682954 105914 711002
rect 105294 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 105914 682954
rect 105294 682634 105914 682718
rect 105294 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 105914 682634
rect 105294 646954 105914 682398
rect 105294 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 105914 646954
rect 105294 646634 105914 646718
rect 105294 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 105914 646634
rect 105294 610954 105914 646398
rect 105294 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 105914 610954
rect 105294 610634 105914 610718
rect 105294 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 105914 610634
rect 105294 574954 105914 610398
rect 105294 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 105914 574954
rect 105294 574634 105914 574718
rect 105294 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 105914 574634
rect 105294 538954 105914 574398
rect 105294 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 105914 538954
rect 105294 538634 105914 538718
rect 105294 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 105914 538634
rect 105294 502954 105914 538398
rect 105294 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 105914 502954
rect 105294 502634 105914 502718
rect 105294 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 105914 502634
rect 105294 466954 105914 502398
rect 105294 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 105914 466954
rect 105294 466634 105914 466718
rect 105294 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 105914 466634
rect 105294 430954 105914 466398
rect 105294 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 105914 430954
rect 105294 430634 105914 430718
rect 105294 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 105914 430634
rect 105294 394954 105914 430398
rect 105294 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 105914 394954
rect 105294 394634 105914 394718
rect 105294 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 105914 394634
rect 105294 358954 105914 394398
rect 105294 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 105914 358954
rect 105294 358634 105914 358718
rect 105294 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 105914 358634
rect 105294 322954 105914 358398
rect 105294 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 105914 322954
rect 105294 322634 105914 322718
rect 105294 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 105914 322634
rect 105294 286954 105914 322398
rect 105294 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 105914 286954
rect 105294 286634 105914 286718
rect 105294 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 105914 286634
rect 105294 250954 105914 286398
rect 105294 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 105914 250954
rect 105294 250634 105914 250718
rect 105294 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 105914 250634
rect 105294 248684 105914 250398
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 248684 110414 254898
rect 114294 705798 114914 711590
rect 114294 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 114914 705798
rect 114294 705478 114914 705562
rect 114294 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 114914 705478
rect 114294 691954 114914 705242
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 655954 114914 691398
rect 114294 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 114914 655954
rect 114294 655634 114914 655718
rect 114294 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 114914 655634
rect 114294 619954 114914 655398
rect 114294 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 114914 619954
rect 114294 619634 114914 619718
rect 114294 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 114914 619634
rect 114294 583954 114914 619398
rect 114294 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 114914 583954
rect 114294 583634 114914 583718
rect 114294 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 114914 583634
rect 114294 547954 114914 583398
rect 114294 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 114914 547954
rect 114294 547634 114914 547718
rect 114294 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 114914 547634
rect 114294 511954 114914 547398
rect 114294 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 114914 511954
rect 114294 511634 114914 511718
rect 114294 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 114914 511634
rect 114294 475954 114914 511398
rect 114294 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 114914 475954
rect 114294 475634 114914 475718
rect 114294 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 114914 475634
rect 114294 439954 114914 475398
rect 114294 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 114914 439954
rect 114294 439634 114914 439718
rect 114294 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 114914 439634
rect 114294 403954 114914 439398
rect 114294 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 114914 403954
rect 114294 403634 114914 403718
rect 114294 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 114914 403634
rect 114294 367954 114914 403398
rect 114294 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 114914 367954
rect 114294 367634 114914 367718
rect 114294 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 114914 367634
rect 114294 331954 114914 367398
rect 114294 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 114914 331954
rect 114294 331634 114914 331718
rect 114294 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 114914 331634
rect 114294 295954 114914 331398
rect 114294 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 114914 295954
rect 114294 295634 114914 295718
rect 114294 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 114914 295634
rect 114294 259954 114914 295398
rect 114294 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 114914 259954
rect 114294 259634 114914 259718
rect 114294 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 114914 259634
rect 114294 248684 114914 259398
rect 118794 706758 119414 711590
rect 118794 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 119414 706758
rect 118794 706438 119414 706522
rect 118794 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 119414 706438
rect 118794 696454 119414 706202
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 660454 119414 695898
rect 118794 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 119414 660454
rect 118794 660134 119414 660218
rect 118794 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 119414 660134
rect 118794 624454 119414 659898
rect 118794 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 119414 624454
rect 118794 624134 119414 624218
rect 118794 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 119414 624134
rect 118794 588454 119414 623898
rect 118794 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 119414 588454
rect 118794 588134 119414 588218
rect 118794 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 119414 588134
rect 118794 552454 119414 587898
rect 118794 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 119414 552454
rect 118794 552134 119414 552218
rect 118794 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 119414 552134
rect 118794 516454 119414 551898
rect 118794 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 119414 516454
rect 118794 516134 119414 516218
rect 118794 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 119414 516134
rect 118794 480454 119414 515898
rect 118794 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 119414 480454
rect 118794 480134 119414 480218
rect 118794 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 119414 480134
rect 118794 444454 119414 479898
rect 118794 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 119414 444454
rect 118794 444134 119414 444218
rect 118794 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 119414 444134
rect 118794 408454 119414 443898
rect 118794 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 119414 408454
rect 118794 408134 119414 408218
rect 118794 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 119414 408134
rect 118794 372454 119414 407898
rect 118794 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 119414 372454
rect 118794 372134 119414 372218
rect 118794 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 119414 372134
rect 118794 336454 119414 371898
rect 118794 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 119414 336454
rect 118794 336134 119414 336218
rect 118794 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 119414 336134
rect 118794 300454 119414 335898
rect 118794 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 119414 300454
rect 118794 300134 119414 300218
rect 118794 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 119414 300134
rect 118794 264454 119414 299898
rect 118794 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 119414 264454
rect 118794 264134 119414 264218
rect 118794 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 119414 264134
rect 118794 248684 119414 263898
rect 123294 707718 123914 711590
rect 123294 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 123914 707718
rect 123294 707398 123914 707482
rect 123294 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 123914 707398
rect 123294 700954 123914 707162
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 664954 123914 700398
rect 123294 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 123914 664954
rect 123294 664634 123914 664718
rect 123294 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 123914 664634
rect 123294 628954 123914 664398
rect 123294 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 123914 628954
rect 123294 628634 123914 628718
rect 123294 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 123914 628634
rect 123294 592954 123914 628398
rect 123294 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 123914 592954
rect 123294 592634 123914 592718
rect 123294 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 123914 592634
rect 123294 556954 123914 592398
rect 123294 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 123914 556954
rect 123294 556634 123914 556718
rect 123294 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 123914 556634
rect 123294 520954 123914 556398
rect 123294 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 123914 520954
rect 123294 520634 123914 520718
rect 123294 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 123914 520634
rect 123294 484954 123914 520398
rect 123294 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 123914 484954
rect 123294 484634 123914 484718
rect 123294 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 123914 484634
rect 123294 448954 123914 484398
rect 123294 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 123914 448954
rect 123294 448634 123914 448718
rect 123294 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 123914 448634
rect 123294 412954 123914 448398
rect 123294 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 123914 412954
rect 123294 412634 123914 412718
rect 123294 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 123914 412634
rect 123294 376954 123914 412398
rect 123294 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 123914 376954
rect 123294 376634 123914 376718
rect 123294 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 123914 376634
rect 123294 340954 123914 376398
rect 123294 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 123914 340954
rect 123294 340634 123914 340718
rect 123294 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 123914 340634
rect 123294 304954 123914 340398
rect 123294 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 123914 304954
rect 123294 304634 123914 304718
rect 123294 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 123914 304634
rect 123294 268954 123914 304398
rect 123294 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 123914 268954
rect 123294 268634 123914 268718
rect 123294 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 123914 268634
rect 123294 248684 123914 268398
rect 127794 708678 128414 711590
rect 127794 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 128414 708678
rect 127794 708358 128414 708442
rect 127794 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 128414 708358
rect 127794 669454 128414 708122
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 248684 128414 272898
rect 132294 709638 132914 711590
rect 132294 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 132914 709638
rect 132294 709318 132914 709402
rect 132294 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 132914 709318
rect 132294 673954 132914 709082
rect 132294 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 132914 673954
rect 132294 673634 132914 673718
rect 132294 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 132914 673634
rect 132294 637954 132914 673398
rect 132294 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 132914 637954
rect 132294 637634 132914 637718
rect 132294 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 132914 637634
rect 132294 601954 132914 637398
rect 132294 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 132914 601954
rect 132294 601634 132914 601718
rect 132294 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 132914 601634
rect 132294 565954 132914 601398
rect 132294 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 132914 565954
rect 132294 565634 132914 565718
rect 132294 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 132914 565634
rect 132294 529954 132914 565398
rect 132294 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 132914 529954
rect 132294 529634 132914 529718
rect 132294 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 132914 529634
rect 132294 493954 132914 529398
rect 132294 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 132914 493954
rect 132294 493634 132914 493718
rect 132294 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 132914 493634
rect 132294 457954 132914 493398
rect 132294 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 132914 457954
rect 132294 457634 132914 457718
rect 132294 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 132914 457634
rect 132294 421954 132914 457398
rect 132294 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 132914 421954
rect 132294 421634 132914 421718
rect 132294 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 132914 421634
rect 132294 385954 132914 421398
rect 132294 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 132914 385954
rect 132294 385634 132914 385718
rect 132294 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 132914 385634
rect 132294 349954 132914 385398
rect 132294 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 132914 349954
rect 132294 349634 132914 349718
rect 132294 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 132914 349634
rect 132294 313954 132914 349398
rect 132294 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 132914 313954
rect 132294 313634 132914 313718
rect 132294 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 132914 313634
rect 132294 277954 132914 313398
rect 132294 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 132914 277954
rect 132294 277634 132914 277718
rect 132294 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 132914 277634
rect 132294 248684 132914 277398
rect 136794 710598 137414 711590
rect 136794 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 137414 710598
rect 136794 710278 137414 710362
rect 136794 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 137414 710278
rect 136794 678454 137414 710042
rect 136794 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 137414 678454
rect 136794 678134 137414 678218
rect 136794 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 137414 678134
rect 136794 642454 137414 677898
rect 136794 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 137414 642454
rect 136794 642134 137414 642218
rect 136794 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 137414 642134
rect 136794 606454 137414 641898
rect 136794 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 137414 606454
rect 136794 606134 137414 606218
rect 136794 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 137414 606134
rect 136794 570454 137414 605898
rect 136794 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 137414 570454
rect 136794 570134 137414 570218
rect 136794 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 137414 570134
rect 136794 534454 137414 569898
rect 136794 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 137414 534454
rect 136794 534134 137414 534218
rect 136794 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 137414 534134
rect 136794 498454 137414 533898
rect 136794 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 137414 498454
rect 136794 498134 137414 498218
rect 136794 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 137414 498134
rect 136794 462454 137414 497898
rect 136794 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 137414 462454
rect 136794 462134 137414 462218
rect 136794 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 137414 462134
rect 136794 426454 137414 461898
rect 136794 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 137414 426454
rect 136794 426134 137414 426218
rect 136794 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 137414 426134
rect 136794 390454 137414 425898
rect 136794 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 137414 390454
rect 136794 390134 137414 390218
rect 136794 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 137414 390134
rect 136794 354454 137414 389898
rect 136794 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 137414 354454
rect 136794 354134 137414 354218
rect 136794 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 137414 354134
rect 136794 318454 137414 353898
rect 136794 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 137414 318454
rect 136794 318134 137414 318218
rect 136794 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 137414 318134
rect 136794 282454 137414 317898
rect 136794 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 137414 282454
rect 136794 282134 137414 282218
rect 136794 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 137414 282134
rect 136794 248684 137414 281898
rect 141294 711558 141914 711590
rect 141294 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 141914 711558
rect 141294 711238 141914 711322
rect 141294 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 141914 711238
rect 141294 682954 141914 711002
rect 141294 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 141914 682954
rect 141294 682634 141914 682718
rect 141294 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 141914 682634
rect 141294 646954 141914 682398
rect 141294 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 141914 646954
rect 141294 646634 141914 646718
rect 141294 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 141914 646634
rect 141294 610954 141914 646398
rect 141294 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 141914 610954
rect 141294 610634 141914 610718
rect 141294 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 141914 610634
rect 141294 574954 141914 610398
rect 141294 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 141914 574954
rect 141294 574634 141914 574718
rect 141294 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 141914 574634
rect 141294 538954 141914 574398
rect 141294 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 141914 538954
rect 141294 538634 141914 538718
rect 141294 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 141914 538634
rect 141294 502954 141914 538398
rect 141294 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 141914 502954
rect 141294 502634 141914 502718
rect 141294 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 141914 502634
rect 141294 466954 141914 502398
rect 141294 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 141914 466954
rect 141294 466634 141914 466718
rect 141294 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 141914 466634
rect 141294 430954 141914 466398
rect 141294 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 141914 430954
rect 141294 430634 141914 430718
rect 141294 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 141914 430634
rect 141294 394954 141914 430398
rect 141294 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 141914 394954
rect 141294 394634 141914 394718
rect 141294 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 141914 394634
rect 141294 358954 141914 394398
rect 141294 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 141914 358954
rect 141294 358634 141914 358718
rect 141294 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 141914 358634
rect 141294 322954 141914 358398
rect 141294 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 141914 322954
rect 141294 322634 141914 322718
rect 141294 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 141914 322634
rect 141294 286954 141914 322398
rect 141294 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 141914 286954
rect 141294 286634 141914 286718
rect 141294 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 141914 286634
rect 141294 250954 141914 286398
rect 141294 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 141914 250954
rect 141294 250634 141914 250718
rect 141294 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 141914 250634
rect 141294 248684 141914 250398
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 248684 146414 254898
rect 150294 705798 150914 711590
rect 150294 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 150914 705798
rect 150294 705478 150914 705562
rect 150294 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 150914 705478
rect 150294 691954 150914 705242
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 655954 150914 691398
rect 150294 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 150914 655954
rect 150294 655634 150914 655718
rect 150294 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 150914 655634
rect 150294 619954 150914 655398
rect 150294 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 150914 619954
rect 150294 619634 150914 619718
rect 150294 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 150914 619634
rect 150294 583954 150914 619398
rect 150294 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 150914 583954
rect 150294 583634 150914 583718
rect 150294 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 150914 583634
rect 150294 547954 150914 583398
rect 150294 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 150914 547954
rect 150294 547634 150914 547718
rect 150294 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 150914 547634
rect 150294 511954 150914 547398
rect 150294 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 150914 511954
rect 150294 511634 150914 511718
rect 150294 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 150914 511634
rect 150294 475954 150914 511398
rect 150294 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 150914 475954
rect 150294 475634 150914 475718
rect 150294 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 150914 475634
rect 150294 439954 150914 475398
rect 150294 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 150914 439954
rect 150294 439634 150914 439718
rect 150294 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 150914 439634
rect 150294 403954 150914 439398
rect 150294 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 150914 403954
rect 150294 403634 150914 403718
rect 150294 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 150914 403634
rect 150294 367954 150914 403398
rect 150294 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 150914 367954
rect 150294 367634 150914 367718
rect 150294 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 150914 367634
rect 150294 331954 150914 367398
rect 150294 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 150914 331954
rect 150294 331634 150914 331718
rect 150294 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 150914 331634
rect 150294 295954 150914 331398
rect 150294 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 150914 295954
rect 150294 295634 150914 295718
rect 150294 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 150914 295634
rect 150294 259954 150914 295398
rect 150294 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 150914 259954
rect 150294 259634 150914 259718
rect 150294 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 150914 259634
rect 150294 248684 150914 259398
rect 154794 706758 155414 711590
rect 154794 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 155414 706758
rect 154794 706438 155414 706522
rect 154794 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 155414 706438
rect 154794 696454 155414 706202
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 660454 155414 695898
rect 154794 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 155414 660454
rect 154794 660134 155414 660218
rect 154794 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 155414 660134
rect 154794 624454 155414 659898
rect 154794 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 155414 624454
rect 154794 624134 155414 624218
rect 154794 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 155414 624134
rect 154794 588454 155414 623898
rect 154794 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 155414 588454
rect 154794 588134 155414 588218
rect 154794 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 155414 588134
rect 154794 552454 155414 587898
rect 154794 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 155414 552454
rect 154794 552134 155414 552218
rect 154794 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 155414 552134
rect 154794 516454 155414 551898
rect 154794 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 155414 516454
rect 154794 516134 155414 516218
rect 154794 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 155414 516134
rect 154794 480454 155414 515898
rect 154794 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 155414 480454
rect 154794 480134 155414 480218
rect 154794 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 155414 480134
rect 154794 444454 155414 479898
rect 154794 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 155414 444454
rect 154794 444134 155414 444218
rect 154794 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 155414 444134
rect 154794 408454 155414 443898
rect 154794 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 155414 408454
rect 154794 408134 155414 408218
rect 154794 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 155414 408134
rect 154794 372454 155414 407898
rect 154794 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 155414 372454
rect 154794 372134 155414 372218
rect 154794 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 155414 372134
rect 154794 336454 155414 371898
rect 154794 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 155414 336454
rect 154794 336134 155414 336218
rect 154794 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 155414 336134
rect 154794 300454 155414 335898
rect 154794 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 155414 300454
rect 154794 300134 155414 300218
rect 154794 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 155414 300134
rect 154794 264454 155414 299898
rect 154794 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 155414 264454
rect 154794 264134 155414 264218
rect 154794 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 155414 264134
rect 154794 248684 155414 263898
rect 159294 707718 159914 711590
rect 159294 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 159914 707718
rect 159294 707398 159914 707482
rect 159294 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 159914 707398
rect 159294 700954 159914 707162
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 664954 159914 700398
rect 159294 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 159914 664954
rect 159294 664634 159914 664718
rect 159294 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 159914 664634
rect 159294 628954 159914 664398
rect 159294 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 159914 628954
rect 159294 628634 159914 628718
rect 159294 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 159914 628634
rect 159294 592954 159914 628398
rect 159294 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 159914 592954
rect 159294 592634 159914 592718
rect 159294 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 159914 592634
rect 159294 556954 159914 592398
rect 159294 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 159914 556954
rect 159294 556634 159914 556718
rect 159294 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 159914 556634
rect 159294 520954 159914 556398
rect 159294 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 159914 520954
rect 159294 520634 159914 520718
rect 159294 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 159914 520634
rect 159294 484954 159914 520398
rect 159294 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 159914 484954
rect 159294 484634 159914 484718
rect 159294 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 159914 484634
rect 159294 448954 159914 484398
rect 159294 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 159914 448954
rect 159294 448634 159914 448718
rect 159294 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 159914 448634
rect 159294 412954 159914 448398
rect 159294 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 159914 412954
rect 159294 412634 159914 412718
rect 159294 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 159914 412634
rect 159294 376954 159914 412398
rect 159294 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 159914 376954
rect 159294 376634 159914 376718
rect 159294 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 159914 376634
rect 159294 340954 159914 376398
rect 159294 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 159914 340954
rect 159294 340634 159914 340718
rect 159294 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 159914 340634
rect 159294 304954 159914 340398
rect 159294 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 159914 304954
rect 159294 304634 159914 304718
rect 159294 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 159914 304634
rect 159294 268954 159914 304398
rect 159294 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 159914 268954
rect 159294 268634 159914 268718
rect 159294 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 159914 268634
rect 159294 248684 159914 268398
rect 163794 708678 164414 711590
rect 163794 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 164414 708678
rect 163794 708358 164414 708442
rect 163794 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 164414 708358
rect 163794 669454 164414 708122
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 248684 164414 272898
rect 168294 709638 168914 711590
rect 168294 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 168914 709638
rect 168294 709318 168914 709402
rect 168294 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 168914 709318
rect 168294 673954 168914 709082
rect 168294 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 168914 673954
rect 168294 673634 168914 673718
rect 168294 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 168914 673634
rect 168294 637954 168914 673398
rect 168294 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 168914 637954
rect 168294 637634 168914 637718
rect 168294 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 168914 637634
rect 168294 601954 168914 637398
rect 168294 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 168914 601954
rect 168294 601634 168914 601718
rect 168294 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 168914 601634
rect 168294 565954 168914 601398
rect 168294 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 168914 565954
rect 168294 565634 168914 565718
rect 168294 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 168914 565634
rect 168294 529954 168914 565398
rect 168294 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 168914 529954
rect 168294 529634 168914 529718
rect 168294 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 168914 529634
rect 168294 493954 168914 529398
rect 168294 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 168914 493954
rect 168294 493634 168914 493718
rect 168294 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 168914 493634
rect 168294 457954 168914 493398
rect 168294 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 168914 457954
rect 168294 457634 168914 457718
rect 168294 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 168914 457634
rect 168294 421954 168914 457398
rect 168294 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 168914 421954
rect 168294 421634 168914 421718
rect 168294 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 168914 421634
rect 168294 385954 168914 421398
rect 168294 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 168914 385954
rect 168294 385634 168914 385718
rect 168294 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 168914 385634
rect 168294 349954 168914 385398
rect 168294 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 168914 349954
rect 168294 349634 168914 349718
rect 168294 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 168914 349634
rect 168294 313954 168914 349398
rect 168294 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 168914 313954
rect 168294 313634 168914 313718
rect 168294 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 168914 313634
rect 168294 277954 168914 313398
rect 168294 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 168914 277954
rect 168294 277634 168914 277718
rect 168294 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 168914 277634
rect 168294 248684 168914 277398
rect 172794 710598 173414 711590
rect 172794 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 173414 710598
rect 172794 710278 173414 710362
rect 172794 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 173414 710278
rect 172794 678454 173414 710042
rect 172794 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 173414 678454
rect 172794 678134 173414 678218
rect 172794 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 173414 678134
rect 172794 642454 173414 677898
rect 172794 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 173414 642454
rect 172794 642134 173414 642218
rect 172794 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 173414 642134
rect 172794 606454 173414 641898
rect 172794 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 173414 606454
rect 172794 606134 173414 606218
rect 172794 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 173414 606134
rect 172794 570454 173414 605898
rect 172794 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 173414 570454
rect 172794 570134 173414 570218
rect 172794 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 173414 570134
rect 172794 534454 173414 569898
rect 172794 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 173414 534454
rect 172794 534134 173414 534218
rect 172794 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 173414 534134
rect 172794 498454 173414 533898
rect 172794 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 173414 498454
rect 172794 498134 173414 498218
rect 172794 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 173414 498134
rect 172794 462454 173414 497898
rect 172794 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 173414 462454
rect 172794 462134 173414 462218
rect 172794 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 173414 462134
rect 172794 426454 173414 461898
rect 172794 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 173414 426454
rect 172794 426134 173414 426218
rect 172794 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 173414 426134
rect 172794 390454 173414 425898
rect 172794 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 173414 390454
rect 172794 390134 173414 390218
rect 172794 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 173414 390134
rect 172794 354454 173414 389898
rect 172794 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 173414 354454
rect 172794 354134 173414 354218
rect 172794 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 173414 354134
rect 172794 318454 173414 353898
rect 172794 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 173414 318454
rect 172794 318134 173414 318218
rect 172794 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 173414 318134
rect 172794 282454 173414 317898
rect 172794 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 173414 282454
rect 172794 282134 173414 282218
rect 172794 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 173414 282134
rect 172794 248684 173414 281898
rect 177294 711558 177914 711590
rect 177294 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 177914 711558
rect 177294 711238 177914 711322
rect 177294 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 177914 711238
rect 177294 682954 177914 711002
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 177294 646954 177914 682398
rect 177294 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 177914 646954
rect 177294 646634 177914 646718
rect 177294 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 177914 646634
rect 177294 610954 177914 646398
rect 177294 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 177914 610954
rect 177294 610634 177914 610718
rect 177294 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 177914 610634
rect 177294 574954 177914 610398
rect 177294 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 177914 574954
rect 177294 574634 177914 574718
rect 177294 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 177914 574634
rect 177294 538954 177914 574398
rect 177294 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 177914 538954
rect 177294 538634 177914 538718
rect 177294 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 177914 538634
rect 177294 502954 177914 538398
rect 177294 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 177914 502954
rect 177294 502634 177914 502718
rect 177294 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 177914 502634
rect 177294 466954 177914 502398
rect 177294 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 177914 466954
rect 177294 466634 177914 466718
rect 177294 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 177914 466634
rect 177294 430954 177914 466398
rect 177294 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 177914 430954
rect 177294 430634 177914 430718
rect 177294 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 177914 430634
rect 177294 394954 177914 430398
rect 177294 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 177914 394954
rect 177294 394634 177914 394718
rect 177294 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 177914 394634
rect 177294 358954 177914 394398
rect 177294 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 177914 358954
rect 177294 358634 177914 358718
rect 177294 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 177914 358634
rect 177294 322954 177914 358398
rect 177294 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 177914 322954
rect 177294 322634 177914 322718
rect 177294 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 177914 322634
rect 177294 286954 177914 322398
rect 177294 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 177914 286954
rect 177294 286634 177914 286718
rect 177294 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 177914 286634
rect 177294 250954 177914 286398
rect 177294 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 177914 250954
rect 177294 250634 177914 250718
rect 177294 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 177914 250634
rect 177294 248684 177914 250398
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 248684 182414 254898
rect 186294 705798 186914 711590
rect 186294 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 186914 705798
rect 186294 705478 186914 705562
rect 186294 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 186914 705478
rect 186294 691954 186914 705242
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 655954 186914 691398
rect 186294 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 186914 655954
rect 186294 655634 186914 655718
rect 186294 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 186914 655634
rect 186294 619954 186914 655398
rect 186294 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 186914 619954
rect 186294 619634 186914 619718
rect 186294 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 186914 619634
rect 186294 583954 186914 619398
rect 186294 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 186914 583954
rect 186294 583634 186914 583718
rect 186294 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 186914 583634
rect 186294 547954 186914 583398
rect 186294 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 186914 547954
rect 186294 547634 186914 547718
rect 186294 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 186914 547634
rect 186294 511954 186914 547398
rect 186294 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 186914 511954
rect 186294 511634 186914 511718
rect 186294 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 186914 511634
rect 186294 475954 186914 511398
rect 186294 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 186914 475954
rect 186294 475634 186914 475718
rect 186294 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 186914 475634
rect 186294 439954 186914 475398
rect 186294 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 186914 439954
rect 186294 439634 186914 439718
rect 186294 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 186914 439634
rect 186294 403954 186914 439398
rect 186294 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 186914 403954
rect 186294 403634 186914 403718
rect 186294 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 186914 403634
rect 186294 367954 186914 403398
rect 186294 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 186914 367954
rect 186294 367634 186914 367718
rect 186294 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 186914 367634
rect 186294 331954 186914 367398
rect 186294 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 186914 331954
rect 186294 331634 186914 331718
rect 186294 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 186914 331634
rect 186294 295954 186914 331398
rect 186294 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 186914 295954
rect 186294 295634 186914 295718
rect 186294 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 186914 295634
rect 186294 259954 186914 295398
rect 186294 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 186914 259954
rect 186294 259634 186914 259718
rect 186294 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 186914 259634
rect 186294 248684 186914 259398
rect 190794 706758 191414 711590
rect 190794 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 191414 706758
rect 190794 706438 191414 706522
rect 190794 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 191414 706438
rect 190794 696454 191414 706202
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 660454 191414 695898
rect 190794 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 191414 660454
rect 190794 660134 191414 660218
rect 190794 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 191414 660134
rect 190794 624454 191414 659898
rect 190794 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 191414 624454
rect 190794 624134 191414 624218
rect 190794 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 191414 624134
rect 190794 588454 191414 623898
rect 190794 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 191414 588454
rect 190794 588134 191414 588218
rect 190794 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 191414 588134
rect 190794 552454 191414 587898
rect 190794 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 191414 552454
rect 190794 552134 191414 552218
rect 190794 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 191414 552134
rect 190794 516454 191414 551898
rect 190794 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 191414 516454
rect 190794 516134 191414 516218
rect 190794 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 191414 516134
rect 190794 480454 191414 515898
rect 190794 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 191414 480454
rect 190794 480134 191414 480218
rect 190794 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 191414 480134
rect 190794 444454 191414 479898
rect 190794 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 191414 444454
rect 190794 444134 191414 444218
rect 190794 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 191414 444134
rect 190794 408454 191414 443898
rect 190794 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 191414 408454
rect 190794 408134 191414 408218
rect 190794 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 191414 408134
rect 190794 372454 191414 407898
rect 190794 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 191414 372454
rect 190794 372134 191414 372218
rect 190794 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 191414 372134
rect 190794 336454 191414 371898
rect 190794 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 191414 336454
rect 190794 336134 191414 336218
rect 190794 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 191414 336134
rect 190794 300454 191414 335898
rect 190794 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 191414 300454
rect 190794 300134 191414 300218
rect 190794 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 191414 300134
rect 190794 264454 191414 299898
rect 190794 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 191414 264454
rect 190794 264134 191414 264218
rect 190794 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 191414 264134
rect 190794 248684 191414 263898
rect 195294 707718 195914 711590
rect 195294 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 195914 707718
rect 195294 707398 195914 707482
rect 195294 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 195914 707398
rect 195294 700954 195914 707162
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 664954 195914 700398
rect 195294 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 195914 664954
rect 195294 664634 195914 664718
rect 195294 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 195914 664634
rect 195294 628954 195914 664398
rect 195294 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 195914 628954
rect 195294 628634 195914 628718
rect 195294 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 195914 628634
rect 195294 592954 195914 628398
rect 195294 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 195914 592954
rect 195294 592634 195914 592718
rect 195294 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 195914 592634
rect 195294 556954 195914 592398
rect 195294 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 195914 556954
rect 195294 556634 195914 556718
rect 195294 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 195914 556634
rect 195294 520954 195914 556398
rect 195294 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 195914 520954
rect 195294 520634 195914 520718
rect 195294 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 195914 520634
rect 195294 484954 195914 520398
rect 195294 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 195914 484954
rect 195294 484634 195914 484718
rect 195294 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 195914 484634
rect 195294 448954 195914 484398
rect 195294 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 195914 448954
rect 195294 448634 195914 448718
rect 195294 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 195914 448634
rect 195294 412954 195914 448398
rect 195294 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 195914 412954
rect 195294 412634 195914 412718
rect 195294 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 195914 412634
rect 195294 376954 195914 412398
rect 195294 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 195914 376954
rect 195294 376634 195914 376718
rect 195294 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 195914 376634
rect 195294 340954 195914 376398
rect 195294 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 195914 340954
rect 195294 340634 195914 340718
rect 195294 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 195914 340634
rect 195294 304954 195914 340398
rect 195294 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 195914 304954
rect 195294 304634 195914 304718
rect 195294 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 195914 304634
rect 195294 268954 195914 304398
rect 195294 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 195914 268954
rect 195294 268634 195914 268718
rect 195294 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 195914 268634
rect 195294 248684 195914 268398
rect 199794 708678 200414 711590
rect 199794 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 200414 708678
rect 199794 708358 200414 708442
rect 199794 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 200414 708358
rect 199794 669454 200414 708122
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 248684 200414 272898
rect 204294 709638 204914 711590
rect 204294 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 204914 709638
rect 204294 709318 204914 709402
rect 204294 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 204914 709318
rect 204294 673954 204914 709082
rect 204294 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 204914 673954
rect 204294 673634 204914 673718
rect 204294 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 204914 673634
rect 204294 637954 204914 673398
rect 204294 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 204914 637954
rect 204294 637634 204914 637718
rect 204294 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 204914 637634
rect 204294 601954 204914 637398
rect 204294 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 204914 601954
rect 204294 601634 204914 601718
rect 204294 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 204914 601634
rect 204294 565954 204914 601398
rect 204294 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 204914 565954
rect 204294 565634 204914 565718
rect 204294 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 204914 565634
rect 204294 529954 204914 565398
rect 204294 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 204914 529954
rect 204294 529634 204914 529718
rect 204294 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 204914 529634
rect 204294 493954 204914 529398
rect 204294 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 204914 493954
rect 204294 493634 204914 493718
rect 204294 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 204914 493634
rect 204294 457954 204914 493398
rect 204294 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 204914 457954
rect 204294 457634 204914 457718
rect 204294 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 204914 457634
rect 204294 421954 204914 457398
rect 204294 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 204914 421954
rect 204294 421634 204914 421718
rect 204294 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 204914 421634
rect 204294 385954 204914 421398
rect 204294 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 204914 385954
rect 204294 385634 204914 385718
rect 204294 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 204914 385634
rect 204294 349954 204914 385398
rect 204294 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 204914 349954
rect 204294 349634 204914 349718
rect 204294 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 204914 349634
rect 204294 313954 204914 349398
rect 204294 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 204914 313954
rect 204294 313634 204914 313718
rect 204294 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 204914 313634
rect 204294 277954 204914 313398
rect 204294 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 204914 277954
rect 204294 277634 204914 277718
rect 204294 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 204914 277634
rect 204294 248684 204914 277398
rect 208794 710598 209414 711590
rect 208794 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 209414 710598
rect 208794 710278 209414 710362
rect 208794 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 209414 710278
rect 208794 678454 209414 710042
rect 208794 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 209414 678454
rect 208794 678134 209414 678218
rect 208794 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 209414 678134
rect 208794 642454 209414 677898
rect 208794 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 209414 642454
rect 208794 642134 209414 642218
rect 208794 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 209414 642134
rect 208794 606454 209414 641898
rect 208794 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 209414 606454
rect 208794 606134 209414 606218
rect 208794 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 209414 606134
rect 208794 570454 209414 605898
rect 208794 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 209414 570454
rect 208794 570134 209414 570218
rect 208794 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 209414 570134
rect 208794 534454 209414 569898
rect 208794 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 209414 534454
rect 208794 534134 209414 534218
rect 208794 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 209414 534134
rect 208794 498454 209414 533898
rect 208794 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 209414 498454
rect 208794 498134 209414 498218
rect 208794 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 209414 498134
rect 208794 462454 209414 497898
rect 208794 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 209414 462454
rect 208794 462134 209414 462218
rect 208794 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 209414 462134
rect 208794 426454 209414 461898
rect 208794 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 209414 426454
rect 208794 426134 209414 426218
rect 208794 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 209414 426134
rect 208794 390454 209414 425898
rect 208794 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 209414 390454
rect 208794 390134 209414 390218
rect 208794 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 209414 390134
rect 208794 354454 209414 389898
rect 208794 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 209414 354454
rect 208794 354134 209414 354218
rect 208794 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 209414 354134
rect 208794 318454 209414 353898
rect 208794 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 209414 318454
rect 208794 318134 209414 318218
rect 208794 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 209414 318134
rect 208794 282454 209414 317898
rect 208794 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 209414 282454
rect 208794 282134 209414 282218
rect 208794 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 209414 282134
rect 208794 248684 209414 281898
rect 213294 711558 213914 711590
rect 213294 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 213914 711558
rect 213294 711238 213914 711322
rect 213294 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 213914 711238
rect 213294 682954 213914 711002
rect 213294 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 213914 682954
rect 213294 682634 213914 682718
rect 213294 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 213914 682634
rect 213294 646954 213914 682398
rect 213294 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 213914 646954
rect 213294 646634 213914 646718
rect 213294 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 213914 646634
rect 213294 610954 213914 646398
rect 213294 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 213914 610954
rect 213294 610634 213914 610718
rect 213294 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 213914 610634
rect 213294 574954 213914 610398
rect 213294 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 213914 574954
rect 213294 574634 213914 574718
rect 213294 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 213914 574634
rect 213294 538954 213914 574398
rect 213294 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 213914 538954
rect 213294 538634 213914 538718
rect 213294 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 213914 538634
rect 213294 502954 213914 538398
rect 213294 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 213914 502954
rect 213294 502634 213914 502718
rect 213294 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 213914 502634
rect 213294 466954 213914 502398
rect 213294 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 213914 466954
rect 213294 466634 213914 466718
rect 213294 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 213914 466634
rect 213294 430954 213914 466398
rect 213294 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 213914 430954
rect 213294 430634 213914 430718
rect 213294 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 213914 430634
rect 213294 394954 213914 430398
rect 213294 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 213914 394954
rect 213294 394634 213914 394718
rect 213294 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 213914 394634
rect 213294 358954 213914 394398
rect 213294 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 213914 358954
rect 213294 358634 213914 358718
rect 213294 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 213914 358634
rect 213294 322954 213914 358398
rect 213294 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 213914 322954
rect 213294 322634 213914 322718
rect 213294 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 213914 322634
rect 213294 286954 213914 322398
rect 213294 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 213914 286954
rect 213294 286634 213914 286718
rect 213294 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 213914 286634
rect 213294 250954 213914 286398
rect 213294 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 213914 250954
rect 213294 250634 213914 250718
rect 213294 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 213914 250634
rect 213294 248684 213914 250398
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 248684 218414 254898
rect 222294 705798 222914 711590
rect 222294 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 222914 705798
rect 222294 705478 222914 705562
rect 222294 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 222914 705478
rect 222294 691954 222914 705242
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 655954 222914 691398
rect 222294 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 222914 655954
rect 222294 655634 222914 655718
rect 222294 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 222914 655634
rect 222294 619954 222914 655398
rect 222294 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 222914 619954
rect 222294 619634 222914 619718
rect 222294 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 222914 619634
rect 222294 583954 222914 619398
rect 222294 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 222914 583954
rect 222294 583634 222914 583718
rect 222294 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 222914 583634
rect 222294 547954 222914 583398
rect 222294 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 222914 547954
rect 222294 547634 222914 547718
rect 222294 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 222914 547634
rect 222294 511954 222914 547398
rect 222294 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 222914 511954
rect 222294 511634 222914 511718
rect 222294 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 222914 511634
rect 222294 475954 222914 511398
rect 222294 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 222914 475954
rect 222294 475634 222914 475718
rect 222294 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 222914 475634
rect 222294 439954 222914 475398
rect 222294 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 222914 439954
rect 222294 439634 222914 439718
rect 222294 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 222914 439634
rect 222294 403954 222914 439398
rect 222294 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 222914 403954
rect 222294 403634 222914 403718
rect 222294 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 222914 403634
rect 222294 367954 222914 403398
rect 222294 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 222914 367954
rect 222294 367634 222914 367718
rect 222294 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 222914 367634
rect 222294 331954 222914 367398
rect 222294 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 222914 331954
rect 222294 331634 222914 331718
rect 222294 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 222914 331634
rect 222294 295954 222914 331398
rect 222294 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 222914 295954
rect 222294 295634 222914 295718
rect 222294 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 222914 295634
rect 222294 259954 222914 295398
rect 222294 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 222914 259954
rect 222294 259634 222914 259718
rect 222294 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 222914 259634
rect 222294 248684 222914 259398
rect 226794 706758 227414 711590
rect 226794 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 227414 706758
rect 226794 706438 227414 706522
rect 226794 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 227414 706438
rect 226794 696454 227414 706202
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 660454 227414 695898
rect 226794 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 227414 660454
rect 226794 660134 227414 660218
rect 226794 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 227414 660134
rect 226794 624454 227414 659898
rect 226794 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 227414 624454
rect 226794 624134 227414 624218
rect 226794 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 227414 624134
rect 226794 588454 227414 623898
rect 226794 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 227414 588454
rect 226794 588134 227414 588218
rect 226794 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 227414 588134
rect 226794 552454 227414 587898
rect 226794 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 227414 552454
rect 226794 552134 227414 552218
rect 226794 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 227414 552134
rect 226794 516454 227414 551898
rect 226794 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 227414 516454
rect 226794 516134 227414 516218
rect 226794 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 227414 516134
rect 226794 480454 227414 515898
rect 226794 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 227414 480454
rect 226794 480134 227414 480218
rect 226794 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 227414 480134
rect 226794 444454 227414 479898
rect 226794 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 227414 444454
rect 226794 444134 227414 444218
rect 226794 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 227414 444134
rect 226794 408454 227414 443898
rect 226794 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 227414 408454
rect 226794 408134 227414 408218
rect 226794 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 227414 408134
rect 226794 372454 227414 407898
rect 226794 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 227414 372454
rect 226794 372134 227414 372218
rect 226794 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 227414 372134
rect 226794 336454 227414 371898
rect 226794 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 227414 336454
rect 226794 336134 227414 336218
rect 226794 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 227414 336134
rect 226794 300454 227414 335898
rect 226794 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 227414 300454
rect 226794 300134 227414 300218
rect 226794 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 227414 300134
rect 226794 264454 227414 299898
rect 226794 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 227414 264454
rect 226794 264134 227414 264218
rect 226794 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 227414 264134
rect 226794 248684 227414 263898
rect 231294 707718 231914 711590
rect 231294 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 231914 707718
rect 231294 707398 231914 707482
rect 231294 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 231914 707398
rect 231294 700954 231914 707162
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 664954 231914 700398
rect 231294 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 231914 664954
rect 231294 664634 231914 664718
rect 231294 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 231914 664634
rect 231294 628954 231914 664398
rect 231294 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 231914 628954
rect 231294 628634 231914 628718
rect 231294 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 231914 628634
rect 231294 592954 231914 628398
rect 231294 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 231914 592954
rect 231294 592634 231914 592718
rect 231294 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 231914 592634
rect 231294 556954 231914 592398
rect 231294 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 231914 556954
rect 231294 556634 231914 556718
rect 231294 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 231914 556634
rect 231294 520954 231914 556398
rect 231294 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 231914 520954
rect 231294 520634 231914 520718
rect 231294 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 231914 520634
rect 231294 484954 231914 520398
rect 231294 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 231914 484954
rect 231294 484634 231914 484718
rect 231294 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 231914 484634
rect 231294 448954 231914 484398
rect 231294 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 231914 448954
rect 231294 448634 231914 448718
rect 231294 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 231914 448634
rect 231294 412954 231914 448398
rect 231294 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 231914 412954
rect 231294 412634 231914 412718
rect 231294 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 231914 412634
rect 231294 376954 231914 412398
rect 231294 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 231914 376954
rect 231294 376634 231914 376718
rect 231294 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 231914 376634
rect 231294 340954 231914 376398
rect 231294 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 231914 340954
rect 231294 340634 231914 340718
rect 231294 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 231914 340634
rect 231294 304954 231914 340398
rect 231294 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 231914 304954
rect 231294 304634 231914 304718
rect 231294 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 231914 304634
rect 231294 268954 231914 304398
rect 231294 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 231914 268954
rect 231294 268634 231914 268718
rect 231294 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 231914 268634
rect 231294 248684 231914 268398
rect 235794 708678 236414 711590
rect 235794 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 236414 708678
rect 235794 708358 236414 708442
rect 235794 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 236414 708358
rect 235794 669454 236414 708122
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 248684 236414 272898
rect 240294 709638 240914 711590
rect 240294 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 240914 709638
rect 240294 709318 240914 709402
rect 240294 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 240914 709318
rect 240294 673954 240914 709082
rect 240294 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 240914 673954
rect 240294 673634 240914 673718
rect 240294 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 240914 673634
rect 240294 637954 240914 673398
rect 240294 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 240914 637954
rect 240294 637634 240914 637718
rect 240294 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 240914 637634
rect 240294 601954 240914 637398
rect 240294 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 240914 601954
rect 240294 601634 240914 601718
rect 240294 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 240914 601634
rect 240294 565954 240914 601398
rect 240294 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 240914 565954
rect 240294 565634 240914 565718
rect 240294 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 240914 565634
rect 240294 529954 240914 565398
rect 240294 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 240914 529954
rect 240294 529634 240914 529718
rect 240294 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 240914 529634
rect 240294 493954 240914 529398
rect 240294 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 240914 493954
rect 240294 493634 240914 493718
rect 240294 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 240914 493634
rect 240294 457954 240914 493398
rect 240294 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 240914 457954
rect 240294 457634 240914 457718
rect 240294 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 240914 457634
rect 240294 421954 240914 457398
rect 240294 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 240914 421954
rect 240294 421634 240914 421718
rect 240294 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 240914 421634
rect 240294 385954 240914 421398
rect 240294 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 240914 385954
rect 240294 385634 240914 385718
rect 240294 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 240914 385634
rect 240294 349954 240914 385398
rect 240294 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 240914 349954
rect 240294 349634 240914 349718
rect 240294 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 240914 349634
rect 240294 313954 240914 349398
rect 240294 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 240914 313954
rect 240294 313634 240914 313718
rect 240294 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 240914 313634
rect 240294 277954 240914 313398
rect 240294 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 240914 277954
rect 240294 277634 240914 277718
rect 240294 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 240914 277634
rect 240294 248684 240914 277398
rect 244794 710598 245414 711590
rect 244794 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 245414 710598
rect 244794 710278 245414 710362
rect 244794 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 245414 710278
rect 244794 678454 245414 710042
rect 244794 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 245414 678454
rect 244794 678134 245414 678218
rect 244794 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 245414 678134
rect 244794 642454 245414 677898
rect 244794 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 245414 642454
rect 244794 642134 245414 642218
rect 244794 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 245414 642134
rect 244794 606454 245414 641898
rect 244794 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 245414 606454
rect 244794 606134 245414 606218
rect 244794 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 245414 606134
rect 244794 570454 245414 605898
rect 244794 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 245414 570454
rect 244794 570134 245414 570218
rect 244794 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 245414 570134
rect 244794 534454 245414 569898
rect 244794 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 245414 534454
rect 244794 534134 245414 534218
rect 244794 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 245414 534134
rect 244794 498454 245414 533898
rect 244794 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 245414 498454
rect 244794 498134 245414 498218
rect 244794 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 245414 498134
rect 244794 462454 245414 497898
rect 244794 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 245414 462454
rect 244794 462134 245414 462218
rect 244794 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 245414 462134
rect 244794 426454 245414 461898
rect 244794 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 245414 426454
rect 244794 426134 245414 426218
rect 244794 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 245414 426134
rect 244794 390454 245414 425898
rect 244794 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 245414 390454
rect 244794 390134 245414 390218
rect 244794 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 245414 390134
rect 244794 354454 245414 389898
rect 244794 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 245414 354454
rect 244794 354134 245414 354218
rect 244794 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 245414 354134
rect 244794 318454 245414 353898
rect 244794 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 245414 318454
rect 244794 318134 245414 318218
rect 244794 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 245414 318134
rect 244794 282454 245414 317898
rect 244794 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 245414 282454
rect 244794 282134 245414 282218
rect 244794 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 245414 282134
rect 244794 248684 245414 281898
rect 249294 711558 249914 711590
rect 249294 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 249914 711558
rect 249294 711238 249914 711322
rect 249294 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 249914 711238
rect 249294 682954 249914 711002
rect 249294 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 249914 682954
rect 249294 682634 249914 682718
rect 249294 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 249914 682634
rect 249294 646954 249914 682398
rect 249294 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 249914 646954
rect 249294 646634 249914 646718
rect 249294 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 249914 646634
rect 249294 610954 249914 646398
rect 249294 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 249914 610954
rect 249294 610634 249914 610718
rect 249294 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 249914 610634
rect 249294 574954 249914 610398
rect 249294 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 249914 574954
rect 249294 574634 249914 574718
rect 249294 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 249914 574634
rect 249294 538954 249914 574398
rect 249294 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 249914 538954
rect 249294 538634 249914 538718
rect 249294 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 249914 538634
rect 249294 502954 249914 538398
rect 249294 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 249914 502954
rect 249294 502634 249914 502718
rect 249294 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 249914 502634
rect 249294 466954 249914 502398
rect 249294 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 249914 466954
rect 249294 466634 249914 466718
rect 249294 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 249914 466634
rect 249294 430954 249914 466398
rect 249294 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 249914 430954
rect 249294 430634 249914 430718
rect 249294 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 249914 430634
rect 249294 394954 249914 430398
rect 249294 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 249914 394954
rect 249294 394634 249914 394718
rect 249294 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 249914 394634
rect 249294 358954 249914 394398
rect 249294 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 249914 358954
rect 249294 358634 249914 358718
rect 249294 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 249914 358634
rect 249294 322954 249914 358398
rect 249294 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 249914 322954
rect 249294 322634 249914 322718
rect 249294 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 249914 322634
rect 249294 286954 249914 322398
rect 249294 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 249914 286954
rect 249294 286634 249914 286718
rect 249294 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 249914 286634
rect 249294 250954 249914 286398
rect 249294 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 249914 250954
rect 249294 250634 249914 250718
rect 249294 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 249914 250634
rect 249294 248684 249914 250398
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 248684 254414 254898
rect 258294 705798 258914 711590
rect 258294 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 258914 705798
rect 258294 705478 258914 705562
rect 258294 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 258914 705478
rect 258294 691954 258914 705242
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 655954 258914 691398
rect 258294 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 258914 655954
rect 258294 655634 258914 655718
rect 258294 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 258914 655634
rect 258294 619954 258914 655398
rect 258294 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 258914 619954
rect 258294 619634 258914 619718
rect 258294 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 258914 619634
rect 258294 583954 258914 619398
rect 258294 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 258914 583954
rect 258294 583634 258914 583718
rect 258294 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 258914 583634
rect 258294 547954 258914 583398
rect 258294 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 258914 547954
rect 258294 547634 258914 547718
rect 258294 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 258914 547634
rect 258294 511954 258914 547398
rect 258294 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 258914 511954
rect 258294 511634 258914 511718
rect 258294 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 258914 511634
rect 258294 475954 258914 511398
rect 258294 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 258914 475954
rect 258294 475634 258914 475718
rect 258294 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 258914 475634
rect 258294 439954 258914 475398
rect 258294 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 258914 439954
rect 258294 439634 258914 439718
rect 258294 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 258914 439634
rect 258294 403954 258914 439398
rect 258294 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 258914 403954
rect 258294 403634 258914 403718
rect 258294 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 258914 403634
rect 258294 367954 258914 403398
rect 258294 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 258914 367954
rect 258294 367634 258914 367718
rect 258294 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 258914 367634
rect 258294 331954 258914 367398
rect 258294 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 258914 331954
rect 258294 331634 258914 331718
rect 258294 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 258914 331634
rect 258294 295954 258914 331398
rect 258294 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 258914 295954
rect 258294 295634 258914 295718
rect 258294 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 258914 295634
rect 258294 259954 258914 295398
rect 258294 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 258914 259954
rect 258294 259634 258914 259718
rect 258294 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 258914 259634
rect 258294 248684 258914 259398
rect 262794 706758 263414 711590
rect 262794 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 263414 706758
rect 262794 706438 263414 706522
rect 262794 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 263414 706438
rect 262794 696454 263414 706202
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 660454 263414 695898
rect 262794 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 263414 660454
rect 262794 660134 263414 660218
rect 262794 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 263414 660134
rect 262794 624454 263414 659898
rect 262794 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 263414 624454
rect 262794 624134 263414 624218
rect 262794 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 263414 624134
rect 262794 588454 263414 623898
rect 262794 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 263414 588454
rect 262794 588134 263414 588218
rect 262794 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 263414 588134
rect 262794 552454 263414 587898
rect 262794 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 263414 552454
rect 262794 552134 263414 552218
rect 262794 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 263414 552134
rect 262794 516454 263414 551898
rect 262794 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 263414 516454
rect 262794 516134 263414 516218
rect 262794 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 263414 516134
rect 262794 480454 263414 515898
rect 262794 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 263414 480454
rect 262794 480134 263414 480218
rect 262794 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 263414 480134
rect 262794 444454 263414 479898
rect 262794 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 263414 444454
rect 262794 444134 263414 444218
rect 262794 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 263414 444134
rect 262794 408454 263414 443898
rect 262794 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 263414 408454
rect 262794 408134 263414 408218
rect 262794 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 263414 408134
rect 262794 372454 263414 407898
rect 262794 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 263414 372454
rect 262794 372134 263414 372218
rect 262794 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 263414 372134
rect 262794 336454 263414 371898
rect 262794 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 263414 336454
rect 262794 336134 263414 336218
rect 262794 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 263414 336134
rect 262794 300454 263414 335898
rect 262794 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 263414 300454
rect 262794 300134 263414 300218
rect 262794 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 263414 300134
rect 262794 264454 263414 299898
rect 262794 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 263414 264454
rect 262794 264134 263414 264218
rect 262794 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 263414 264134
rect 262794 248684 263414 263898
rect 267294 707718 267914 711590
rect 267294 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 267914 707718
rect 267294 707398 267914 707482
rect 267294 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 267914 707398
rect 267294 700954 267914 707162
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 664954 267914 700398
rect 267294 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 267914 664954
rect 267294 664634 267914 664718
rect 267294 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 267914 664634
rect 267294 628954 267914 664398
rect 267294 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 267914 628954
rect 267294 628634 267914 628718
rect 267294 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 267914 628634
rect 267294 592954 267914 628398
rect 267294 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 267914 592954
rect 267294 592634 267914 592718
rect 267294 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 267914 592634
rect 267294 556954 267914 592398
rect 267294 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 267914 556954
rect 267294 556634 267914 556718
rect 267294 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 267914 556634
rect 267294 520954 267914 556398
rect 267294 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 267914 520954
rect 267294 520634 267914 520718
rect 267294 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 267914 520634
rect 267294 484954 267914 520398
rect 267294 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 267914 484954
rect 267294 484634 267914 484718
rect 267294 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 267914 484634
rect 267294 448954 267914 484398
rect 267294 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 267914 448954
rect 267294 448634 267914 448718
rect 267294 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 267914 448634
rect 267294 412954 267914 448398
rect 267294 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 267914 412954
rect 267294 412634 267914 412718
rect 267294 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 267914 412634
rect 267294 376954 267914 412398
rect 267294 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 267914 376954
rect 267294 376634 267914 376718
rect 267294 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 267914 376634
rect 267294 340954 267914 376398
rect 267294 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 267914 340954
rect 267294 340634 267914 340718
rect 267294 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 267914 340634
rect 267294 304954 267914 340398
rect 267294 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 267914 304954
rect 267294 304634 267914 304718
rect 267294 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 267914 304634
rect 267294 268954 267914 304398
rect 267294 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 267914 268954
rect 267294 268634 267914 268718
rect 267294 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 267914 268634
rect 267294 248684 267914 268398
rect 271794 708678 272414 711590
rect 271794 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 272414 708678
rect 271794 708358 272414 708442
rect 271794 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 272414 708358
rect 271794 669454 272414 708122
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 248684 272414 272898
rect 276294 709638 276914 711590
rect 276294 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 276914 709638
rect 276294 709318 276914 709402
rect 276294 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 276914 709318
rect 276294 673954 276914 709082
rect 276294 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 276914 673954
rect 276294 673634 276914 673718
rect 276294 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 276914 673634
rect 276294 637954 276914 673398
rect 276294 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 276914 637954
rect 276294 637634 276914 637718
rect 276294 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 276914 637634
rect 276294 601954 276914 637398
rect 276294 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 276914 601954
rect 276294 601634 276914 601718
rect 276294 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 276914 601634
rect 276294 565954 276914 601398
rect 276294 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 276914 565954
rect 276294 565634 276914 565718
rect 276294 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 276914 565634
rect 276294 529954 276914 565398
rect 276294 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 276914 529954
rect 276294 529634 276914 529718
rect 276294 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 276914 529634
rect 276294 493954 276914 529398
rect 276294 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 276914 493954
rect 276294 493634 276914 493718
rect 276294 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 276914 493634
rect 276294 457954 276914 493398
rect 276294 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 276914 457954
rect 276294 457634 276914 457718
rect 276294 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 276914 457634
rect 276294 421954 276914 457398
rect 276294 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 276914 421954
rect 276294 421634 276914 421718
rect 276294 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 276914 421634
rect 276294 385954 276914 421398
rect 276294 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 276914 385954
rect 276294 385634 276914 385718
rect 276294 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 276914 385634
rect 276294 349954 276914 385398
rect 276294 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 276914 349954
rect 276294 349634 276914 349718
rect 276294 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 276914 349634
rect 276294 313954 276914 349398
rect 276294 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 276914 313954
rect 276294 313634 276914 313718
rect 276294 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 276914 313634
rect 276294 277954 276914 313398
rect 276294 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 276914 277954
rect 276294 277634 276914 277718
rect 276294 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 276914 277634
rect 276294 248684 276914 277398
rect 280794 710598 281414 711590
rect 280794 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 281414 710598
rect 280794 710278 281414 710362
rect 280794 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 281414 710278
rect 280794 678454 281414 710042
rect 280794 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 281414 678454
rect 280794 678134 281414 678218
rect 280794 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 281414 678134
rect 280794 642454 281414 677898
rect 280794 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 281414 642454
rect 280794 642134 281414 642218
rect 280794 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 281414 642134
rect 280794 606454 281414 641898
rect 280794 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 281414 606454
rect 280794 606134 281414 606218
rect 280794 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 281414 606134
rect 280794 570454 281414 605898
rect 280794 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 281414 570454
rect 280794 570134 281414 570218
rect 280794 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 281414 570134
rect 280794 534454 281414 569898
rect 280794 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 281414 534454
rect 280794 534134 281414 534218
rect 280794 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 281414 534134
rect 280794 498454 281414 533898
rect 280794 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 281414 498454
rect 280794 498134 281414 498218
rect 280794 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 281414 498134
rect 280794 462454 281414 497898
rect 280794 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 281414 462454
rect 280794 462134 281414 462218
rect 280794 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 281414 462134
rect 280794 426454 281414 461898
rect 280794 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 281414 426454
rect 280794 426134 281414 426218
rect 280794 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 281414 426134
rect 280794 390454 281414 425898
rect 280794 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 281414 390454
rect 280794 390134 281414 390218
rect 280794 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 281414 390134
rect 280794 354454 281414 389898
rect 280794 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 281414 354454
rect 280794 354134 281414 354218
rect 280794 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 281414 354134
rect 280794 318454 281414 353898
rect 280794 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 281414 318454
rect 280794 318134 281414 318218
rect 280794 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 281414 318134
rect 280794 282454 281414 317898
rect 280794 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 281414 282454
rect 280794 282134 281414 282218
rect 280794 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 281414 282134
rect 280794 248684 281414 281898
rect 285294 711558 285914 711590
rect 285294 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 285914 711558
rect 285294 711238 285914 711322
rect 285294 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 285914 711238
rect 285294 682954 285914 711002
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 285294 646954 285914 682398
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 285294 610954 285914 646398
rect 285294 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 285914 610954
rect 285294 610634 285914 610718
rect 285294 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 285914 610634
rect 285294 574954 285914 610398
rect 285294 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 285914 574954
rect 285294 574634 285914 574718
rect 285294 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 285914 574634
rect 285294 538954 285914 574398
rect 285294 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 285914 538954
rect 285294 538634 285914 538718
rect 285294 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 285914 538634
rect 285294 502954 285914 538398
rect 285294 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 285914 502954
rect 285294 502634 285914 502718
rect 285294 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 285914 502634
rect 285294 466954 285914 502398
rect 285294 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 285914 466954
rect 285294 466634 285914 466718
rect 285294 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 285914 466634
rect 285294 430954 285914 466398
rect 285294 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 285914 430954
rect 285294 430634 285914 430718
rect 285294 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 285914 430634
rect 285294 394954 285914 430398
rect 285294 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 285914 394954
rect 285294 394634 285914 394718
rect 285294 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 285914 394634
rect 285294 358954 285914 394398
rect 285294 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 285914 358954
rect 285294 358634 285914 358718
rect 285294 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 285914 358634
rect 285294 322954 285914 358398
rect 285294 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 285914 322954
rect 285294 322634 285914 322718
rect 285294 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 285914 322634
rect 285294 286954 285914 322398
rect 285294 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 285914 286954
rect 285294 286634 285914 286718
rect 285294 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 285914 286634
rect 285294 250954 285914 286398
rect 285294 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 285914 250954
rect 285294 250634 285914 250718
rect 285294 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 285914 250634
rect 285294 248684 285914 250398
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 248684 290414 254898
rect 294294 705798 294914 711590
rect 294294 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 294914 705798
rect 294294 705478 294914 705562
rect 294294 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 294914 705478
rect 294294 691954 294914 705242
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 619954 294914 655398
rect 294294 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 294914 619954
rect 294294 619634 294914 619718
rect 294294 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 294914 619634
rect 294294 583954 294914 619398
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 294294 547954 294914 583398
rect 294294 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 294914 547954
rect 294294 547634 294914 547718
rect 294294 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 294914 547634
rect 294294 511954 294914 547398
rect 294294 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 294914 511954
rect 294294 511634 294914 511718
rect 294294 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 294914 511634
rect 294294 475954 294914 511398
rect 294294 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 294914 475954
rect 294294 475634 294914 475718
rect 294294 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 294914 475634
rect 294294 439954 294914 475398
rect 294294 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 294914 439954
rect 294294 439634 294914 439718
rect 294294 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 294914 439634
rect 294294 403954 294914 439398
rect 294294 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 294914 403954
rect 294294 403634 294914 403718
rect 294294 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 294914 403634
rect 294294 367954 294914 403398
rect 294294 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 294914 367954
rect 294294 367634 294914 367718
rect 294294 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 294914 367634
rect 294294 331954 294914 367398
rect 294294 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 294914 331954
rect 294294 331634 294914 331718
rect 294294 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 294914 331634
rect 294294 295954 294914 331398
rect 294294 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 294914 295954
rect 294294 295634 294914 295718
rect 294294 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 294914 295634
rect 294294 259954 294914 295398
rect 294294 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 294914 259954
rect 294294 259634 294914 259718
rect 294294 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 294914 259634
rect 294294 248684 294914 259398
rect 298794 706758 299414 711590
rect 298794 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 299414 706758
rect 298794 706438 299414 706522
rect 298794 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 299414 706438
rect 298794 696454 299414 706202
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 660454 299414 695898
rect 298794 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 299414 660454
rect 298794 660134 299414 660218
rect 298794 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 299414 660134
rect 298794 624454 299414 659898
rect 298794 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 299414 624454
rect 298794 624134 299414 624218
rect 298794 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 299414 624134
rect 298794 588454 299414 623898
rect 298794 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 299414 588454
rect 298794 588134 299414 588218
rect 298794 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 299414 588134
rect 298794 552454 299414 587898
rect 298794 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 299414 552454
rect 298794 552134 299414 552218
rect 298794 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 299414 552134
rect 298794 516454 299414 551898
rect 298794 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 299414 516454
rect 298794 516134 299414 516218
rect 298794 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 299414 516134
rect 298794 480454 299414 515898
rect 298794 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 299414 480454
rect 298794 480134 299414 480218
rect 298794 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 299414 480134
rect 298794 444454 299414 479898
rect 298794 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 299414 444454
rect 298794 444134 299414 444218
rect 298794 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 299414 444134
rect 298794 408454 299414 443898
rect 298794 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 299414 408454
rect 298794 408134 299414 408218
rect 298794 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 299414 408134
rect 298794 372454 299414 407898
rect 298794 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 299414 372454
rect 298794 372134 299414 372218
rect 298794 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 299414 372134
rect 298794 336454 299414 371898
rect 298794 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 299414 336454
rect 298794 336134 299414 336218
rect 298794 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 299414 336134
rect 298794 300454 299414 335898
rect 298794 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 299414 300454
rect 298794 300134 299414 300218
rect 298794 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 299414 300134
rect 298794 264454 299414 299898
rect 298794 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 299414 264454
rect 298794 264134 299414 264218
rect 298794 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 299414 264134
rect 298794 248684 299414 263898
rect 303294 707718 303914 711590
rect 303294 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 303914 707718
rect 303294 707398 303914 707482
rect 303294 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 303914 707398
rect 303294 700954 303914 707162
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 664954 303914 700398
rect 303294 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 303914 664954
rect 303294 664634 303914 664718
rect 303294 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 303914 664634
rect 303294 628954 303914 664398
rect 303294 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 303914 628954
rect 303294 628634 303914 628718
rect 303294 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 303914 628634
rect 303294 592954 303914 628398
rect 303294 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 303914 592954
rect 303294 592634 303914 592718
rect 303294 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 303914 592634
rect 303294 556954 303914 592398
rect 303294 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 303914 556954
rect 303294 556634 303914 556718
rect 303294 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 303914 556634
rect 303294 520954 303914 556398
rect 303294 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 303914 520954
rect 303294 520634 303914 520718
rect 303294 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 303914 520634
rect 303294 484954 303914 520398
rect 303294 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 303914 484954
rect 303294 484634 303914 484718
rect 303294 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 303914 484634
rect 303294 448954 303914 484398
rect 303294 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 303914 448954
rect 303294 448634 303914 448718
rect 303294 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 303914 448634
rect 303294 412954 303914 448398
rect 303294 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 303914 412954
rect 303294 412634 303914 412718
rect 303294 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 303914 412634
rect 303294 376954 303914 412398
rect 303294 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 303914 376954
rect 303294 376634 303914 376718
rect 303294 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 303914 376634
rect 303294 340954 303914 376398
rect 303294 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 303914 340954
rect 303294 340634 303914 340718
rect 303294 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 303914 340634
rect 303294 304954 303914 340398
rect 303294 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 303914 304954
rect 303294 304634 303914 304718
rect 303294 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 303914 304634
rect 303294 268954 303914 304398
rect 303294 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 303914 268954
rect 303294 268634 303914 268718
rect 303294 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 303914 268634
rect 303294 248684 303914 268398
rect 307794 708678 308414 711590
rect 307794 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 308414 708678
rect 307794 708358 308414 708442
rect 307794 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 308414 708358
rect 307794 669454 308414 708122
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 248684 308414 272898
rect 312294 709638 312914 711590
rect 312294 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 312914 709638
rect 312294 709318 312914 709402
rect 312294 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 312914 709318
rect 312294 673954 312914 709082
rect 312294 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 312914 673954
rect 312294 673634 312914 673718
rect 312294 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 312914 673634
rect 312294 637954 312914 673398
rect 312294 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 312914 637954
rect 312294 637634 312914 637718
rect 312294 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 312914 637634
rect 312294 601954 312914 637398
rect 312294 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 312914 601954
rect 312294 601634 312914 601718
rect 312294 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 312914 601634
rect 312294 565954 312914 601398
rect 312294 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 312914 565954
rect 312294 565634 312914 565718
rect 312294 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 312914 565634
rect 312294 529954 312914 565398
rect 312294 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 312914 529954
rect 312294 529634 312914 529718
rect 312294 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 312914 529634
rect 312294 493954 312914 529398
rect 312294 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 312914 493954
rect 312294 493634 312914 493718
rect 312294 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 312914 493634
rect 312294 457954 312914 493398
rect 312294 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 312914 457954
rect 312294 457634 312914 457718
rect 312294 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 312914 457634
rect 312294 421954 312914 457398
rect 312294 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 312914 421954
rect 312294 421634 312914 421718
rect 312294 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 312914 421634
rect 312294 385954 312914 421398
rect 312294 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 312914 385954
rect 312294 385634 312914 385718
rect 312294 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 312914 385634
rect 312294 349954 312914 385398
rect 312294 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 312914 349954
rect 312294 349634 312914 349718
rect 312294 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 312914 349634
rect 312294 313954 312914 349398
rect 312294 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 312914 313954
rect 312294 313634 312914 313718
rect 312294 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 312914 313634
rect 312294 277954 312914 313398
rect 312294 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 312914 277954
rect 312294 277634 312914 277718
rect 312294 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 312914 277634
rect 312294 248684 312914 277398
rect 316794 710598 317414 711590
rect 316794 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 317414 710598
rect 316794 710278 317414 710362
rect 316794 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 317414 710278
rect 316794 678454 317414 710042
rect 316794 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 317414 678454
rect 316794 678134 317414 678218
rect 316794 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 317414 678134
rect 316794 642454 317414 677898
rect 316794 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 317414 642454
rect 316794 642134 317414 642218
rect 316794 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 317414 642134
rect 316794 606454 317414 641898
rect 316794 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 317414 606454
rect 316794 606134 317414 606218
rect 316794 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 317414 606134
rect 316794 570454 317414 605898
rect 316794 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 317414 570454
rect 316794 570134 317414 570218
rect 316794 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 317414 570134
rect 316794 534454 317414 569898
rect 316794 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 317414 534454
rect 316794 534134 317414 534218
rect 316794 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 317414 534134
rect 316794 498454 317414 533898
rect 316794 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 317414 498454
rect 316794 498134 317414 498218
rect 316794 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 317414 498134
rect 316794 462454 317414 497898
rect 316794 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 317414 462454
rect 316794 462134 317414 462218
rect 316794 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 317414 462134
rect 316794 426454 317414 461898
rect 316794 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 317414 426454
rect 316794 426134 317414 426218
rect 316794 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 317414 426134
rect 316794 390454 317414 425898
rect 316794 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 317414 390454
rect 316794 390134 317414 390218
rect 316794 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 317414 390134
rect 316794 354454 317414 389898
rect 316794 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 317414 354454
rect 316794 354134 317414 354218
rect 316794 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 317414 354134
rect 316794 318454 317414 353898
rect 316794 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 317414 318454
rect 316794 318134 317414 318218
rect 316794 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 317414 318134
rect 316794 282454 317414 317898
rect 316794 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 317414 282454
rect 316794 282134 317414 282218
rect 316794 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 317414 282134
rect 316794 248684 317414 281898
rect 321294 711558 321914 711590
rect 321294 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 321914 711558
rect 321294 711238 321914 711322
rect 321294 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 321914 711238
rect 321294 682954 321914 711002
rect 321294 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 321914 682954
rect 321294 682634 321914 682718
rect 321294 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 321914 682634
rect 321294 646954 321914 682398
rect 321294 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 321914 646954
rect 321294 646634 321914 646718
rect 321294 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 321914 646634
rect 321294 610954 321914 646398
rect 321294 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 321914 610954
rect 321294 610634 321914 610718
rect 321294 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 321914 610634
rect 321294 574954 321914 610398
rect 321294 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 321914 574954
rect 321294 574634 321914 574718
rect 321294 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 321914 574634
rect 321294 538954 321914 574398
rect 321294 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 321914 538954
rect 321294 538634 321914 538718
rect 321294 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 321914 538634
rect 321294 502954 321914 538398
rect 321294 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 321914 502954
rect 321294 502634 321914 502718
rect 321294 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 321914 502634
rect 321294 466954 321914 502398
rect 321294 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 321914 466954
rect 321294 466634 321914 466718
rect 321294 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 321914 466634
rect 321294 430954 321914 466398
rect 321294 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 321914 430954
rect 321294 430634 321914 430718
rect 321294 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 321914 430634
rect 321294 394954 321914 430398
rect 321294 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 321914 394954
rect 321294 394634 321914 394718
rect 321294 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 321914 394634
rect 321294 358954 321914 394398
rect 321294 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 321914 358954
rect 321294 358634 321914 358718
rect 321294 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 321914 358634
rect 321294 322954 321914 358398
rect 321294 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 321914 322954
rect 321294 322634 321914 322718
rect 321294 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 321914 322634
rect 321294 286954 321914 322398
rect 321294 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 321914 286954
rect 321294 286634 321914 286718
rect 321294 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 321914 286634
rect 321294 250954 321914 286398
rect 321294 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 321914 250954
rect 321294 250634 321914 250718
rect 321294 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 321914 250634
rect 321294 248684 321914 250398
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 248684 326414 254898
rect 330294 705798 330914 711590
rect 330294 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 330914 705798
rect 330294 705478 330914 705562
rect 330294 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 330914 705478
rect 330294 691954 330914 705242
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 655954 330914 691398
rect 330294 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 330914 655954
rect 330294 655634 330914 655718
rect 330294 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 330914 655634
rect 330294 619954 330914 655398
rect 330294 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 330914 619954
rect 330294 619634 330914 619718
rect 330294 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 330914 619634
rect 330294 583954 330914 619398
rect 330294 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 330914 583954
rect 330294 583634 330914 583718
rect 330294 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 330914 583634
rect 330294 547954 330914 583398
rect 330294 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 330914 547954
rect 330294 547634 330914 547718
rect 330294 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 330914 547634
rect 330294 511954 330914 547398
rect 330294 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 330914 511954
rect 330294 511634 330914 511718
rect 330294 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 330914 511634
rect 330294 475954 330914 511398
rect 330294 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 330914 475954
rect 330294 475634 330914 475718
rect 330294 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 330914 475634
rect 330294 439954 330914 475398
rect 330294 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 330914 439954
rect 330294 439634 330914 439718
rect 330294 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 330914 439634
rect 330294 403954 330914 439398
rect 330294 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 330914 403954
rect 330294 403634 330914 403718
rect 330294 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 330914 403634
rect 330294 367954 330914 403398
rect 330294 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 330914 367954
rect 330294 367634 330914 367718
rect 330294 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 330914 367634
rect 330294 331954 330914 367398
rect 330294 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 330914 331954
rect 330294 331634 330914 331718
rect 330294 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 330914 331634
rect 330294 295954 330914 331398
rect 330294 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 330914 295954
rect 330294 295634 330914 295718
rect 330294 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 330914 295634
rect 330294 259954 330914 295398
rect 330294 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 330914 259954
rect 330294 259634 330914 259718
rect 330294 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 330914 259634
rect 330294 248684 330914 259398
rect 334794 706758 335414 711590
rect 334794 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 335414 706758
rect 334794 706438 335414 706522
rect 334794 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 335414 706438
rect 334794 696454 335414 706202
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 660454 335414 695898
rect 334794 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 335414 660454
rect 334794 660134 335414 660218
rect 334794 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 335414 660134
rect 334794 624454 335414 659898
rect 334794 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 335414 624454
rect 334794 624134 335414 624218
rect 334794 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 335414 624134
rect 334794 588454 335414 623898
rect 334794 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 335414 588454
rect 334794 588134 335414 588218
rect 334794 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 335414 588134
rect 334794 552454 335414 587898
rect 334794 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 335414 552454
rect 334794 552134 335414 552218
rect 334794 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 335414 552134
rect 334794 516454 335414 551898
rect 334794 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 335414 516454
rect 334794 516134 335414 516218
rect 334794 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 335414 516134
rect 334794 480454 335414 515898
rect 334794 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 335414 480454
rect 334794 480134 335414 480218
rect 334794 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 335414 480134
rect 334794 444454 335414 479898
rect 334794 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 335414 444454
rect 334794 444134 335414 444218
rect 334794 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 335414 444134
rect 334794 408454 335414 443898
rect 334794 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 335414 408454
rect 334794 408134 335414 408218
rect 334794 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 335414 408134
rect 334794 372454 335414 407898
rect 334794 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 335414 372454
rect 334794 372134 335414 372218
rect 334794 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 335414 372134
rect 334794 336454 335414 371898
rect 334794 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 335414 336454
rect 334794 336134 335414 336218
rect 334794 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 335414 336134
rect 334794 300454 335414 335898
rect 334794 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 335414 300454
rect 334794 300134 335414 300218
rect 334794 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 335414 300134
rect 334794 264454 335414 299898
rect 334794 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 335414 264454
rect 334794 264134 335414 264218
rect 334794 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 335414 264134
rect 334794 248684 335414 263898
rect 339294 707718 339914 711590
rect 339294 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 339914 707718
rect 339294 707398 339914 707482
rect 339294 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 339914 707398
rect 339294 700954 339914 707162
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 664954 339914 700398
rect 339294 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 339914 664954
rect 339294 664634 339914 664718
rect 339294 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 339914 664634
rect 339294 628954 339914 664398
rect 339294 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 339914 628954
rect 339294 628634 339914 628718
rect 339294 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 339914 628634
rect 339294 592954 339914 628398
rect 339294 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 339914 592954
rect 339294 592634 339914 592718
rect 339294 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 339914 592634
rect 339294 556954 339914 592398
rect 339294 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 339914 556954
rect 339294 556634 339914 556718
rect 339294 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 339914 556634
rect 339294 520954 339914 556398
rect 339294 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 339914 520954
rect 339294 520634 339914 520718
rect 339294 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 339914 520634
rect 339294 484954 339914 520398
rect 339294 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 339914 484954
rect 339294 484634 339914 484718
rect 339294 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 339914 484634
rect 339294 448954 339914 484398
rect 339294 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 339914 448954
rect 339294 448634 339914 448718
rect 339294 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 339914 448634
rect 339294 412954 339914 448398
rect 339294 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 339914 412954
rect 339294 412634 339914 412718
rect 339294 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 339914 412634
rect 339294 376954 339914 412398
rect 339294 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 339914 376954
rect 339294 376634 339914 376718
rect 339294 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 339914 376634
rect 339294 340954 339914 376398
rect 339294 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 339914 340954
rect 339294 340634 339914 340718
rect 339294 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 339914 340634
rect 339294 304954 339914 340398
rect 339294 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 339914 304954
rect 339294 304634 339914 304718
rect 339294 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 339914 304634
rect 339294 268954 339914 304398
rect 339294 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 339914 268954
rect 339294 268634 339914 268718
rect 339294 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 339914 268634
rect 339294 248684 339914 268398
rect 343794 708678 344414 711590
rect 343794 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 344414 708678
rect 343794 708358 344414 708442
rect 343794 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 344414 708358
rect 343794 669454 344414 708122
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 248684 344414 272898
rect 348294 709638 348914 711590
rect 348294 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 348914 709638
rect 348294 709318 348914 709402
rect 348294 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 348914 709318
rect 348294 673954 348914 709082
rect 348294 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 348914 673954
rect 348294 673634 348914 673718
rect 348294 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 348914 673634
rect 348294 637954 348914 673398
rect 348294 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 348914 637954
rect 348294 637634 348914 637718
rect 348294 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 348914 637634
rect 348294 601954 348914 637398
rect 348294 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 348914 601954
rect 348294 601634 348914 601718
rect 348294 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 348914 601634
rect 348294 565954 348914 601398
rect 348294 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 348914 565954
rect 348294 565634 348914 565718
rect 348294 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 348914 565634
rect 348294 529954 348914 565398
rect 348294 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 348914 529954
rect 348294 529634 348914 529718
rect 348294 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 348914 529634
rect 348294 493954 348914 529398
rect 348294 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 348914 493954
rect 348294 493634 348914 493718
rect 348294 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 348914 493634
rect 348294 457954 348914 493398
rect 348294 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 348914 457954
rect 348294 457634 348914 457718
rect 348294 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 348914 457634
rect 348294 421954 348914 457398
rect 348294 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 348914 421954
rect 348294 421634 348914 421718
rect 348294 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 348914 421634
rect 348294 385954 348914 421398
rect 348294 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 348914 385954
rect 348294 385634 348914 385718
rect 348294 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 348914 385634
rect 348294 349954 348914 385398
rect 348294 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 348914 349954
rect 348294 349634 348914 349718
rect 348294 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 348914 349634
rect 348294 313954 348914 349398
rect 348294 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 348914 313954
rect 348294 313634 348914 313718
rect 348294 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 348914 313634
rect 348294 277954 348914 313398
rect 348294 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 348914 277954
rect 348294 277634 348914 277718
rect 348294 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 348914 277634
rect 348294 248684 348914 277398
rect 352794 710598 353414 711590
rect 352794 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 353414 710598
rect 352794 710278 353414 710362
rect 352794 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 353414 710278
rect 352794 678454 353414 710042
rect 352794 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 353414 678454
rect 352794 678134 353414 678218
rect 352794 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 353414 678134
rect 352794 642454 353414 677898
rect 352794 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 353414 642454
rect 352794 642134 353414 642218
rect 352794 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 353414 642134
rect 352794 606454 353414 641898
rect 352794 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 353414 606454
rect 352794 606134 353414 606218
rect 352794 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 353414 606134
rect 352794 570454 353414 605898
rect 352794 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 353414 570454
rect 352794 570134 353414 570218
rect 352794 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 353414 570134
rect 352794 534454 353414 569898
rect 352794 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 353414 534454
rect 352794 534134 353414 534218
rect 352794 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 353414 534134
rect 352794 498454 353414 533898
rect 352794 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 353414 498454
rect 352794 498134 353414 498218
rect 352794 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 353414 498134
rect 352794 462454 353414 497898
rect 352794 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 353414 462454
rect 352794 462134 353414 462218
rect 352794 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 353414 462134
rect 352794 426454 353414 461898
rect 352794 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 353414 426454
rect 352794 426134 353414 426218
rect 352794 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 353414 426134
rect 352794 390454 353414 425898
rect 352794 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 353414 390454
rect 352794 390134 353414 390218
rect 352794 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 353414 390134
rect 352794 354454 353414 389898
rect 352794 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 353414 354454
rect 352794 354134 353414 354218
rect 352794 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 353414 354134
rect 352794 318454 353414 353898
rect 352794 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 353414 318454
rect 352794 318134 353414 318218
rect 352794 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 353414 318134
rect 352794 282454 353414 317898
rect 352794 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 353414 282454
rect 352794 282134 353414 282218
rect 352794 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 353414 282134
rect 352794 248684 353414 281898
rect 357294 711558 357914 711590
rect 357294 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 357914 711558
rect 357294 711238 357914 711322
rect 357294 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 357914 711238
rect 357294 682954 357914 711002
rect 357294 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 357914 682954
rect 357294 682634 357914 682718
rect 357294 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 357914 682634
rect 357294 646954 357914 682398
rect 357294 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 357914 646954
rect 357294 646634 357914 646718
rect 357294 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 357914 646634
rect 357294 610954 357914 646398
rect 357294 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 357914 610954
rect 357294 610634 357914 610718
rect 357294 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 357914 610634
rect 357294 574954 357914 610398
rect 357294 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 357914 574954
rect 357294 574634 357914 574718
rect 357294 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 357914 574634
rect 357294 538954 357914 574398
rect 357294 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 357914 538954
rect 357294 538634 357914 538718
rect 357294 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 357914 538634
rect 357294 502954 357914 538398
rect 357294 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 357914 502954
rect 357294 502634 357914 502718
rect 357294 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 357914 502634
rect 357294 466954 357914 502398
rect 357294 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 357914 466954
rect 357294 466634 357914 466718
rect 357294 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 357914 466634
rect 357294 430954 357914 466398
rect 357294 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 357914 430954
rect 357294 430634 357914 430718
rect 357294 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 357914 430634
rect 357294 394954 357914 430398
rect 357294 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 357914 394954
rect 357294 394634 357914 394718
rect 357294 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 357914 394634
rect 357294 358954 357914 394398
rect 357294 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 357914 358954
rect 357294 358634 357914 358718
rect 357294 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 357914 358634
rect 357294 322954 357914 358398
rect 357294 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 357914 322954
rect 357294 322634 357914 322718
rect 357294 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 357914 322634
rect 357294 286954 357914 322398
rect 357294 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 357914 286954
rect 357294 286634 357914 286718
rect 357294 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 357914 286634
rect 357294 250954 357914 286398
rect 357294 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 357914 250954
rect 357294 250634 357914 250718
rect 357294 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 357914 250634
rect 357294 248684 357914 250398
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 248684 362414 254898
rect 366294 705798 366914 711590
rect 366294 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 366914 705798
rect 366294 705478 366914 705562
rect 366294 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 366914 705478
rect 366294 691954 366914 705242
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 655954 366914 691398
rect 366294 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 366914 655954
rect 366294 655634 366914 655718
rect 366294 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 366914 655634
rect 366294 619954 366914 655398
rect 366294 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 366914 619954
rect 366294 619634 366914 619718
rect 366294 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 366914 619634
rect 366294 583954 366914 619398
rect 366294 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 366914 583954
rect 366294 583634 366914 583718
rect 366294 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 366914 583634
rect 366294 547954 366914 583398
rect 366294 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 366914 547954
rect 366294 547634 366914 547718
rect 366294 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 366914 547634
rect 366294 511954 366914 547398
rect 366294 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 366914 511954
rect 366294 511634 366914 511718
rect 366294 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 366914 511634
rect 366294 475954 366914 511398
rect 366294 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 366914 475954
rect 366294 475634 366914 475718
rect 366294 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 366914 475634
rect 366294 439954 366914 475398
rect 366294 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 366914 439954
rect 366294 439634 366914 439718
rect 366294 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 366914 439634
rect 366294 403954 366914 439398
rect 366294 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 366914 403954
rect 366294 403634 366914 403718
rect 366294 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 366914 403634
rect 366294 367954 366914 403398
rect 366294 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 366914 367954
rect 366294 367634 366914 367718
rect 366294 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 366914 367634
rect 366294 331954 366914 367398
rect 366294 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 366914 331954
rect 366294 331634 366914 331718
rect 366294 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 366914 331634
rect 366294 295954 366914 331398
rect 366294 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 366914 295954
rect 366294 295634 366914 295718
rect 366294 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 366914 295634
rect 366294 259954 366914 295398
rect 366294 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 366914 259954
rect 366294 259634 366914 259718
rect 366294 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 366914 259634
rect 366294 248684 366914 259398
rect 370794 706758 371414 711590
rect 370794 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 371414 706758
rect 370794 706438 371414 706522
rect 370794 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 371414 706438
rect 370794 696454 371414 706202
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 660454 371414 695898
rect 370794 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 371414 660454
rect 370794 660134 371414 660218
rect 370794 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 371414 660134
rect 370794 624454 371414 659898
rect 370794 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 371414 624454
rect 370794 624134 371414 624218
rect 370794 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 371414 624134
rect 370794 588454 371414 623898
rect 370794 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 371414 588454
rect 370794 588134 371414 588218
rect 370794 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 371414 588134
rect 370794 552454 371414 587898
rect 370794 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 371414 552454
rect 370794 552134 371414 552218
rect 370794 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 371414 552134
rect 370794 516454 371414 551898
rect 370794 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 371414 516454
rect 370794 516134 371414 516218
rect 370794 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 371414 516134
rect 370794 480454 371414 515898
rect 370794 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 371414 480454
rect 370794 480134 371414 480218
rect 370794 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 371414 480134
rect 370794 444454 371414 479898
rect 370794 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 371414 444454
rect 370794 444134 371414 444218
rect 370794 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 371414 444134
rect 370794 408454 371414 443898
rect 370794 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 371414 408454
rect 370794 408134 371414 408218
rect 370794 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 371414 408134
rect 370794 372454 371414 407898
rect 370794 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 371414 372454
rect 370794 372134 371414 372218
rect 370794 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 371414 372134
rect 370794 336454 371414 371898
rect 370794 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 371414 336454
rect 370794 336134 371414 336218
rect 370794 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 371414 336134
rect 370794 300454 371414 335898
rect 370794 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 371414 300454
rect 370794 300134 371414 300218
rect 370794 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 371414 300134
rect 370794 264454 371414 299898
rect 370794 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 371414 264454
rect 370794 264134 371414 264218
rect 370794 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 371414 264134
rect 370794 248684 371414 263898
rect 375294 707718 375914 711590
rect 375294 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 375914 707718
rect 375294 707398 375914 707482
rect 375294 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 375914 707398
rect 375294 700954 375914 707162
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 664954 375914 700398
rect 375294 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 375914 664954
rect 375294 664634 375914 664718
rect 375294 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 375914 664634
rect 375294 628954 375914 664398
rect 375294 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 375914 628954
rect 375294 628634 375914 628718
rect 375294 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 375914 628634
rect 375294 592954 375914 628398
rect 375294 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 375914 592954
rect 375294 592634 375914 592718
rect 375294 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 375914 592634
rect 375294 556954 375914 592398
rect 375294 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 375914 556954
rect 375294 556634 375914 556718
rect 375294 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 375914 556634
rect 375294 520954 375914 556398
rect 375294 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 375914 520954
rect 375294 520634 375914 520718
rect 375294 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 375914 520634
rect 375294 484954 375914 520398
rect 375294 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 375914 484954
rect 375294 484634 375914 484718
rect 375294 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 375914 484634
rect 375294 448954 375914 484398
rect 375294 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 375914 448954
rect 375294 448634 375914 448718
rect 375294 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 375914 448634
rect 375294 412954 375914 448398
rect 375294 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 375914 412954
rect 375294 412634 375914 412718
rect 375294 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 375914 412634
rect 375294 376954 375914 412398
rect 375294 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 375914 376954
rect 375294 376634 375914 376718
rect 375294 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 375914 376634
rect 375294 340954 375914 376398
rect 375294 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 375914 340954
rect 375294 340634 375914 340718
rect 375294 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 375914 340634
rect 375294 304954 375914 340398
rect 375294 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 375914 304954
rect 375294 304634 375914 304718
rect 375294 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 375914 304634
rect 375294 268954 375914 304398
rect 375294 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 375914 268954
rect 375294 268634 375914 268718
rect 375294 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 375914 268634
rect 375294 248684 375914 268398
rect 379794 708678 380414 711590
rect 379794 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 380414 708678
rect 379794 708358 380414 708442
rect 379794 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 380414 708358
rect 379794 669454 380414 708122
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 248684 380414 272898
rect 384294 709638 384914 711590
rect 384294 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 384914 709638
rect 384294 709318 384914 709402
rect 384294 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 384914 709318
rect 384294 673954 384914 709082
rect 384294 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 384914 673954
rect 384294 673634 384914 673718
rect 384294 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 384914 673634
rect 384294 637954 384914 673398
rect 384294 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 384914 637954
rect 384294 637634 384914 637718
rect 384294 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 384914 637634
rect 384294 601954 384914 637398
rect 384294 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 384914 601954
rect 384294 601634 384914 601718
rect 384294 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 384914 601634
rect 384294 565954 384914 601398
rect 384294 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 384914 565954
rect 384294 565634 384914 565718
rect 384294 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 384914 565634
rect 384294 529954 384914 565398
rect 384294 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 384914 529954
rect 384294 529634 384914 529718
rect 384294 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 384914 529634
rect 384294 493954 384914 529398
rect 384294 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 384914 493954
rect 384294 493634 384914 493718
rect 384294 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 384914 493634
rect 384294 457954 384914 493398
rect 384294 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 384914 457954
rect 384294 457634 384914 457718
rect 384294 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 384914 457634
rect 384294 421954 384914 457398
rect 384294 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 384914 421954
rect 384294 421634 384914 421718
rect 384294 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 384914 421634
rect 384294 385954 384914 421398
rect 384294 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 384914 385954
rect 384294 385634 384914 385718
rect 384294 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 384914 385634
rect 384294 349954 384914 385398
rect 384294 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 384914 349954
rect 384294 349634 384914 349718
rect 384294 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 384914 349634
rect 384294 313954 384914 349398
rect 384294 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 384914 313954
rect 384294 313634 384914 313718
rect 384294 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 384914 313634
rect 384294 277954 384914 313398
rect 384294 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 384914 277954
rect 384294 277634 384914 277718
rect 384294 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 384914 277634
rect 384294 248684 384914 277398
rect 388794 710598 389414 711590
rect 388794 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 389414 710598
rect 388794 710278 389414 710362
rect 388794 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 389414 710278
rect 388794 678454 389414 710042
rect 388794 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 389414 678454
rect 388794 678134 389414 678218
rect 388794 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 389414 678134
rect 388794 642454 389414 677898
rect 388794 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 389414 642454
rect 388794 642134 389414 642218
rect 388794 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 389414 642134
rect 388794 606454 389414 641898
rect 388794 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 389414 606454
rect 388794 606134 389414 606218
rect 388794 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 389414 606134
rect 388794 570454 389414 605898
rect 388794 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 389414 570454
rect 388794 570134 389414 570218
rect 388794 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 389414 570134
rect 388794 534454 389414 569898
rect 388794 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 389414 534454
rect 388794 534134 389414 534218
rect 388794 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 389414 534134
rect 388794 498454 389414 533898
rect 388794 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 389414 498454
rect 388794 498134 389414 498218
rect 388794 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 389414 498134
rect 388794 462454 389414 497898
rect 388794 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 389414 462454
rect 388794 462134 389414 462218
rect 388794 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 389414 462134
rect 388794 426454 389414 461898
rect 388794 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 389414 426454
rect 388794 426134 389414 426218
rect 388794 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 389414 426134
rect 388794 390454 389414 425898
rect 388794 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 389414 390454
rect 388794 390134 389414 390218
rect 388794 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 389414 390134
rect 388794 354454 389414 389898
rect 388794 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 389414 354454
rect 388794 354134 389414 354218
rect 388794 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 389414 354134
rect 388794 318454 389414 353898
rect 388794 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 389414 318454
rect 388794 318134 389414 318218
rect 388794 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 389414 318134
rect 388794 282454 389414 317898
rect 388794 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 389414 282454
rect 388794 282134 389414 282218
rect 388794 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 389414 282134
rect 388794 248684 389414 281898
rect 393294 711558 393914 711590
rect 393294 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 393914 711558
rect 393294 711238 393914 711322
rect 393294 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 393914 711238
rect 393294 682954 393914 711002
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 396579 696964 396645 696965
rect 396579 696900 396580 696964
rect 396644 696900 396645 696964
rect 396579 696899 396645 696900
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 393294 646954 393914 682398
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 393294 610954 393914 646398
rect 393294 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 393914 610954
rect 393294 610634 393914 610718
rect 393294 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 393914 610634
rect 393294 574954 393914 610398
rect 393294 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 393914 574954
rect 393294 574634 393914 574718
rect 393294 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 393914 574634
rect 393294 538954 393914 574398
rect 393294 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 393914 538954
rect 393294 538634 393914 538718
rect 393294 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 393914 538634
rect 393294 502954 393914 538398
rect 393294 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 393914 502954
rect 393294 502634 393914 502718
rect 393294 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 393914 502634
rect 393294 466954 393914 502398
rect 393294 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 393914 466954
rect 393294 466634 393914 466718
rect 393294 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 393914 466634
rect 393294 430954 393914 466398
rect 393294 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 393914 430954
rect 393294 430634 393914 430718
rect 393294 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 393914 430634
rect 393294 394954 393914 430398
rect 393294 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 393914 394954
rect 393294 394634 393914 394718
rect 393294 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 393914 394634
rect 393294 358954 393914 394398
rect 393294 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 393914 358954
rect 393294 358634 393914 358718
rect 393294 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 393914 358634
rect 393294 322954 393914 358398
rect 393294 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 393914 322954
rect 393294 322634 393914 322718
rect 393294 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 393914 322634
rect 393294 286954 393914 322398
rect 393294 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 393914 286954
rect 393294 286634 393914 286718
rect 393294 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 393914 286634
rect 393294 250954 393914 286398
rect 393294 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 393914 250954
rect 393294 250634 393914 250718
rect 393294 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 393914 250634
rect 393294 248684 393914 250398
rect 65300 246303 70100 246486
rect 65300 246067 65342 246303
rect 65578 246067 65662 246303
rect 65898 246067 65982 246303
rect 66218 246067 66302 246303
rect 66538 246067 66622 246303
rect 66858 246067 66942 246303
rect 67178 246067 67262 246303
rect 67498 246067 67582 246303
rect 67818 246067 67902 246303
rect 68138 246067 68222 246303
rect 68458 246067 68542 246303
rect 68778 246067 68862 246303
rect 69098 246067 69182 246303
rect 69418 246067 69502 246303
rect 69738 246067 69822 246303
rect 70058 246067 70100 246303
rect 65300 245884 70100 246067
rect 65300 241953 71300 241984
rect 65300 241717 65462 241953
rect 65698 241717 65782 241953
rect 66018 241717 66102 241953
rect 66338 241717 66422 241953
rect 66658 241717 66742 241953
rect 66978 241717 67062 241953
rect 67298 241717 67382 241953
rect 67618 241717 67702 241953
rect 67938 241717 68022 241953
rect 68258 241717 68342 241953
rect 68578 241717 68662 241953
rect 68898 241717 68982 241953
rect 69218 241717 69302 241953
rect 69538 241717 69622 241953
rect 69858 241717 69942 241953
rect 70178 241717 70262 241953
rect 70498 241717 70582 241953
rect 70818 241717 70902 241953
rect 71138 241717 71300 241953
rect 65300 241633 71300 241717
rect 65300 241397 65462 241633
rect 65698 241397 65782 241633
rect 66018 241397 66102 241633
rect 66338 241397 66422 241633
rect 66658 241397 66742 241633
rect 66978 241397 67062 241633
rect 67298 241397 67382 241633
rect 67618 241397 67702 241633
rect 67938 241397 68022 241633
rect 68258 241397 68342 241633
rect 68578 241397 68662 241633
rect 68898 241397 68982 241633
rect 69218 241397 69302 241633
rect 69538 241397 69622 241633
rect 69858 241397 69942 241633
rect 70178 241397 70262 241633
rect 70498 241397 70582 241633
rect 70818 241397 70902 241633
rect 71138 241397 71300 241633
rect 65300 241366 71300 241397
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42294 151954 42914 187398
rect 42294 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 42914 151954
rect 42294 151634 42914 151718
rect 42294 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 42914 151634
rect 42294 115954 42914 151398
rect 42294 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 42914 115954
rect 42294 115634 42914 115718
rect 42294 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 42914 115634
rect 42294 79954 42914 115398
rect 42294 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 42914 79954
rect 42294 79634 42914 79718
rect 42294 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 42914 79634
rect 42294 43954 42914 79398
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1306 42914 7398
rect 42294 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 42914 -1306
rect 42294 -1626 42914 -1542
rect 42294 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 42914 -1626
rect 42294 -7654 42914 -1862
rect 46794 228453 47414 228484
rect 46794 228217 46826 228453
rect 47062 228217 47146 228453
rect 47382 228217 47414 228453
rect 46794 228133 47414 228217
rect 46794 227897 46826 228133
rect 47062 227897 47146 228133
rect 47382 227897 47414 228133
rect 46794 192454 47414 227897
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46794 120454 47414 155898
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 84454 47414 119898
rect 46794 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 47414 84454
rect 46794 84134 47414 84218
rect 46794 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 47414 84134
rect 46794 48454 47414 83898
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2266 47414 11898
rect 46794 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 47414 -2266
rect 46794 -2586 47414 -2502
rect 46794 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 47414 -2586
rect 46794 -7654 47414 -2822
rect 51294 196954 51914 228484
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 51294 160954 51914 196398
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 124954 51914 160398
rect 51294 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 51914 124954
rect 51294 124634 51914 124718
rect 51294 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 51914 124634
rect 51294 88954 51914 124398
rect 51294 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 51914 88954
rect 51294 88634 51914 88718
rect 51294 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 51914 88634
rect 51294 52954 51914 88398
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3226 51914 16398
rect 51294 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 51914 -3226
rect 51294 -3546 51914 -3462
rect 51294 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 51914 -3546
rect 51294 -7654 51914 -3782
rect 55794 201454 56414 228484
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4186 56414 20898
rect 55794 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 56414 -4186
rect 55794 -4506 56414 -4422
rect 55794 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 56414 -4506
rect 55794 -7654 56414 -4742
rect 60294 205954 60914 228484
rect 60294 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 60914 205954
rect 60294 205634 60914 205718
rect 60294 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 60914 205634
rect 60294 169954 60914 205398
rect 60294 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 60914 169954
rect 60294 169634 60914 169718
rect 60294 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 60914 169634
rect 60294 133954 60914 169398
rect 60294 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 60914 133954
rect 60294 133634 60914 133718
rect 60294 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 60914 133634
rect 60294 97954 60914 133398
rect 60294 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 60914 97954
rect 60294 97634 60914 97718
rect 60294 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 60914 97634
rect 60294 61954 60914 97398
rect 60294 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 60914 61954
rect 60294 61634 60914 61718
rect 60294 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 60914 61634
rect 60294 25954 60914 61398
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 60294 -5146 60914 25398
rect 60294 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 60914 -5146
rect 60294 -5466 60914 -5382
rect 60294 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 60914 -5466
rect 60294 -7654 60914 -5702
rect 64794 210454 65414 228484
rect 64794 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 65414 210454
rect 64794 210134 65414 210218
rect 64794 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 65414 210134
rect 64794 174454 65414 209898
rect 64794 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 65414 174454
rect 64794 174134 65414 174218
rect 64794 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 65414 174134
rect 64794 138454 65414 173898
rect 64794 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 65414 138454
rect 64794 138134 65414 138218
rect 64794 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 65414 138134
rect 64794 102454 65414 137898
rect 64794 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 65414 102454
rect 64794 102134 65414 102218
rect 64794 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 65414 102134
rect 64794 66454 65414 101898
rect 64794 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 65414 66454
rect 64794 66134 65414 66218
rect 64794 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 65414 66134
rect 64794 30454 65414 65898
rect 64794 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 65414 30454
rect 64794 30134 65414 30218
rect 64794 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 65414 30134
rect 64794 -6106 65414 29898
rect 64794 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 65414 -6106
rect 64794 -6426 65414 -6342
rect 64794 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 65414 -6426
rect 64794 -7654 65414 -6662
rect 69294 214954 69914 228484
rect 69294 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 69914 214954
rect 69294 214634 69914 214718
rect 69294 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 69914 214634
rect 69294 178954 69914 214398
rect 69294 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 69914 178954
rect 69294 178634 69914 178718
rect 69294 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 69914 178634
rect 69294 142954 69914 178398
rect 69294 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 69914 142954
rect 69294 142634 69914 142718
rect 69294 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 69914 142634
rect 69294 106954 69914 142398
rect 69294 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 69914 106954
rect 69294 106634 69914 106718
rect 69294 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 69914 106634
rect 69294 70954 69914 106398
rect 69294 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 69914 70954
rect 69294 70634 69914 70718
rect 69294 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 69914 70634
rect 69294 34954 69914 70398
rect 69294 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 69914 34954
rect 69294 34634 69914 34718
rect 69294 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 69914 34634
rect 69294 -7066 69914 34398
rect 69294 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 69914 -7066
rect 69294 -7386 69914 -7302
rect 69294 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 69914 -7386
rect 69294 -7654 69914 -7622
rect 73794 219454 74414 228484
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 78294 223954 78914 228484
rect 78294 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 78914 223954
rect 78294 223634 78914 223718
rect 78294 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 78914 223634
rect 78294 187954 78914 223398
rect 78294 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 78914 187954
rect 78294 187634 78914 187718
rect 78294 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 78914 187634
rect 78294 151954 78914 187398
rect 78294 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 78914 151954
rect 78294 151634 78914 151718
rect 78294 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 78914 151634
rect 78294 115954 78914 151398
rect 78294 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 78914 115954
rect 78294 115634 78914 115718
rect 78294 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 78914 115634
rect 78294 79954 78914 115398
rect 78294 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 78914 79954
rect 78294 79634 78914 79718
rect 78294 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 78914 79634
rect 78294 43954 78914 79398
rect 78294 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 78914 43954
rect 78294 43634 78914 43718
rect 78294 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 78914 43634
rect 78294 7954 78914 43398
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1306 78914 7398
rect 78294 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 78914 -1306
rect 78294 -1626 78914 -1542
rect 78294 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 78914 -1626
rect 78294 -7654 78914 -1862
rect 82794 228453 83414 228484
rect 82794 228217 82826 228453
rect 83062 228217 83146 228453
rect 83382 228217 83414 228453
rect 82794 228133 83414 228217
rect 82794 227897 82826 228133
rect 83062 227897 83146 228133
rect 83382 227897 83414 228133
rect 82794 192454 83414 227897
rect 82794 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 83414 192454
rect 82794 192134 83414 192218
rect 82794 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 83414 192134
rect 82794 156454 83414 191898
rect 82794 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 83414 156454
rect 82794 156134 83414 156218
rect 82794 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 83414 156134
rect 82794 120454 83414 155898
rect 82794 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 83414 120454
rect 82794 120134 83414 120218
rect 82794 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 83414 120134
rect 82794 84454 83414 119898
rect 82794 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 83414 84454
rect 82794 84134 83414 84218
rect 82794 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 83414 84134
rect 82794 48454 83414 83898
rect 82794 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 83414 48454
rect 82794 48134 83414 48218
rect 82794 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 83414 48134
rect 82794 12454 83414 47898
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2266 83414 11898
rect 82794 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 83414 -2266
rect 82794 -2586 83414 -2502
rect 82794 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 83414 -2586
rect 82794 -7654 83414 -2822
rect 87294 196954 87914 228484
rect 87294 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 87914 196954
rect 87294 196634 87914 196718
rect 87294 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 87914 196634
rect 87294 160954 87914 196398
rect 87294 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 87914 160954
rect 87294 160634 87914 160718
rect 87294 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 87914 160634
rect 87294 124954 87914 160398
rect 87294 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 87914 124954
rect 87294 124634 87914 124718
rect 87294 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 87914 124634
rect 87294 88954 87914 124398
rect 87294 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 87914 88954
rect 87294 88634 87914 88718
rect 87294 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 87914 88634
rect 87294 52954 87914 88398
rect 87294 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 87914 52954
rect 87294 52634 87914 52718
rect 87294 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 87914 52634
rect 87294 16954 87914 52398
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3226 87914 16398
rect 87294 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 87914 -3226
rect 87294 -3546 87914 -3462
rect 87294 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 87914 -3546
rect 87294 -7654 87914 -3782
rect 91794 201454 92414 228484
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4186 92414 20898
rect 91794 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 92414 -4186
rect 91794 -4506 92414 -4422
rect 91794 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 92414 -4506
rect 91794 -7654 92414 -4742
rect 96294 205954 96914 228484
rect 96294 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 96914 205954
rect 96294 205634 96914 205718
rect 96294 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 96914 205634
rect 96294 169954 96914 205398
rect 96294 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 96914 169954
rect 96294 169634 96914 169718
rect 96294 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 96914 169634
rect 96294 133954 96914 169398
rect 96294 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 96914 133954
rect 96294 133634 96914 133718
rect 96294 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 96914 133634
rect 96294 97954 96914 133398
rect 96294 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 96914 97954
rect 96294 97634 96914 97718
rect 96294 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 96914 97634
rect 96294 61954 96914 97398
rect 96294 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 96914 61954
rect 96294 61634 96914 61718
rect 96294 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 96914 61634
rect 96294 25954 96914 61398
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96294 -5146 96914 25398
rect 96294 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 96914 -5146
rect 96294 -5466 96914 -5382
rect 96294 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 96914 -5466
rect 96294 -7654 96914 -5702
rect 100794 210454 101414 228484
rect 100794 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 101414 210454
rect 100794 210134 101414 210218
rect 100794 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 101414 210134
rect 100794 174454 101414 209898
rect 100794 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 101414 174454
rect 100794 174134 101414 174218
rect 100794 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 101414 174134
rect 100794 138454 101414 173898
rect 100794 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 101414 138454
rect 100794 138134 101414 138218
rect 100794 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 101414 138134
rect 100794 102454 101414 137898
rect 100794 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 101414 102454
rect 100794 102134 101414 102218
rect 100794 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 101414 102134
rect 100794 66454 101414 101898
rect 100794 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 101414 66454
rect 100794 66134 101414 66218
rect 100794 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 101414 66134
rect 100794 30454 101414 65898
rect 100794 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 101414 30454
rect 100794 30134 101414 30218
rect 100794 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 101414 30134
rect 100794 -6106 101414 29898
rect 100794 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 101414 -6106
rect 100794 -6426 101414 -6342
rect 100794 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 101414 -6426
rect 100794 -7654 101414 -6662
rect 105294 214954 105914 228484
rect 105294 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 105914 214954
rect 105294 214634 105914 214718
rect 105294 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 105914 214634
rect 105294 178954 105914 214398
rect 105294 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 105914 178954
rect 105294 178634 105914 178718
rect 105294 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 105914 178634
rect 105294 142954 105914 178398
rect 105294 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 105914 142954
rect 105294 142634 105914 142718
rect 105294 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 105914 142634
rect 105294 106954 105914 142398
rect 105294 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 105914 106954
rect 105294 106634 105914 106718
rect 105294 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 105914 106634
rect 105294 70954 105914 106398
rect 105294 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 105914 70954
rect 105294 70634 105914 70718
rect 105294 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 105914 70634
rect 105294 34954 105914 70398
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 105294 -7066 105914 34398
rect 105294 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 105914 -7066
rect 105294 -7386 105914 -7302
rect 105294 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 105914 -7386
rect 105294 -7654 105914 -7622
rect 109794 219454 110414 228484
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 114294 223954 114914 228484
rect 114294 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 114914 223954
rect 114294 223634 114914 223718
rect 114294 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 114914 223634
rect 114294 187954 114914 223398
rect 114294 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 114914 187954
rect 114294 187634 114914 187718
rect 114294 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 114914 187634
rect 114294 151954 114914 187398
rect 114294 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 114914 151954
rect 114294 151634 114914 151718
rect 114294 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 114914 151634
rect 114294 115954 114914 151398
rect 118794 228453 119414 228484
rect 118794 228217 118826 228453
rect 119062 228217 119146 228453
rect 119382 228217 119414 228453
rect 118794 228133 119414 228217
rect 118794 227897 118826 228133
rect 119062 227897 119146 228133
rect 119382 227897 119414 228133
rect 118794 192454 119414 227897
rect 118794 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 119414 192454
rect 118794 192134 119414 192218
rect 118794 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 119414 192134
rect 118794 156454 119414 191898
rect 118794 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 119414 156454
rect 118794 156134 119414 156218
rect 118794 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 119414 156134
rect 118794 142000 119414 155898
rect 123294 196954 123914 228484
rect 123294 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 123914 196954
rect 123294 196634 123914 196718
rect 123294 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 123914 196634
rect 123294 160954 123914 196398
rect 123294 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 123914 160954
rect 123294 160634 123914 160718
rect 123294 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 123914 160634
rect 123294 142000 123914 160398
rect 127794 201454 128414 228484
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 142000 128414 164898
rect 132294 205954 132914 228484
rect 172794 210454 173414 228484
rect 172794 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 173414 210454
rect 172794 210134 173414 210218
rect 172794 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 173414 210134
rect 132294 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 132914 205954
rect 132294 205634 132914 205718
rect 132294 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 132914 205634
rect 135914 205861 165514 205986
rect 135914 205625 136036 205861
rect 136272 205625 136356 205861
rect 136592 205625 136676 205861
rect 136912 205625 136996 205861
rect 137232 205625 137316 205861
rect 137552 205625 137636 205861
rect 137872 205625 137956 205861
rect 138192 205625 138276 205861
rect 138512 205625 138596 205861
rect 138832 205625 138916 205861
rect 139152 205625 139236 205861
rect 139472 205625 139556 205861
rect 139792 205625 139876 205861
rect 140112 205625 140196 205861
rect 140432 205625 140516 205861
rect 140752 205625 140836 205861
rect 141072 205625 141156 205861
rect 141392 205625 141476 205861
rect 141712 205625 141796 205861
rect 142032 205625 142116 205861
rect 142352 205625 142436 205861
rect 142672 205625 142756 205861
rect 142992 205625 143076 205861
rect 143312 205625 143396 205861
rect 143632 205625 143716 205861
rect 143952 205625 144036 205861
rect 144272 205625 144356 205861
rect 144592 205625 144676 205861
rect 144912 205625 144996 205861
rect 145232 205625 145316 205861
rect 145552 205625 145636 205861
rect 145872 205625 145956 205861
rect 146192 205625 146276 205861
rect 146512 205625 146596 205861
rect 146832 205625 146916 205861
rect 147152 205625 147236 205861
rect 147472 205625 147556 205861
rect 147792 205625 147876 205861
rect 148112 205625 148196 205861
rect 148432 205625 148516 205861
rect 148752 205625 148836 205861
rect 149072 205625 149156 205861
rect 149392 205625 149476 205861
rect 149712 205625 149796 205861
rect 150032 205625 150116 205861
rect 150352 205625 150436 205861
rect 150672 205625 150756 205861
rect 150992 205625 151076 205861
rect 151312 205625 151396 205861
rect 151632 205625 151716 205861
rect 151952 205625 152036 205861
rect 152272 205625 152356 205861
rect 152592 205625 152676 205861
rect 152912 205625 152996 205861
rect 153232 205625 153316 205861
rect 153552 205625 153636 205861
rect 153872 205625 153956 205861
rect 154192 205625 154276 205861
rect 154512 205625 154596 205861
rect 154832 205625 154916 205861
rect 155152 205625 155236 205861
rect 155472 205625 155556 205861
rect 155792 205625 155876 205861
rect 156112 205625 156196 205861
rect 156432 205625 156516 205861
rect 156752 205625 156836 205861
rect 157072 205625 157156 205861
rect 157392 205625 157476 205861
rect 157712 205625 157796 205861
rect 158032 205625 158116 205861
rect 158352 205625 158436 205861
rect 158672 205625 158756 205861
rect 158992 205625 159076 205861
rect 159312 205625 159396 205861
rect 159632 205625 159716 205861
rect 159952 205625 160036 205861
rect 160272 205625 160356 205861
rect 160592 205625 160676 205861
rect 160912 205625 160996 205861
rect 161232 205625 161316 205861
rect 161552 205625 161636 205861
rect 161872 205625 161956 205861
rect 162192 205625 162276 205861
rect 162512 205625 162596 205861
rect 162832 205625 162916 205861
rect 163152 205625 163236 205861
rect 163472 205625 163556 205861
rect 163792 205625 163876 205861
rect 164112 205625 164196 205861
rect 164432 205625 164516 205861
rect 164752 205625 164836 205861
rect 165072 205625 165156 205861
rect 165392 205625 165514 205861
rect 135914 205500 165514 205625
rect 132294 169954 132914 205398
rect 137314 201411 165514 201486
rect 137314 201175 137376 201411
rect 137612 201175 137696 201411
rect 137932 201175 138016 201411
rect 138252 201175 138336 201411
rect 138572 201175 138656 201411
rect 138892 201175 138976 201411
rect 139212 201175 139296 201411
rect 139532 201175 139616 201411
rect 139852 201175 139936 201411
rect 140172 201175 140256 201411
rect 140492 201175 140576 201411
rect 140812 201175 140896 201411
rect 141132 201175 141216 201411
rect 141452 201175 141536 201411
rect 141772 201175 141856 201411
rect 142092 201175 142176 201411
rect 142412 201175 142496 201411
rect 142732 201175 142816 201411
rect 143052 201175 143136 201411
rect 143372 201175 143456 201411
rect 143692 201175 143776 201411
rect 144012 201175 144096 201411
rect 144332 201175 144416 201411
rect 144652 201175 144736 201411
rect 144972 201175 145056 201411
rect 145292 201175 145376 201411
rect 145612 201175 145696 201411
rect 145932 201175 146016 201411
rect 146252 201175 146336 201411
rect 146572 201175 146656 201411
rect 146892 201175 146976 201411
rect 147212 201175 147296 201411
rect 147532 201175 147616 201411
rect 147852 201175 147936 201411
rect 148172 201175 148256 201411
rect 148492 201175 148576 201411
rect 148812 201175 148896 201411
rect 149132 201175 149216 201411
rect 149452 201175 149536 201411
rect 149772 201175 149856 201411
rect 150092 201175 150176 201411
rect 150412 201175 150496 201411
rect 150732 201175 150816 201411
rect 151052 201175 151136 201411
rect 151372 201175 151456 201411
rect 151692 201175 151776 201411
rect 152012 201175 152096 201411
rect 152332 201175 152416 201411
rect 152652 201175 152736 201411
rect 152972 201175 153056 201411
rect 153292 201175 153376 201411
rect 153612 201175 153696 201411
rect 153932 201175 154016 201411
rect 154252 201175 154336 201411
rect 154572 201175 154656 201411
rect 154892 201175 154976 201411
rect 155212 201175 155296 201411
rect 155532 201175 155616 201411
rect 155852 201175 155936 201411
rect 156172 201175 156256 201411
rect 156492 201175 156576 201411
rect 156812 201175 156896 201411
rect 157132 201175 157216 201411
rect 157452 201175 157536 201411
rect 157772 201175 157856 201411
rect 158092 201175 158176 201411
rect 158412 201175 158496 201411
rect 158732 201175 158816 201411
rect 159052 201175 159136 201411
rect 159372 201175 159456 201411
rect 159692 201175 159776 201411
rect 160012 201175 160096 201411
rect 160332 201175 160416 201411
rect 160652 201175 160736 201411
rect 160972 201175 161056 201411
rect 161292 201175 161376 201411
rect 161612 201175 161696 201411
rect 161932 201175 162016 201411
rect 162252 201175 162336 201411
rect 162572 201175 162656 201411
rect 162892 201175 162976 201411
rect 163212 201175 163296 201411
rect 163532 201175 163616 201411
rect 163852 201175 163936 201411
rect 164172 201175 164256 201411
rect 164492 201175 164576 201411
rect 164812 201175 164896 201411
rect 165132 201175 165216 201411
rect 165452 201175 165514 201411
rect 137314 201100 165514 201175
rect 144499 191044 144565 191045
rect 144499 190980 144500 191044
rect 144564 190980 144565 191044
rect 144499 190979 144565 190980
rect 144502 186013 144562 190979
rect 146155 188596 146221 188597
rect 146155 188532 146156 188596
rect 146220 188532 146221 188596
rect 146155 188531 146221 188532
rect 144499 186012 144565 186013
rect 144499 185948 144500 186012
rect 144564 185948 144565 186012
rect 144499 185947 144565 185948
rect 142843 184380 142909 184381
rect 142843 184316 142844 184380
rect 142908 184316 142909 184380
rect 142843 184315 142909 184316
rect 141003 184244 141069 184245
rect 141003 184180 141004 184244
rect 141068 184180 141069 184244
rect 141003 184179 141069 184180
rect 141006 178805 141066 184179
rect 142475 181116 142541 181117
rect 142475 181052 142476 181116
rect 142540 181052 142541 181116
rect 142475 181051 142541 181052
rect 141003 178804 141069 178805
rect 141003 178740 141004 178804
rect 141068 178740 141069 178804
rect 141003 178739 141069 178740
rect 137014 174454 141514 174486
rect 137014 174218 137066 174454
rect 137302 174218 137386 174454
rect 137622 174218 137706 174454
rect 137942 174218 138026 174454
rect 138262 174218 138346 174454
rect 138582 174218 138666 174454
rect 138902 174218 138986 174454
rect 139222 174218 139306 174454
rect 139542 174218 139626 174454
rect 139862 174218 139946 174454
rect 140182 174218 140266 174454
rect 140502 174218 140586 174454
rect 140822 174218 140906 174454
rect 141142 174218 141226 174454
rect 141462 174218 141514 174454
rect 137014 174134 141514 174218
rect 137014 173898 137066 174134
rect 137302 173898 137386 174134
rect 137622 173898 137706 174134
rect 137942 173898 138026 174134
rect 138262 173898 138346 174134
rect 138582 173898 138666 174134
rect 138902 173898 138986 174134
rect 139222 173898 139306 174134
rect 139542 173898 139626 174134
rect 139862 173898 139946 174134
rect 140182 173898 140266 174134
rect 140502 173898 140586 174134
rect 140822 173898 140906 174134
rect 141142 173898 141226 174134
rect 141462 173898 141514 174134
rect 137014 173866 141514 173898
rect 142478 172957 142538 181051
rect 142846 178805 142906 184315
rect 143027 184108 143093 184109
rect 143027 184044 143028 184108
rect 143092 184044 143093 184108
rect 143027 184043 143093 184044
rect 143030 178941 143090 184043
rect 143027 178940 143093 178941
rect 143027 178876 143028 178940
rect 143092 178876 143093 178940
rect 143027 178875 143093 178876
rect 142843 178804 142909 178805
rect 142843 178740 142844 178804
rect 142908 178740 142909 178804
rect 142843 178739 142909 178740
rect 142475 172956 142541 172957
rect 142475 172892 142476 172956
rect 142540 172892 142541 172956
rect 142475 172891 142541 172892
rect 132294 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 132914 169954
rect 132294 169634 132914 169718
rect 132294 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 132914 169634
rect 132294 142000 132914 169398
rect 146158 142765 146218 188531
rect 146339 186012 146405 186013
rect 146339 185948 146340 186012
rect 146404 185948 146405 186012
rect 146339 185947 146405 185948
rect 146342 175405 146402 185947
rect 158483 176492 158549 176493
rect 158483 176428 158484 176492
rect 158548 176428 158549 176492
rect 158483 176427 158549 176428
rect 146339 175404 146405 175405
rect 146339 175340 146340 175404
rect 146404 175340 146405 175404
rect 146339 175339 146405 175340
rect 158486 172957 158546 176427
rect 172794 174454 173414 209898
rect 172794 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 173414 174454
rect 172794 174134 173414 174218
rect 172794 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 173414 174134
rect 158483 172956 158549 172957
rect 158483 172892 158484 172956
rect 158548 172892 158549 172956
rect 158483 172891 158549 172892
rect 146155 142764 146221 142765
rect 146155 142700 146156 142764
rect 146220 142700 146221 142764
rect 146155 142699 146221 142700
rect 172794 142000 173414 173898
rect 177294 214954 177914 228484
rect 177294 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 177914 214954
rect 177294 214634 177914 214718
rect 177294 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 177914 214634
rect 177294 178954 177914 214398
rect 177294 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 177914 178954
rect 177294 178634 177914 178718
rect 177294 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 177914 178634
rect 177294 142954 177914 178398
rect 177294 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 177914 142954
rect 177294 142634 177914 142718
rect 177294 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 177914 142634
rect 177294 142000 177914 142398
rect 181794 219454 182414 228484
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 142000 182414 146898
rect 186294 223954 186914 228484
rect 186294 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 186914 223954
rect 186294 223634 186914 223718
rect 186294 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 186914 223634
rect 186294 187954 186914 223398
rect 186294 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 186914 187954
rect 186294 187634 186914 187718
rect 186294 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 186914 187634
rect 186294 151954 186914 187398
rect 186294 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 186914 151954
rect 186294 151634 186914 151718
rect 186294 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 186914 151634
rect 114294 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 114914 115954
rect 114294 115634 114914 115718
rect 114294 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 114914 115634
rect 114294 79954 114914 115398
rect 139568 115954 139888 115986
rect 139568 115718 139610 115954
rect 139846 115718 139888 115954
rect 139568 115634 139888 115718
rect 139568 115398 139610 115634
rect 139846 115398 139888 115634
rect 139568 115366 139888 115398
rect 170288 115954 170608 115986
rect 170288 115718 170330 115954
rect 170566 115718 170608 115954
rect 170288 115634 170608 115718
rect 170288 115398 170330 115634
rect 170566 115398 170608 115634
rect 170288 115366 170608 115398
rect 186294 115954 186914 151398
rect 186294 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 186914 115954
rect 186294 115634 186914 115718
rect 186294 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 186914 115634
rect 124208 111454 124528 111486
rect 124208 111218 124250 111454
rect 124486 111218 124528 111454
rect 124208 111134 124528 111218
rect 124208 110898 124250 111134
rect 124486 110898 124528 111134
rect 124208 110866 124528 110898
rect 154928 111454 155248 111486
rect 154928 111218 154970 111454
rect 155206 111218 155248 111454
rect 154928 111134 155248 111218
rect 154928 110898 154970 111134
rect 155206 110898 155248 111134
rect 154928 110866 155248 110898
rect 173571 81292 173637 81293
rect 173571 81228 173572 81292
rect 173636 81228 173637 81292
rect 173571 81227 173637 81228
rect 171547 81156 171613 81157
rect 171547 81092 171548 81156
rect 171612 81092 171613 81156
rect 171547 81091 171613 81092
rect 171179 80748 171245 80749
rect 171179 80684 171180 80748
rect 171244 80684 171245 80748
rect 171179 80683 171245 80684
rect 166211 80612 166277 80613
rect 166211 80548 166212 80612
rect 166276 80548 166277 80612
rect 166211 80547 166277 80548
rect 166214 80205 166274 80547
rect 131803 80204 131869 80205
rect 131803 80140 131804 80204
rect 131868 80140 131869 80204
rect 131803 80139 131869 80140
rect 142843 80204 142909 80205
rect 142843 80140 142844 80204
rect 142908 80140 142909 80204
rect 142843 80139 142909 80140
rect 159219 80204 159285 80205
rect 159219 80140 159220 80204
rect 159284 80140 159285 80204
rect 159219 80139 159285 80140
rect 166211 80204 166277 80205
rect 166211 80140 166212 80204
rect 166276 80140 166277 80204
rect 166211 80139 166277 80140
rect 114294 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 114914 79954
rect 125731 79932 125797 79933
rect 125731 79868 125732 79932
rect 125796 79868 125797 79932
rect 125731 79867 125797 79868
rect 125915 79932 125981 79933
rect 125915 79868 125916 79932
rect 125980 79868 125981 79932
rect 125915 79867 125981 79868
rect 128491 79932 128557 79933
rect 128491 79868 128492 79932
rect 128556 79868 128557 79932
rect 128491 79867 128557 79868
rect 129043 79932 129109 79933
rect 129043 79868 129044 79932
rect 129108 79868 129109 79932
rect 129043 79867 129109 79868
rect 129963 79932 130029 79933
rect 129963 79868 129964 79932
rect 130028 79868 130029 79932
rect 129963 79867 130029 79868
rect 131619 79932 131685 79933
rect 131619 79868 131620 79932
rect 131684 79868 131685 79932
rect 131619 79867 131685 79868
rect 114294 79634 114914 79718
rect 114294 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 114914 79634
rect 114294 43954 114914 79398
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114294 7954 114914 43398
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1306 114914 7398
rect 114294 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 114914 -1306
rect 114294 -1626 114914 -1542
rect 114294 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 114914 -1626
rect 114294 -7654 114914 -1862
rect 118794 48454 119414 78000
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 118794 12454 119414 47898
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2266 119414 11898
rect 118794 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 119414 -2266
rect 118794 -2586 119414 -2502
rect 118794 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 119414 -2586
rect 118794 -7654 119414 -2822
rect 123294 52954 123914 78000
rect 125734 75173 125794 79867
rect 125918 78845 125978 79867
rect 127387 79660 127453 79661
rect 127387 79596 127388 79660
rect 127452 79596 127453 79660
rect 127387 79595 127453 79596
rect 125915 78844 125981 78845
rect 125915 78780 125916 78844
rect 125980 78780 125981 78844
rect 125915 78779 125981 78780
rect 125915 78708 125981 78709
rect 125915 78644 125916 78708
rect 125980 78644 125981 78708
rect 125915 78643 125981 78644
rect 125731 75172 125797 75173
rect 125731 75108 125732 75172
rect 125796 75108 125797 75172
rect 125731 75107 125797 75108
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3226 123914 16398
rect 125918 4861 125978 78643
rect 127390 77621 127450 79595
rect 127387 77620 127453 77621
rect 127387 77556 127388 77620
rect 127452 77556 127453 77620
rect 127387 77555 127453 77556
rect 127387 77484 127453 77485
rect 127387 77420 127388 77484
rect 127452 77420 127453 77484
rect 127387 77419 127453 77420
rect 127203 77348 127269 77349
rect 127203 77284 127204 77348
rect 127268 77284 127269 77348
rect 127203 77283 127269 77284
rect 127206 43485 127266 77283
rect 127203 43484 127269 43485
rect 127203 43420 127204 43484
rect 127268 43420 127269 43484
rect 127203 43419 127269 43420
rect 125915 4860 125981 4861
rect 125915 4796 125916 4860
rect 125980 4796 125981 4860
rect 125915 4795 125981 4796
rect 127390 3365 127450 77419
rect 127794 57454 128414 78000
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127387 3364 127453 3365
rect 127387 3300 127388 3364
rect 127452 3300 127453 3364
rect 127387 3299 127453 3300
rect 123294 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 123914 -3226
rect 123294 -3546 123914 -3462
rect 123294 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 123914 -3546
rect 123294 -7654 123914 -3782
rect 127794 -4186 128414 20898
rect 128494 7850 128554 79867
rect 128859 79660 128925 79661
rect 128859 79596 128860 79660
rect 128924 79596 128925 79660
rect 128859 79595 128925 79596
rect 128675 78844 128741 78845
rect 128675 78780 128676 78844
rect 128740 78780 128741 78844
rect 128675 78779 128741 78780
rect 128678 16590 128738 78779
rect 128862 73813 128922 79595
rect 129046 78573 129106 79867
rect 129779 79660 129845 79661
rect 129779 79596 129780 79660
rect 129844 79596 129845 79660
rect 129779 79595 129845 79596
rect 129043 78572 129109 78573
rect 129043 78508 129044 78572
rect 129108 78508 129109 78572
rect 129043 78507 129109 78508
rect 129782 75445 129842 79595
rect 129779 75444 129845 75445
rect 129779 75380 129780 75444
rect 129844 75380 129845 75444
rect 129779 75379 129845 75380
rect 128859 73812 128925 73813
rect 128859 73748 128860 73812
rect 128924 73748 128925 73812
rect 128859 73747 128925 73748
rect 128678 16530 128922 16590
rect 128494 7790 128738 7850
rect 128678 7717 128738 7790
rect 128675 7716 128741 7717
rect 128675 7652 128676 7716
rect 128740 7652 128741 7716
rect 128675 7651 128741 7652
rect 128862 7581 128922 16530
rect 129966 8941 130026 79867
rect 130883 79796 130949 79797
rect 130883 79732 130884 79796
rect 130948 79732 130949 79796
rect 130883 79731 130949 79732
rect 130331 78844 130397 78845
rect 130331 78780 130332 78844
rect 130396 78780 130397 78844
rect 130331 78779 130397 78780
rect 130147 78708 130213 78709
rect 130147 78644 130148 78708
rect 130212 78644 130213 78708
rect 130147 78643 130213 78644
rect 129963 8940 130029 8941
rect 129963 8876 129964 8940
rect 130028 8876 130029 8940
rect 129963 8875 130029 8876
rect 130150 7853 130210 78643
rect 130334 75581 130394 78779
rect 130886 78573 130946 79731
rect 131622 78845 131682 79867
rect 131619 78844 131685 78845
rect 131619 78780 131620 78844
rect 131684 78780 131685 78844
rect 131619 78779 131685 78780
rect 130883 78572 130949 78573
rect 130883 78508 130884 78572
rect 130948 78508 130949 78572
rect 130883 78507 130949 78508
rect 131435 78436 131501 78437
rect 131435 78372 131436 78436
rect 131500 78372 131501 78436
rect 131435 78371 131501 78372
rect 131251 77076 131317 77077
rect 131251 77012 131252 77076
rect 131316 77012 131317 77076
rect 131251 77011 131317 77012
rect 130331 75580 130397 75581
rect 130331 75516 130332 75580
rect 130396 75516 130397 75580
rect 130331 75515 130397 75516
rect 131067 73268 131133 73269
rect 131067 73204 131068 73268
rect 131132 73204 131133 73268
rect 131067 73203 131133 73204
rect 130147 7852 130213 7853
rect 130147 7788 130148 7852
rect 130212 7788 130213 7852
rect 130147 7787 130213 7788
rect 128859 7580 128925 7581
rect 128859 7516 128860 7580
rect 128924 7516 128925 7580
rect 128859 7515 128925 7516
rect 131070 3501 131130 73203
rect 131254 6221 131314 77011
rect 131438 9077 131498 78371
rect 131806 76805 131866 80139
rect 133459 79932 133525 79933
rect 133459 79868 133460 79932
rect 133524 79868 133525 79932
rect 133459 79867 133525 79868
rect 134011 79932 134077 79933
rect 134011 79868 134012 79932
rect 134076 79868 134077 79932
rect 134011 79867 134077 79868
rect 134563 79932 134629 79933
rect 134563 79868 134564 79932
rect 134628 79868 134629 79932
rect 134563 79867 134629 79868
rect 135483 79932 135549 79933
rect 135483 79868 135484 79932
rect 135548 79868 135549 79932
rect 135483 79867 135549 79868
rect 136403 79932 136469 79933
rect 136403 79868 136404 79932
rect 136468 79868 136469 79932
rect 136403 79867 136469 79868
rect 136955 79932 137021 79933
rect 136955 79868 136956 79932
rect 137020 79868 137021 79932
rect 136955 79867 137021 79868
rect 138059 79932 138125 79933
rect 138059 79868 138060 79932
rect 138124 79868 138125 79932
rect 138059 79867 138125 79868
rect 140267 79932 140333 79933
rect 140267 79868 140268 79932
rect 140332 79868 140333 79932
rect 140267 79867 140333 79868
rect 133091 79796 133157 79797
rect 133091 79732 133092 79796
rect 133156 79732 133157 79796
rect 133091 79731 133157 79732
rect 133275 79796 133341 79797
rect 133275 79732 133276 79796
rect 133340 79732 133341 79796
rect 133275 79731 133341 79732
rect 131987 77756 132053 77757
rect 131987 77692 131988 77756
rect 132052 77692 132053 77756
rect 131987 77691 132053 77692
rect 131803 76804 131869 76805
rect 131803 76740 131804 76804
rect 131868 76740 131869 76804
rect 131803 76739 131869 76740
rect 131435 9076 131501 9077
rect 131435 9012 131436 9076
rect 131500 9012 131501 9076
rect 131435 9011 131501 9012
rect 131990 6221 132050 77691
rect 132294 61954 132914 78000
rect 132294 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 132914 61954
rect 132294 61634 132914 61718
rect 132294 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 132914 61634
rect 132294 25954 132914 61398
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 131251 6220 131317 6221
rect 131251 6156 131252 6220
rect 131316 6156 131317 6220
rect 131251 6155 131317 6156
rect 131987 6220 132053 6221
rect 131987 6156 131988 6220
rect 132052 6156 132053 6220
rect 131987 6155 132053 6156
rect 131067 3500 131133 3501
rect 131067 3436 131068 3500
rect 131132 3436 131133 3500
rect 131067 3435 131133 3436
rect 127794 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 128414 -4186
rect 127794 -4506 128414 -4422
rect 127794 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 128414 -4506
rect 127794 -7654 128414 -4742
rect 132294 -5146 132914 25398
rect 133094 10301 133154 79731
rect 133278 76941 133338 79731
rect 133275 76940 133341 76941
rect 133275 76876 133276 76940
rect 133340 76876 133341 76940
rect 133275 76875 133341 76876
rect 133462 76669 133522 79867
rect 133827 77076 133893 77077
rect 133827 77012 133828 77076
rect 133892 77012 133893 77076
rect 133827 77011 133893 77012
rect 133459 76668 133525 76669
rect 133459 76604 133460 76668
rect 133524 76604 133525 76668
rect 133459 76603 133525 76604
rect 133275 75852 133341 75853
rect 133275 75788 133276 75852
rect 133340 75788 133341 75852
rect 133275 75787 133341 75788
rect 133278 44845 133338 75787
rect 133275 44844 133341 44845
rect 133275 44780 133276 44844
rect 133340 44780 133341 44844
rect 133275 44779 133341 44780
rect 133091 10300 133157 10301
rect 133091 10236 133092 10300
rect 133156 10236 133157 10300
rect 133091 10235 133157 10236
rect 133830 6357 133890 77011
rect 134014 7989 134074 79867
rect 134566 76669 134626 79867
rect 134195 76668 134261 76669
rect 134195 76604 134196 76668
rect 134260 76604 134261 76668
rect 134195 76603 134261 76604
rect 134563 76668 134629 76669
rect 134563 76604 134564 76668
rect 134628 76604 134629 76668
rect 134563 76603 134629 76604
rect 134198 10437 134258 76603
rect 135486 73170 135546 79867
rect 136406 76669 136466 79867
rect 136958 78165 137018 79867
rect 136955 78164 137021 78165
rect 136955 78100 136956 78164
rect 137020 78100 137021 78164
rect 136955 78099 137021 78100
rect 136403 76668 136469 76669
rect 136403 76604 136404 76668
rect 136468 76604 136469 76668
rect 136403 76603 136469 76604
rect 136403 76532 136469 76533
rect 136403 76468 136404 76532
rect 136468 76468 136469 76532
rect 136403 76467 136469 76468
rect 135302 73110 135546 73170
rect 135302 44981 135362 73110
rect 135299 44980 135365 44981
rect 135299 44916 135300 44980
rect 135364 44916 135365 44980
rect 135299 44915 135365 44916
rect 134195 10436 134261 10437
rect 134195 10372 134196 10436
rect 134260 10372 134261 10436
rect 134195 10371 134261 10372
rect 134011 7988 134077 7989
rect 134011 7924 134012 7988
rect 134076 7924 134077 7988
rect 134011 7923 134077 7924
rect 133827 6356 133893 6357
rect 133827 6292 133828 6356
rect 133892 6292 133893 6356
rect 133827 6291 133893 6292
rect 136406 3365 136466 76467
rect 136794 66454 137414 78000
rect 137691 76804 137757 76805
rect 137691 76740 137692 76804
rect 137756 76740 137757 76804
rect 137691 76739 137757 76740
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 136794 30454 137414 65898
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 136403 3364 136469 3365
rect 136403 3300 136404 3364
rect 136468 3300 136469 3364
rect 136403 3299 136469 3300
rect 132294 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 132914 -5146
rect 132294 -5466 132914 -5382
rect 132294 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 132914 -5466
rect 132294 -7654 132914 -5702
rect 136794 -6106 137414 29898
rect 137694 19957 137754 76739
rect 138062 76669 138122 79867
rect 138795 79796 138861 79797
rect 138795 79732 138796 79796
rect 138860 79732 138861 79796
rect 138795 79731 138861 79732
rect 139163 79796 139229 79797
rect 139163 79732 139164 79796
rect 139228 79732 139229 79796
rect 139163 79731 139229 79732
rect 140083 79796 140149 79797
rect 140083 79732 140084 79796
rect 140148 79732 140149 79796
rect 140083 79731 140149 79732
rect 137875 76668 137941 76669
rect 137875 76604 137876 76668
rect 137940 76604 137941 76668
rect 137875 76603 137941 76604
rect 138059 76668 138125 76669
rect 138059 76604 138060 76668
rect 138124 76604 138125 76668
rect 138059 76603 138125 76604
rect 137691 19956 137757 19957
rect 137691 19892 137692 19956
rect 137756 19892 137757 19956
rect 137691 19891 137757 19892
rect 137878 4861 137938 76603
rect 138798 60077 138858 79731
rect 138979 78708 139045 78709
rect 138979 78644 138980 78708
rect 139044 78644 139045 78708
rect 138979 78643 139045 78644
rect 138982 69597 139042 78643
rect 139166 75717 139226 79731
rect 139163 75716 139229 75717
rect 139163 75652 139164 75716
rect 139228 75652 139229 75716
rect 139163 75651 139229 75652
rect 138979 69596 139045 69597
rect 138979 69532 138980 69596
rect 139044 69532 139045 69596
rect 138979 69531 139045 69532
rect 138795 60076 138861 60077
rect 138795 60012 138796 60076
rect 138860 60012 138861 60076
rect 138795 60011 138861 60012
rect 140086 19005 140146 79731
rect 140270 65517 140330 79867
rect 140451 76396 140517 76397
rect 140451 76332 140452 76396
rect 140516 76332 140517 76396
rect 140451 76331 140517 76332
rect 140267 65516 140333 65517
rect 140267 65452 140268 65516
rect 140332 65452 140333 65516
rect 140267 65451 140333 65452
rect 140454 28525 140514 76331
rect 141003 75988 141069 75989
rect 141003 75924 141004 75988
rect 141068 75924 141069 75988
rect 141003 75923 141069 75924
rect 140451 28524 140517 28525
rect 140451 28460 140452 28524
rect 140516 28460 140517 28524
rect 140451 28459 140517 28460
rect 140083 19004 140149 19005
rect 140083 18940 140084 19004
rect 140148 18940 140149 19004
rect 140083 18939 140149 18940
rect 141006 10709 141066 75923
rect 141294 70954 141914 78000
rect 141294 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 141914 70954
rect 141294 70634 141914 70718
rect 141294 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 141914 70634
rect 141294 34954 141914 70398
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141003 10708 141069 10709
rect 141003 10644 141004 10708
rect 141068 10644 141069 10708
rect 141003 10643 141069 10644
rect 137875 4860 137941 4861
rect 137875 4796 137876 4860
rect 137940 4796 137941 4860
rect 137875 4795 137941 4796
rect 136794 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 137414 -6106
rect 136794 -6426 137414 -6342
rect 136794 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 137414 -6426
rect 136794 -7654 137414 -6662
rect 141294 -7066 141914 34398
rect 142846 28389 142906 80139
rect 144499 79932 144565 79933
rect 144499 79868 144500 79932
rect 144564 79868 144565 79932
rect 144499 79867 144565 79868
rect 145603 79932 145669 79933
rect 145603 79868 145604 79932
rect 145668 79868 145669 79932
rect 145603 79867 145669 79868
rect 146707 79932 146773 79933
rect 146707 79868 146708 79932
rect 146772 79868 146773 79932
rect 146707 79867 146773 79868
rect 147075 79932 147141 79933
rect 147075 79868 147076 79932
rect 147140 79868 147141 79932
rect 147075 79867 147141 79868
rect 147811 79932 147877 79933
rect 147811 79868 147812 79932
rect 147876 79868 147877 79932
rect 147811 79867 147877 79868
rect 148915 79932 148981 79933
rect 148915 79868 148916 79932
rect 148980 79868 148981 79932
rect 148915 79867 148981 79868
rect 149651 79932 149717 79933
rect 149651 79868 149652 79932
rect 149716 79868 149717 79932
rect 149651 79867 149717 79868
rect 151675 79932 151741 79933
rect 151675 79868 151676 79932
rect 151740 79930 151741 79932
rect 152779 79932 152845 79933
rect 152779 79930 152780 79932
rect 151740 79870 151922 79930
rect 151740 79868 151741 79870
rect 151675 79867 151741 79868
rect 144315 79660 144381 79661
rect 144315 79596 144316 79660
rect 144380 79596 144381 79660
rect 144315 79595 144381 79596
rect 144318 78845 144378 79595
rect 144315 78844 144381 78845
rect 144315 78780 144316 78844
rect 144380 78780 144381 78844
rect 144315 78779 144381 78780
rect 144131 76124 144197 76125
rect 144131 76060 144132 76124
rect 144196 76060 144197 76124
rect 144131 76059 144197 76060
rect 143211 75988 143277 75989
rect 143211 75924 143212 75988
rect 143276 75924 143277 75988
rect 143211 75923 143277 75924
rect 143027 75852 143093 75853
rect 143027 75788 143028 75852
rect 143092 75788 143093 75852
rect 143027 75787 143093 75788
rect 143030 59941 143090 75787
rect 143027 59940 143093 59941
rect 143027 59876 143028 59940
rect 143092 59876 143093 59940
rect 143027 59875 143093 59876
rect 143214 34101 143274 75923
rect 143211 34100 143277 34101
rect 143211 34036 143212 34100
rect 143276 34036 143277 34100
rect 143211 34035 143277 34036
rect 142843 28388 142909 28389
rect 142843 28324 142844 28388
rect 142908 28324 142909 28388
rect 142843 28323 142909 28324
rect 144134 7717 144194 76059
rect 144502 20229 144562 79867
rect 145235 78572 145301 78573
rect 145235 78508 145236 78572
rect 145300 78508 145301 78572
rect 145235 78507 145301 78508
rect 145238 33965 145298 78507
rect 145419 75988 145485 75989
rect 145419 75924 145420 75988
rect 145484 75924 145485 75988
rect 145419 75923 145485 75924
rect 145235 33964 145301 33965
rect 145235 33900 145236 33964
rect 145300 33900 145301 33964
rect 145235 33899 145301 33900
rect 144499 20228 144565 20229
rect 144499 20164 144500 20228
rect 144564 20164 144565 20228
rect 144499 20163 144565 20164
rect 145422 9213 145482 75923
rect 145419 9212 145485 9213
rect 145419 9148 145420 9212
rect 145484 9148 145485 9212
rect 145419 9147 145485 9148
rect 144131 7716 144197 7717
rect 144131 7652 144132 7716
rect 144196 7652 144197 7716
rect 144131 7651 144197 7652
rect 145606 7581 145666 79867
rect 146155 79660 146221 79661
rect 146155 79596 146156 79660
rect 146220 79596 146221 79660
rect 146155 79595 146221 79596
rect 146158 78845 146218 79595
rect 146155 78844 146221 78845
rect 146155 78780 146156 78844
rect 146220 78780 146221 78844
rect 146155 78779 146221 78780
rect 146710 78029 146770 79867
rect 147078 78029 147138 79867
rect 146707 78028 146773 78029
rect 145794 75454 146414 78000
rect 146707 77964 146708 78028
rect 146772 77964 146773 78028
rect 146707 77963 146773 77964
rect 147075 78028 147141 78029
rect 147075 77964 147076 78028
rect 147140 77964 147141 78028
rect 147075 77963 147141 77964
rect 147259 78028 147325 78029
rect 147259 77964 147260 78028
rect 147324 77964 147325 78028
rect 147259 77963 147325 77964
rect 147075 77348 147141 77349
rect 147075 77284 147076 77348
rect 147140 77284 147141 77348
rect 147075 77283 147141 77284
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145603 7580 145669 7581
rect 145603 7516 145604 7580
rect 145668 7516 145669 7580
rect 145603 7515 145669 7516
rect 141294 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 141914 -7066
rect 141294 -7386 141914 -7302
rect 141294 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 141914 -7386
rect 141294 -7654 141914 -7622
rect 145794 3454 146414 38898
rect 147078 10573 147138 77283
rect 147262 44845 147322 77963
rect 147814 75989 147874 79867
rect 148547 78436 148613 78437
rect 148547 78372 148548 78436
rect 148612 78372 148613 78436
rect 148547 78371 148613 78372
rect 148363 77892 148429 77893
rect 148363 77828 148364 77892
rect 148428 77828 148429 77892
rect 148363 77827 148429 77828
rect 147811 75988 147877 75989
rect 147811 75924 147812 75988
rect 147876 75924 147877 75988
rect 147811 75923 147877 75924
rect 148366 72453 148426 77827
rect 148363 72452 148429 72453
rect 148363 72388 148364 72452
rect 148428 72388 148429 72452
rect 148363 72387 148429 72388
rect 147259 44844 147325 44845
rect 147259 44780 147260 44844
rect 147324 44780 147325 44844
rect 147259 44779 147325 44780
rect 148550 13293 148610 78371
rect 148731 75988 148797 75989
rect 148731 75924 148732 75988
rect 148796 75924 148797 75988
rect 148731 75923 148797 75924
rect 148547 13292 148613 13293
rect 148547 13228 148548 13292
rect 148612 13228 148613 13292
rect 148547 13227 148613 13228
rect 147075 10572 147141 10573
rect 147075 10508 147076 10572
rect 147140 10508 147141 10572
rect 147075 10507 147141 10508
rect 148734 10437 148794 75923
rect 148731 10436 148797 10437
rect 148731 10372 148732 10436
rect 148796 10372 148797 10436
rect 148731 10371 148797 10372
rect 148918 9077 148978 79867
rect 149467 78572 149533 78573
rect 149467 78508 149468 78572
rect 149532 78508 149533 78572
rect 149467 78507 149533 78508
rect 149470 53141 149530 78507
rect 149467 53140 149533 53141
rect 149467 53076 149468 53140
rect 149532 53076 149533 53140
rect 149467 53075 149533 53076
rect 149654 29613 149714 79867
rect 149835 79796 149901 79797
rect 149835 79732 149836 79796
rect 149900 79732 149901 79796
rect 149835 79731 149901 79732
rect 151491 79796 151557 79797
rect 151491 79732 151492 79796
rect 151556 79732 151557 79796
rect 151491 79731 151557 79732
rect 149651 29612 149717 29613
rect 149651 29548 149652 29612
rect 149716 29548 149717 29612
rect 149651 29547 149717 29548
rect 149838 16285 149898 79731
rect 150019 78708 150085 78709
rect 150019 78644 150020 78708
rect 150084 78644 150085 78708
rect 150019 78643 150085 78644
rect 149835 16284 149901 16285
rect 149835 16220 149836 16284
rect 149900 16220 149901 16284
rect 149835 16219 149901 16220
rect 148915 9076 148981 9077
rect 148915 9012 148916 9076
rect 148980 9012 148981 9076
rect 148915 9011 148981 9012
rect 150022 5133 150082 78643
rect 150294 43954 150914 78000
rect 151307 76532 151373 76533
rect 151307 76468 151308 76532
rect 151372 76468 151373 76532
rect 151307 76467 151373 76468
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 150294 7954 150914 43398
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150019 5132 150085 5133
rect 150019 5068 150020 5132
rect 150084 5068 150085 5132
rect 150019 5067 150085 5068
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 150294 -1306 150914 7398
rect 151310 6493 151370 76467
rect 151307 6492 151373 6493
rect 151307 6428 151308 6492
rect 151372 6428 151373 6492
rect 151307 6427 151373 6428
rect 151494 6357 151554 79731
rect 151675 76668 151741 76669
rect 151675 76604 151676 76668
rect 151740 76604 151741 76668
rect 151675 76603 151741 76604
rect 151491 6356 151557 6357
rect 151491 6292 151492 6356
rect 151556 6292 151557 6356
rect 151491 6291 151557 6292
rect 151678 3637 151738 76603
rect 151862 76397 151922 79870
rect 152414 79870 152780 79930
rect 151859 76396 151925 76397
rect 151859 76332 151860 76396
rect 151924 76332 151925 76396
rect 151859 76331 151925 76332
rect 152414 13157 152474 79870
rect 152779 79868 152780 79870
rect 152844 79868 152845 79932
rect 152779 79867 152845 79868
rect 154067 79932 154133 79933
rect 154067 79868 154068 79932
rect 154132 79868 154133 79932
rect 154067 79867 154133 79868
rect 154251 79932 154317 79933
rect 154251 79868 154252 79932
rect 154316 79868 154317 79932
rect 154251 79867 154317 79868
rect 154987 79932 155053 79933
rect 154987 79868 154988 79932
rect 155052 79868 155053 79932
rect 154987 79867 155053 79868
rect 155723 79932 155789 79933
rect 155723 79868 155724 79932
rect 155788 79868 155789 79932
rect 155723 79867 155789 79868
rect 156091 79932 156157 79933
rect 156091 79868 156092 79932
rect 156156 79868 156157 79932
rect 156091 79867 156157 79868
rect 156827 79932 156893 79933
rect 156827 79868 156828 79932
rect 156892 79868 156893 79932
rect 156827 79867 156893 79868
rect 157747 79932 157813 79933
rect 157747 79868 157748 79932
rect 157812 79868 157813 79932
rect 157747 79867 157813 79868
rect 158115 79932 158181 79933
rect 158115 79868 158116 79932
rect 158180 79868 158181 79932
rect 158115 79867 158181 79868
rect 153883 79796 153949 79797
rect 153883 79732 153884 79796
rect 153948 79732 153949 79796
rect 153883 79731 153949 79732
rect 152595 77076 152661 77077
rect 152595 77012 152596 77076
rect 152660 77012 152661 77076
rect 152595 77011 152661 77012
rect 152598 47565 152658 77011
rect 152963 76668 153029 76669
rect 152963 76604 152964 76668
rect 153028 76604 153029 76668
rect 152963 76603 153029 76604
rect 152779 76532 152845 76533
rect 152779 76468 152780 76532
rect 152844 76468 152845 76532
rect 152779 76467 152845 76468
rect 152595 47564 152661 47565
rect 152595 47500 152596 47564
rect 152660 47500 152661 47564
rect 152595 47499 152661 47500
rect 152782 18869 152842 76467
rect 152966 71229 153026 76603
rect 152963 71228 153029 71229
rect 152963 71164 152964 71228
rect 153028 71164 153029 71228
rect 152963 71163 153029 71164
rect 153886 40629 153946 79731
rect 154070 76669 154130 79867
rect 154067 76668 154133 76669
rect 154067 76604 154068 76668
rect 154132 76604 154133 76668
rect 154067 76603 154133 76604
rect 154067 76532 154133 76533
rect 154067 76468 154068 76532
rect 154132 76468 154133 76532
rect 154067 76467 154133 76468
rect 153883 40628 153949 40629
rect 153883 40564 153884 40628
rect 153948 40564 153949 40628
rect 153883 40563 153949 40564
rect 154070 35189 154130 76467
rect 154067 35188 154133 35189
rect 154067 35124 154068 35188
rect 154132 35124 154133 35188
rect 154067 35123 154133 35124
rect 152779 18868 152845 18869
rect 152779 18804 152780 18868
rect 152844 18804 152845 18868
rect 152779 18803 152845 18804
rect 154254 16149 154314 79867
rect 154990 78165 155050 79867
rect 154987 78164 155053 78165
rect 154987 78100 154988 78164
rect 155052 78100 155053 78164
rect 154987 78099 155053 78100
rect 154435 76668 154501 76669
rect 154435 76604 154436 76668
rect 154500 76604 154501 76668
rect 154435 76603 154501 76604
rect 154251 16148 154317 16149
rect 154251 16084 154252 16148
rect 154316 16084 154317 16148
rect 154251 16083 154317 16084
rect 154438 14789 154498 76603
rect 154794 48454 155414 78000
rect 155539 76668 155605 76669
rect 155539 76604 155540 76668
rect 155604 76604 155605 76668
rect 155539 76603 155605 76604
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 154435 14788 154501 14789
rect 154435 14724 154436 14788
rect 154500 14724 154501 14788
rect 154435 14723 154501 14724
rect 152411 13156 152477 13157
rect 152411 13092 152412 13156
rect 152476 13092 152477 13156
rect 152411 13091 152477 13092
rect 154794 12454 155414 47898
rect 155542 25533 155602 76603
rect 155539 25532 155605 25533
rect 155539 25468 155540 25532
rect 155604 25468 155605 25532
rect 155539 25467 155605 25468
rect 155726 16013 155786 79867
rect 156094 76669 156154 79867
rect 156091 76668 156157 76669
rect 156091 76604 156092 76668
rect 156156 76604 156157 76668
rect 156091 76603 156157 76604
rect 156643 76668 156709 76669
rect 156643 76604 156644 76668
rect 156708 76604 156709 76668
rect 156643 76603 156709 76604
rect 155723 16012 155789 16013
rect 155723 15948 155724 16012
rect 155788 15948 155789 16012
rect 155723 15947 155789 15948
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 151675 3636 151741 3637
rect 151675 3572 151676 3636
rect 151740 3572 151741 3636
rect 151675 3571 151741 3572
rect 150294 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 150914 -1306
rect 150294 -1626 150914 -1542
rect 150294 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 150914 -1626
rect 150294 -7654 150914 -1862
rect 154794 -2266 155414 11898
rect 156646 8941 156706 76603
rect 156830 17373 156890 79867
rect 157011 79796 157077 79797
rect 157011 79732 157012 79796
rect 157076 79732 157077 79796
rect 157011 79731 157077 79732
rect 156827 17372 156893 17373
rect 156827 17308 156828 17372
rect 156892 17308 156893 17372
rect 156827 17307 156893 17308
rect 157014 14653 157074 79731
rect 157750 76669 157810 79867
rect 157747 76668 157813 76669
rect 157747 76604 157748 76668
rect 157812 76604 157813 76668
rect 157747 76603 157813 76604
rect 157931 76532 157997 76533
rect 157931 76468 157932 76532
rect 157996 76468 157997 76532
rect 157931 76467 157997 76468
rect 157934 24173 157994 76467
rect 157931 24172 157997 24173
rect 157931 24108 157932 24172
rect 157996 24108 157997 24172
rect 157931 24107 157997 24108
rect 158118 18733 158178 79867
rect 158299 79796 158365 79797
rect 158299 79732 158300 79796
rect 158364 79732 158365 79796
rect 158299 79731 158365 79732
rect 159035 79796 159101 79797
rect 159035 79732 159036 79796
rect 159100 79732 159101 79796
rect 159035 79731 159101 79732
rect 158115 18732 158181 18733
rect 158115 18668 158116 18732
rect 158180 18668 158181 18732
rect 158115 18667 158181 18668
rect 158302 15877 158362 79731
rect 158483 76668 158549 76669
rect 158483 76604 158484 76668
rect 158548 76604 158549 76668
rect 158483 76603 158549 76604
rect 158299 15876 158365 15877
rect 158299 15812 158300 15876
rect 158364 15812 158365 15876
rect 158299 15811 158365 15812
rect 157011 14652 157077 14653
rect 157011 14588 157012 14652
rect 157076 14588 157077 14652
rect 157011 14587 157077 14588
rect 158486 11797 158546 76603
rect 158851 76260 158917 76261
rect 158851 76196 158852 76260
rect 158916 76196 158917 76260
rect 158851 76195 158917 76196
rect 158854 21589 158914 76195
rect 158851 21588 158917 21589
rect 158851 21524 158852 21588
rect 158916 21524 158917 21588
rect 158851 21523 158917 21524
rect 158483 11796 158549 11797
rect 158483 11732 158484 11796
rect 158548 11732 158549 11796
rect 158483 11731 158549 11732
rect 156643 8940 156709 8941
rect 156643 8876 156644 8940
rect 156708 8876 156709 8940
rect 156643 8875 156709 8876
rect 159038 4997 159098 79731
rect 159222 79117 159282 80139
rect 171182 79933 171242 80683
rect 171363 80612 171429 80613
rect 171363 80548 171364 80612
rect 171428 80548 171429 80612
rect 171363 80547 171429 80548
rect 161243 79932 161309 79933
rect 161243 79868 161244 79932
rect 161308 79868 161309 79932
rect 161243 79867 161309 79868
rect 162715 79932 162781 79933
rect 162715 79868 162716 79932
rect 162780 79868 162781 79932
rect 162715 79867 162781 79868
rect 163451 79932 163517 79933
rect 163451 79868 163452 79932
rect 163516 79868 163517 79932
rect 163451 79867 163517 79868
rect 164923 79932 164989 79933
rect 164923 79868 164924 79932
rect 164988 79868 164989 79932
rect 164923 79867 164989 79868
rect 165107 79932 165173 79933
rect 165107 79868 165108 79932
rect 165172 79868 165173 79932
rect 165107 79867 165173 79868
rect 166395 79932 166461 79933
rect 166395 79868 166396 79932
rect 166460 79868 166461 79932
rect 166395 79867 166461 79868
rect 167499 79932 167565 79933
rect 167499 79868 167500 79932
rect 167564 79868 167565 79932
rect 167499 79867 167565 79868
rect 169155 79932 169221 79933
rect 169155 79868 169156 79932
rect 169220 79868 169221 79932
rect 169155 79867 169221 79868
rect 169339 79932 169405 79933
rect 169339 79868 169340 79932
rect 169404 79868 169405 79932
rect 169339 79867 169405 79868
rect 170443 79932 170509 79933
rect 170443 79868 170444 79932
rect 170508 79868 170509 79932
rect 170443 79867 170509 79868
rect 171179 79932 171245 79933
rect 171179 79868 171180 79932
rect 171244 79868 171245 79932
rect 171179 79867 171245 79868
rect 160139 79660 160205 79661
rect 160139 79596 160140 79660
rect 160204 79596 160205 79660
rect 160139 79595 160205 79596
rect 159219 79116 159285 79117
rect 159219 79052 159220 79116
rect 159284 79052 159285 79116
rect 159219 79051 159285 79052
rect 160142 78573 160202 79595
rect 161246 79117 161306 79867
rect 162347 79796 162413 79797
rect 162347 79732 162348 79796
rect 162412 79732 162413 79796
rect 162347 79731 162413 79732
rect 161243 79116 161309 79117
rect 161243 79052 161244 79116
rect 161308 79052 161309 79116
rect 161243 79051 161309 79052
rect 160139 78572 160205 78573
rect 160139 78508 160140 78572
rect 160204 78508 160205 78572
rect 160139 78507 160205 78508
rect 159294 52954 159914 78000
rect 161243 77348 161309 77349
rect 161243 77284 161244 77348
rect 161308 77284 161309 77348
rect 161243 77283 161309 77284
rect 160875 76668 160941 76669
rect 160875 76604 160876 76668
rect 160940 76604 160941 76668
rect 160875 76603 160941 76604
rect 160691 76532 160757 76533
rect 160691 76468 160692 76532
rect 160756 76468 160757 76532
rect 160691 76467 160757 76468
rect 160694 61437 160754 76467
rect 160691 61436 160757 61437
rect 160691 61372 160692 61436
rect 160756 61372 160757 61436
rect 160691 61371 160757 61372
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159294 16954 159914 52398
rect 160878 21453 160938 76603
rect 161059 76396 161125 76397
rect 161059 76332 161060 76396
rect 161124 76332 161125 76396
rect 161059 76331 161125 76332
rect 160875 21452 160941 21453
rect 160875 21388 160876 21452
rect 160940 21388 160941 21452
rect 160875 21387 160941 21388
rect 161062 20093 161122 76331
rect 161059 20092 161125 20093
rect 161059 20028 161060 20092
rect 161124 20028 161125 20092
rect 161059 20027 161125 20028
rect 161246 17237 161306 77283
rect 162350 21317 162410 79731
rect 162531 79660 162597 79661
rect 162531 79596 162532 79660
rect 162596 79596 162597 79660
rect 162531 79595 162597 79596
rect 162347 21316 162413 21317
rect 162347 21252 162348 21316
rect 162412 21252 162413 21316
rect 162347 21251 162413 21252
rect 161243 17236 161309 17237
rect 161243 17172 161244 17236
rect 161308 17172 161309 17236
rect 161243 17171 161309 17172
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 159035 4996 159101 4997
rect 159035 4932 159036 4996
rect 159100 4932 159101 4996
rect 159035 4931 159101 4932
rect 154794 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 155414 -2266
rect 154794 -2586 155414 -2502
rect 154794 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 155414 -2586
rect 154794 -7654 155414 -2822
rect 159294 -3226 159914 16398
rect 162534 14517 162594 79595
rect 162531 14516 162597 14517
rect 162531 14452 162532 14516
rect 162596 14452 162597 14516
rect 162531 14451 162597 14452
rect 162718 11661 162778 79867
rect 163454 71093 163514 79867
rect 164371 79660 164437 79661
rect 164371 79596 164372 79660
rect 164436 79596 164437 79660
rect 164371 79595 164437 79596
rect 163635 79116 163701 79117
rect 163635 79052 163636 79116
rect 163700 79052 163701 79116
rect 163635 79051 163701 79052
rect 163451 71092 163517 71093
rect 163451 71028 163452 71092
rect 163516 71028 163517 71092
rect 163451 71027 163517 71028
rect 163638 19957 163698 79051
rect 164374 78570 164434 79595
rect 164374 78510 164618 78570
rect 163794 57454 164414 78000
rect 164558 75309 164618 78510
rect 164926 76669 164986 79867
rect 164923 76668 164989 76669
rect 164923 76604 164924 76668
rect 164988 76604 164989 76668
rect 164923 76603 164989 76604
rect 164923 76532 164989 76533
rect 164923 76468 164924 76532
rect 164988 76468 164989 76532
rect 164923 76467 164989 76468
rect 164555 75308 164621 75309
rect 164555 75244 164556 75308
rect 164620 75244 164621 75308
rect 164555 75243 164621 75244
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163635 19956 163701 19957
rect 163635 19892 163636 19956
rect 163700 19892 163701 19956
rect 163635 19891 163701 19892
rect 162715 11660 162781 11661
rect 162715 11596 162716 11660
rect 162780 11596 162781 11660
rect 162715 11595 162781 11596
rect 159294 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 159914 -3226
rect 159294 -3546 159914 -3462
rect 159294 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 159914 -3546
rect 159294 -7654 159914 -3782
rect 163794 -4186 164414 20898
rect 164926 10301 164986 76467
rect 165110 28253 165170 79867
rect 165291 79796 165357 79797
rect 165291 79732 165292 79796
rect 165356 79732 165357 79796
rect 165291 79731 165357 79732
rect 165107 28252 165173 28253
rect 165107 28188 165108 28252
rect 165172 28188 165173 28252
rect 165107 28187 165173 28188
rect 165294 27029 165354 79731
rect 165475 76668 165541 76669
rect 165475 76604 165476 76668
rect 165540 76604 165541 76668
rect 165475 76603 165541 76604
rect 165478 68237 165538 76603
rect 165475 68236 165541 68237
rect 165475 68172 165476 68236
rect 165540 68172 165541 68236
rect 165475 68171 165541 68172
rect 166398 62933 166458 79867
rect 166579 79796 166645 79797
rect 166579 79732 166580 79796
rect 166644 79732 166645 79796
rect 166579 79731 166645 79732
rect 166395 62932 166461 62933
rect 166395 62868 166396 62932
rect 166460 62868 166461 62932
rect 166395 62867 166461 62868
rect 166582 32605 166642 79731
rect 166763 76668 166829 76669
rect 166763 76604 166764 76668
rect 166828 76604 166829 76668
rect 166763 76603 166829 76604
rect 166579 32604 166645 32605
rect 166579 32540 166580 32604
rect 166644 32540 166645 32604
rect 166579 32539 166645 32540
rect 165291 27028 165357 27029
rect 165291 26964 165292 27028
rect 165356 26964 165357 27028
rect 165291 26963 165357 26964
rect 166766 13021 166826 76603
rect 167502 76397 167562 79867
rect 167867 79660 167933 79661
rect 167867 79596 167868 79660
rect 167932 79596 167933 79660
rect 167867 79595 167933 79596
rect 167683 78708 167749 78709
rect 167683 78644 167684 78708
rect 167748 78644 167749 78708
rect 167683 78643 167749 78644
rect 167499 76396 167565 76397
rect 167499 76332 167500 76396
rect 167564 76332 167565 76396
rect 167499 76331 167565 76332
rect 167686 30973 167746 78643
rect 167683 30972 167749 30973
rect 167683 30908 167684 30972
rect 167748 30908 167749 30972
rect 167683 30907 167749 30908
rect 167870 18597 167930 79595
rect 168051 76668 168117 76669
rect 168051 76604 168052 76668
rect 168116 76604 168117 76668
rect 168051 76603 168117 76604
rect 167867 18596 167933 18597
rect 167867 18532 167868 18596
rect 167932 18532 167933 18596
rect 167867 18531 167933 18532
rect 166763 13020 166829 13021
rect 166763 12956 166764 13020
rect 166828 12956 166829 13020
rect 166763 12955 166829 12956
rect 164923 10300 164989 10301
rect 164923 10236 164924 10300
rect 164988 10236 164989 10300
rect 164923 10235 164989 10236
rect 168054 4861 168114 76603
rect 168294 61954 168914 78000
rect 169158 77349 169218 79867
rect 169155 77348 169221 77349
rect 169155 77284 169156 77348
rect 169220 77284 169221 77348
rect 169155 77283 169221 77284
rect 169342 76533 169402 79867
rect 170075 78708 170141 78709
rect 170075 78644 170076 78708
rect 170140 78644 170141 78708
rect 170075 78643 170141 78644
rect 169339 76532 169405 76533
rect 169339 76468 169340 76532
rect 169404 76468 169405 76532
rect 169339 76467 169405 76468
rect 169339 76124 169405 76125
rect 169339 76060 169340 76124
rect 169404 76060 169405 76124
rect 169339 76059 169405 76060
rect 168294 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 168914 61954
rect 168294 61634 168914 61718
rect 168294 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 168914 61634
rect 168294 25954 168914 61398
rect 169342 32469 169402 76059
rect 170078 75853 170138 78643
rect 170075 75852 170141 75853
rect 170075 75788 170076 75852
rect 170140 75788 170141 75852
rect 170075 75787 170141 75788
rect 169339 32468 169405 32469
rect 169339 32404 169340 32468
rect 169404 32404 169405 32468
rect 169339 32403 169405 32404
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168051 4860 168117 4861
rect 168051 4796 168052 4860
rect 168116 4796 168117 4860
rect 168051 4795 168117 4796
rect 163794 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 164414 -4186
rect 163794 -4506 164414 -4422
rect 163794 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 164414 -4506
rect 163794 -7654 164414 -4742
rect 168294 -5146 168914 25398
rect 170446 21725 170506 79867
rect 171366 79797 171426 80547
rect 171363 79796 171429 79797
rect 171363 79732 171364 79796
rect 171428 79732 171429 79796
rect 171363 79731 171429 79732
rect 170627 79660 170693 79661
rect 170627 79596 170628 79660
rect 170692 79596 170693 79660
rect 170627 79595 170693 79596
rect 170630 33829 170690 79595
rect 171550 78845 171610 81091
rect 173203 80476 173269 80477
rect 173203 80412 173204 80476
rect 173268 80412 173269 80476
rect 173203 80411 173269 80412
rect 171915 79932 171981 79933
rect 171915 79868 171916 79932
rect 171980 79868 171981 79932
rect 171915 79867 171981 79868
rect 172421 79932 172487 79933
rect 172421 79868 172422 79932
rect 172486 79930 172487 79932
rect 172486 79868 172530 79930
rect 172421 79867 172530 79868
rect 171918 78981 171978 79867
rect 171915 78980 171981 78981
rect 171915 78916 171916 78980
rect 171980 78916 171981 78980
rect 171915 78915 171981 78916
rect 171547 78844 171613 78845
rect 171547 78780 171548 78844
rect 171612 78780 171613 78844
rect 171547 78779 171613 78780
rect 172470 78709 172530 79867
rect 173206 79525 173266 80411
rect 173574 79661 173634 81227
rect 186294 79954 186914 115398
rect 186294 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 186914 79954
rect 173571 79660 173637 79661
rect 173571 79596 173572 79660
rect 173636 79596 173637 79660
rect 173571 79595 173637 79596
rect 186294 79634 186914 79718
rect 173203 79524 173269 79525
rect 173203 79460 173204 79524
rect 173268 79460 173269 79524
rect 173203 79459 173269 79460
rect 186294 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 186914 79634
rect 170995 78708 171061 78709
rect 170995 78644 170996 78708
rect 171060 78644 171061 78708
rect 170995 78643 171061 78644
rect 172467 78708 172533 78709
rect 172467 78644 172468 78708
rect 172532 78644 172533 78708
rect 172467 78643 172533 78644
rect 170811 76260 170877 76261
rect 170811 76196 170812 76260
rect 170876 76196 170877 76260
rect 170811 76195 170877 76196
rect 170627 33828 170693 33829
rect 170627 33764 170628 33828
rect 170692 33764 170693 33828
rect 170627 33763 170693 33764
rect 170814 26893 170874 76195
rect 170998 76125 171058 78643
rect 171179 77348 171245 77349
rect 171179 77284 171180 77348
rect 171244 77284 171245 77348
rect 171179 77283 171245 77284
rect 170995 76124 171061 76125
rect 170995 76060 170996 76124
rect 171060 76060 171061 76124
rect 170995 76059 171061 76060
rect 171182 62797 171242 77283
rect 171731 75988 171797 75989
rect 171731 75924 171732 75988
rect 171796 75924 171797 75988
rect 171731 75923 171797 75924
rect 171179 62796 171245 62797
rect 171179 62732 171180 62796
rect 171244 62732 171245 62796
rect 171179 62731 171245 62732
rect 170811 26892 170877 26893
rect 170811 26828 170812 26892
rect 170876 26828 170877 26892
rect 170811 26827 170877 26828
rect 170443 21724 170509 21725
rect 170443 21660 170444 21724
rect 170508 21660 170509 21724
rect 170443 21659 170509 21660
rect 171734 3501 171794 75923
rect 171915 75852 171981 75853
rect 171915 75788 171916 75852
rect 171980 75788 171981 75852
rect 171915 75787 171981 75788
rect 171731 3500 171797 3501
rect 171731 3436 171732 3500
rect 171796 3436 171797 3500
rect 171731 3435 171797 3436
rect 171918 3365 171978 75787
rect 172794 66454 173414 78000
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 172794 30454 173414 65898
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 171915 3364 171981 3365
rect 171915 3300 171916 3364
rect 171980 3300 171981 3364
rect 171915 3299 171981 3300
rect 168294 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 168914 -5146
rect 168294 -5466 168914 -5382
rect 168294 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 168914 -5466
rect 168294 -7654 168914 -5702
rect 172794 -6106 173414 29898
rect 172794 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 173414 -6106
rect 172794 -6426 173414 -6342
rect 172794 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 173414 -6426
rect 172794 -7654 173414 -6662
rect 177294 70954 177914 78000
rect 177294 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 177914 70954
rect 177294 70634 177914 70718
rect 177294 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 177914 70634
rect 177294 34954 177914 70398
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 177294 -7066 177914 34398
rect 177294 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 177914 -7066
rect 177294 -7386 177914 -7302
rect 177294 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 177914 -7386
rect 177294 -7654 177914 -7622
rect 181794 75454 182414 78000
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 186294 43954 186914 79398
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 186294 7954 186914 43398
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1306 186914 7398
rect 186294 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 186914 -1306
rect 186294 -1626 186914 -1542
rect 186294 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 186914 -1626
rect 186294 -7654 186914 -1862
rect 190794 228453 191414 228484
rect 190794 228217 190826 228453
rect 191062 228217 191146 228453
rect 191382 228217 191414 228453
rect 190794 228133 191414 228217
rect 190794 227897 190826 228133
rect 191062 227897 191146 228133
rect 191382 227897 191414 228133
rect 190794 192454 191414 227897
rect 190794 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 191414 192454
rect 190794 192134 191414 192218
rect 190794 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 191414 192134
rect 190794 156454 191414 191898
rect 190794 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 191414 156454
rect 190794 156134 191414 156218
rect 190794 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 191414 156134
rect 190794 120454 191414 155898
rect 190794 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 191414 120454
rect 190794 120134 191414 120218
rect 190794 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 191414 120134
rect 190794 84454 191414 119898
rect 190794 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 191414 84454
rect 190794 84134 191414 84218
rect 190794 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 191414 84134
rect 190794 48454 191414 83898
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 190794 12454 191414 47898
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2266 191414 11898
rect 190794 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 191414 -2266
rect 190794 -2586 191414 -2502
rect 190794 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 191414 -2586
rect 190794 -7654 191414 -2822
rect 195294 196954 195914 228484
rect 195294 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 195914 196954
rect 195294 196634 195914 196718
rect 195294 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 195914 196634
rect 195294 160954 195914 196398
rect 195294 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 195914 160954
rect 195294 160634 195914 160718
rect 195294 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 195914 160634
rect 195294 124954 195914 160398
rect 195294 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 195914 124954
rect 195294 124634 195914 124718
rect 195294 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 195914 124634
rect 195294 88954 195914 124398
rect 195294 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 195914 88954
rect 195294 88634 195914 88718
rect 195294 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 195914 88634
rect 195294 52954 195914 88398
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 195294 16954 195914 52398
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3226 195914 16398
rect 195294 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 195914 -3226
rect 195294 -3546 195914 -3462
rect 195294 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 195914 -3546
rect 195294 -7654 195914 -3782
rect 199794 201454 200414 228484
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4186 200414 20898
rect 199794 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 200414 -4186
rect 199794 -4506 200414 -4422
rect 199794 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 200414 -4506
rect 199794 -7654 200414 -4742
rect 204294 205954 204914 228484
rect 204294 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 204914 205954
rect 204294 205634 204914 205718
rect 204294 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 204914 205634
rect 204294 169954 204914 205398
rect 204294 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 204914 169954
rect 204294 169634 204914 169718
rect 204294 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 204914 169634
rect 204294 133954 204914 169398
rect 204294 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 204914 133954
rect 204294 133634 204914 133718
rect 204294 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 204914 133634
rect 204294 97954 204914 133398
rect 204294 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 204914 97954
rect 204294 97634 204914 97718
rect 204294 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 204914 97634
rect 204294 61954 204914 97398
rect 204294 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 204914 61954
rect 204294 61634 204914 61718
rect 204294 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 204914 61634
rect 204294 25954 204914 61398
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5146 204914 25398
rect 204294 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 204914 -5146
rect 204294 -5466 204914 -5382
rect 204294 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 204914 -5466
rect 204294 -7654 204914 -5702
rect 208794 210454 209414 228484
rect 208794 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 209414 210454
rect 208794 210134 209414 210218
rect 208794 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 209414 210134
rect 208794 174454 209414 209898
rect 208794 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 209414 174454
rect 208794 174134 209414 174218
rect 208794 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 209414 174134
rect 208794 138454 209414 173898
rect 208794 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 209414 138454
rect 208794 138134 209414 138218
rect 208794 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 209414 138134
rect 208794 102454 209414 137898
rect 208794 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 209414 102454
rect 208794 102134 209414 102218
rect 208794 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 209414 102134
rect 208794 66454 209414 101898
rect 208794 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 209414 66454
rect 208794 66134 209414 66218
rect 208794 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 209414 66134
rect 208794 30454 209414 65898
rect 208794 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 209414 30454
rect 208794 30134 209414 30218
rect 208794 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 209414 30134
rect 208794 -6106 209414 29898
rect 208794 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 209414 -6106
rect 208794 -6426 209414 -6342
rect 208794 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 209414 -6426
rect 208794 -7654 209414 -6662
rect 213294 214954 213914 228484
rect 213294 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 213914 214954
rect 213294 214634 213914 214718
rect 213294 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 213914 214634
rect 213294 178954 213914 214398
rect 213294 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 213914 178954
rect 213294 178634 213914 178718
rect 213294 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 213914 178634
rect 213294 142954 213914 178398
rect 213294 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 213914 142954
rect 213294 142634 213914 142718
rect 213294 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 213914 142634
rect 213294 106954 213914 142398
rect 213294 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 213914 106954
rect 213294 106634 213914 106718
rect 213294 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 213914 106634
rect 213294 70954 213914 106398
rect 213294 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 213914 70954
rect 213294 70634 213914 70718
rect 213294 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 213914 70634
rect 213294 34954 213914 70398
rect 213294 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 213914 34954
rect 213294 34634 213914 34718
rect 213294 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 213914 34634
rect 213294 -7066 213914 34398
rect 213294 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 213914 -7066
rect 213294 -7386 213914 -7302
rect 213294 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 213914 -7386
rect 213294 -7654 213914 -7622
rect 217794 219454 218414 228484
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 222294 223954 222914 228484
rect 222294 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 222914 223954
rect 222294 223634 222914 223718
rect 222294 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 222914 223634
rect 222294 187954 222914 223398
rect 222294 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 222914 187954
rect 222294 187634 222914 187718
rect 222294 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 222914 187634
rect 222294 151954 222914 187398
rect 222294 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 222914 151954
rect 222294 151634 222914 151718
rect 222294 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 222914 151634
rect 222294 115954 222914 151398
rect 222294 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 222914 115954
rect 222294 115634 222914 115718
rect 222294 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 222914 115634
rect 222294 79954 222914 115398
rect 222294 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 222914 79954
rect 222294 79634 222914 79718
rect 222294 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 222914 79634
rect 222294 43954 222914 79398
rect 222294 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 222914 43954
rect 222294 43634 222914 43718
rect 222294 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 222914 43634
rect 222294 7954 222914 43398
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 222294 -1306 222914 7398
rect 222294 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 222914 -1306
rect 222294 -1626 222914 -1542
rect 222294 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 222914 -1626
rect 222294 -7654 222914 -1862
rect 226794 228453 227414 228484
rect 226794 228217 226826 228453
rect 227062 228217 227146 228453
rect 227382 228217 227414 228453
rect 226794 228133 227414 228217
rect 226794 227897 226826 228133
rect 227062 227897 227146 228133
rect 227382 227897 227414 228133
rect 226794 192454 227414 227897
rect 226794 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 227414 192454
rect 226794 192134 227414 192218
rect 226794 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 227414 192134
rect 226794 156454 227414 191898
rect 226794 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 227414 156454
rect 226794 156134 227414 156218
rect 226794 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 227414 156134
rect 226794 120454 227414 155898
rect 226794 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 227414 120454
rect 226794 120134 227414 120218
rect 226794 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 227414 120134
rect 226794 84454 227414 119898
rect 226794 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 227414 84454
rect 226794 84134 227414 84218
rect 226794 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 227414 84134
rect 226794 48454 227414 83898
rect 226794 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 227414 48454
rect 226794 48134 227414 48218
rect 226794 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 227414 48134
rect 226794 12454 227414 47898
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2266 227414 11898
rect 226794 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 227414 -2266
rect 226794 -2586 227414 -2502
rect 226794 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 227414 -2586
rect 226794 -7654 227414 -2822
rect 231294 196954 231914 228484
rect 231294 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 231914 196954
rect 231294 196634 231914 196718
rect 231294 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 231914 196634
rect 231294 160954 231914 196398
rect 231294 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 231914 160954
rect 231294 160634 231914 160718
rect 231294 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 231914 160634
rect 231294 124954 231914 160398
rect 231294 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 231914 124954
rect 231294 124634 231914 124718
rect 231294 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 231914 124634
rect 231294 88954 231914 124398
rect 231294 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 231914 88954
rect 231294 88634 231914 88718
rect 231294 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 231914 88634
rect 231294 52954 231914 88398
rect 231294 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 231914 52954
rect 231294 52634 231914 52718
rect 231294 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 231914 52634
rect 231294 16954 231914 52398
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3226 231914 16398
rect 231294 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 231914 -3226
rect 231294 -3546 231914 -3462
rect 231294 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 231914 -3546
rect 231294 -7654 231914 -3782
rect 235794 201454 236414 228484
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4186 236414 20898
rect 235794 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 236414 -4186
rect 235794 -4506 236414 -4422
rect 235794 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 236414 -4506
rect 235794 -7654 236414 -4742
rect 240294 205954 240914 228484
rect 240294 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 240914 205954
rect 240294 205634 240914 205718
rect 240294 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 240914 205634
rect 240294 169954 240914 205398
rect 240294 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 240914 169954
rect 240294 169634 240914 169718
rect 240294 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 240914 169634
rect 240294 133954 240914 169398
rect 240294 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 240914 133954
rect 240294 133634 240914 133718
rect 240294 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 240914 133634
rect 240294 97954 240914 133398
rect 240294 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 240914 97954
rect 240294 97634 240914 97718
rect 240294 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 240914 97634
rect 240294 61954 240914 97398
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 25954 240914 61398
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 240294 -5146 240914 25398
rect 240294 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 240914 -5146
rect 240294 -5466 240914 -5382
rect 240294 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 240914 -5466
rect 240294 -7654 240914 -5702
rect 244794 210454 245414 228484
rect 244794 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 245414 210454
rect 244794 210134 245414 210218
rect 244794 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 245414 210134
rect 244794 174454 245414 209898
rect 244794 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 245414 174454
rect 244794 174134 245414 174218
rect 244794 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 245414 174134
rect 244794 138454 245414 173898
rect 244794 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 245414 138454
rect 244794 138134 245414 138218
rect 244794 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 245414 138134
rect 244794 102454 245414 137898
rect 244794 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 245414 102454
rect 244794 102134 245414 102218
rect 244794 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 245414 102134
rect 244794 66454 245414 101898
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 30454 245414 65898
rect 244794 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 245414 30454
rect 244794 30134 245414 30218
rect 244794 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 245414 30134
rect 244794 -6106 245414 29898
rect 244794 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 245414 -6106
rect 244794 -6426 245414 -6342
rect 244794 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 245414 -6426
rect 244794 -7654 245414 -6662
rect 249294 214954 249914 228484
rect 249294 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 249914 214954
rect 249294 214634 249914 214718
rect 249294 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 249914 214634
rect 249294 178954 249914 214398
rect 249294 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 249914 178954
rect 249294 178634 249914 178718
rect 249294 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 249914 178634
rect 249294 142954 249914 178398
rect 249294 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 249914 142954
rect 249294 142634 249914 142718
rect 249294 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 249914 142634
rect 249294 106954 249914 142398
rect 249294 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 249914 106954
rect 249294 106634 249914 106718
rect 249294 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 249914 106634
rect 249294 70954 249914 106398
rect 249294 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 249914 70954
rect 249294 70634 249914 70718
rect 249294 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 249914 70634
rect 249294 34954 249914 70398
rect 249294 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 249914 34954
rect 249294 34634 249914 34718
rect 249294 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 249914 34634
rect 249294 -7066 249914 34398
rect 249294 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 249914 -7066
rect 249294 -7386 249914 -7302
rect 249294 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 249914 -7386
rect 249294 -7654 249914 -7622
rect 253794 219454 254414 228484
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 258294 223954 258914 228484
rect 258294 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 258914 223954
rect 258294 223634 258914 223718
rect 258294 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 258914 223634
rect 258294 187954 258914 223398
rect 258294 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 258914 187954
rect 258294 187634 258914 187718
rect 258294 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 258914 187634
rect 258294 151954 258914 187398
rect 258294 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 258914 151954
rect 258294 151634 258914 151718
rect 258294 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 258914 151634
rect 258294 115954 258914 151398
rect 258294 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 258914 115954
rect 258294 115634 258914 115718
rect 258294 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 258914 115634
rect 258294 79954 258914 115398
rect 258294 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 258914 79954
rect 258294 79634 258914 79718
rect 258294 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 258914 79634
rect 258294 43954 258914 79398
rect 258294 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 258914 43954
rect 258294 43634 258914 43718
rect 258294 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 258914 43634
rect 258294 7954 258914 43398
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258294 -1306 258914 7398
rect 258294 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 258914 -1306
rect 258294 -1626 258914 -1542
rect 258294 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 258914 -1626
rect 258294 -7654 258914 -1862
rect 262794 228453 263414 228484
rect 262794 228217 262826 228453
rect 263062 228217 263146 228453
rect 263382 228217 263414 228453
rect 262794 228133 263414 228217
rect 262794 227897 262826 228133
rect 263062 227897 263146 228133
rect 263382 227897 263414 228133
rect 262794 192454 263414 227897
rect 262794 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 263414 192454
rect 262794 192134 263414 192218
rect 262794 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 263414 192134
rect 262794 156454 263414 191898
rect 262794 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 263414 156454
rect 262794 156134 263414 156218
rect 262794 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 263414 156134
rect 262794 120454 263414 155898
rect 262794 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 263414 120454
rect 262794 120134 263414 120218
rect 262794 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 263414 120134
rect 262794 84454 263414 119898
rect 262794 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 263414 84454
rect 262794 84134 263414 84218
rect 262794 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 263414 84134
rect 262794 48454 263414 83898
rect 262794 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 263414 48454
rect 262794 48134 263414 48218
rect 262794 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 263414 48134
rect 262794 12454 263414 47898
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2266 263414 11898
rect 262794 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 263414 -2266
rect 262794 -2586 263414 -2502
rect 262794 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 263414 -2586
rect 262794 -7654 263414 -2822
rect 267294 196954 267914 228484
rect 267294 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 267914 196954
rect 267294 196634 267914 196718
rect 267294 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 267914 196634
rect 267294 160954 267914 196398
rect 267294 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 267914 160954
rect 267294 160634 267914 160718
rect 267294 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 267914 160634
rect 267294 124954 267914 160398
rect 267294 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 267914 124954
rect 267294 124634 267914 124718
rect 267294 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 267914 124634
rect 267294 88954 267914 124398
rect 267294 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 267914 88954
rect 267294 88634 267914 88718
rect 267294 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 267914 88634
rect 267294 52954 267914 88398
rect 267294 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 267914 52954
rect 267294 52634 267914 52718
rect 267294 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 267914 52634
rect 267294 16954 267914 52398
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3226 267914 16398
rect 267294 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 267914 -3226
rect 267294 -3546 267914 -3462
rect 267294 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 267914 -3546
rect 267294 -7654 267914 -3782
rect 271794 201454 272414 228484
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4186 272414 20898
rect 271794 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 272414 -4186
rect 271794 -4506 272414 -4422
rect 271794 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 272414 -4506
rect 271794 -7654 272414 -4742
rect 276294 205954 276914 228484
rect 276294 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 276914 205954
rect 276294 205634 276914 205718
rect 276294 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 276914 205634
rect 276294 169954 276914 205398
rect 276294 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 276914 169954
rect 276294 169634 276914 169718
rect 276294 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 276914 169634
rect 276294 133954 276914 169398
rect 276294 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 276914 133954
rect 276294 133634 276914 133718
rect 276294 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 276914 133634
rect 276294 97954 276914 133398
rect 276294 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 276914 97954
rect 276294 97634 276914 97718
rect 276294 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 276914 97634
rect 276294 61954 276914 97398
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 25954 276914 61398
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 276294 -5146 276914 25398
rect 276294 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 276914 -5146
rect 276294 -5466 276914 -5382
rect 276294 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 276914 -5466
rect 276294 -7654 276914 -5702
rect 280794 210454 281414 228484
rect 280794 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 281414 210454
rect 280794 210134 281414 210218
rect 280794 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 281414 210134
rect 280794 174454 281414 209898
rect 280794 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 281414 174454
rect 280794 174134 281414 174218
rect 280794 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 281414 174134
rect 280794 138454 281414 173898
rect 280794 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 281414 138454
rect 280794 138134 281414 138218
rect 280794 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 281414 138134
rect 280794 102454 281414 137898
rect 280794 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 281414 102454
rect 280794 102134 281414 102218
rect 280794 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 281414 102134
rect 280794 66454 281414 101898
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 30454 281414 65898
rect 280794 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 281414 30454
rect 280794 30134 281414 30218
rect 280794 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 281414 30134
rect 280794 -6106 281414 29898
rect 280794 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 281414 -6106
rect 280794 -6426 281414 -6342
rect 280794 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 281414 -6426
rect 280794 -7654 281414 -6662
rect 285294 214954 285914 228484
rect 285294 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 285914 214954
rect 285294 214634 285914 214718
rect 285294 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 285914 214634
rect 285294 178954 285914 214398
rect 285294 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 285914 178954
rect 285294 178634 285914 178718
rect 285294 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 285914 178634
rect 285294 142954 285914 178398
rect 285294 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 285914 142954
rect 285294 142634 285914 142718
rect 285294 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 285914 142634
rect 285294 106954 285914 142398
rect 285294 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 285914 106954
rect 285294 106634 285914 106718
rect 285294 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 285914 106634
rect 285294 70954 285914 106398
rect 285294 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 285914 70954
rect 285294 70634 285914 70718
rect 285294 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 285914 70634
rect 285294 34954 285914 70398
rect 285294 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 285914 34954
rect 285294 34634 285914 34718
rect 285294 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 285914 34634
rect 285294 -7066 285914 34398
rect 285294 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 285914 -7066
rect 285294 -7386 285914 -7302
rect 285294 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 285914 -7386
rect 285294 -7654 285914 -7622
rect 289794 219454 290414 228484
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 294294 223954 294914 228484
rect 294294 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 294914 223954
rect 294294 223634 294914 223718
rect 294294 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 294914 223634
rect 294294 187954 294914 223398
rect 294294 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 294914 187954
rect 294294 187634 294914 187718
rect 294294 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 294914 187634
rect 294294 151954 294914 187398
rect 294294 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 294914 151954
rect 294294 151634 294914 151718
rect 294294 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 294914 151634
rect 294294 115954 294914 151398
rect 294294 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 294914 115954
rect 294294 115634 294914 115718
rect 294294 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 294914 115634
rect 294294 79954 294914 115398
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 294294 43954 294914 79398
rect 294294 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 294914 43954
rect 294294 43634 294914 43718
rect 294294 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 294914 43634
rect 294294 7954 294914 43398
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1306 294914 7398
rect 294294 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 294914 -1306
rect 294294 -1626 294914 -1542
rect 294294 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 294914 -1626
rect 294294 -7654 294914 -1862
rect 298794 228453 299414 228484
rect 298794 228217 298826 228453
rect 299062 228217 299146 228453
rect 299382 228217 299414 228453
rect 298794 228133 299414 228217
rect 298794 227897 298826 228133
rect 299062 227897 299146 228133
rect 299382 227897 299414 228133
rect 298794 192454 299414 227897
rect 298794 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 299414 192454
rect 298794 192134 299414 192218
rect 298794 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 299414 192134
rect 298794 156454 299414 191898
rect 298794 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 299414 156454
rect 298794 156134 299414 156218
rect 298794 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 299414 156134
rect 298794 120454 299414 155898
rect 298794 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 299414 120454
rect 298794 120134 299414 120218
rect 298794 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 299414 120134
rect 298794 84454 299414 119898
rect 298794 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 299414 84454
rect 298794 84134 299414 84218
rect 298794 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 299414 84134
rect 298794 48454 299414 83898
rect 298794 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 299414 48454
rect 298794 48134 299414 48218
rect 298794 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 299414 48134
rect 298794 12454 299414 47898
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298794 -2266 299414 11898
rect 298794 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 299414 -2266
rect 298794 -2586 299414 -2502
rect 298794 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 299414 -2586
rect 298794 -7654 299414 -2822
rect 303294 196954 303914 228484
rect 303294 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 303914 196954
rect 303294 196634 303914 196718
rect 303294 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 303914 196634
rect 303294 160954 303914 196398
rect 303294 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 303914 160954
rect 303294 160634 303914 160718
rect 303294 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 303914 160634
rect 303294 124954 303914 160398
rect 303294 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 303914 124954
rect 303294 124634 303914 124718
rect 303294 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 303914 124634
rect 303294 88954 303914 124398
rect 303294 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 303914 88954
rect 303294 88634 303914 88718
rect 303294 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 303914 88634
rect 303294 52954 303914 88398
rect 303294 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 303914 52954
rect 303294 52634 303914 52718
rect 303294 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 303914 52634
rect 303294 16954 303914 52398
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 303294 -3226 303914 16398
rect 303294 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 303914 -3226
rect 303294 -3546 303914 -3462
rect 303294 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 303914 -3546
rect 303294 -7654 303914 -3782
rect 307794 201454 308414 228484
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4186 308414 20898
rect 307794 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 308414 -4186
rect 307794 -4506 308414 -4422
rect 307794 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 308414 -4506
rect 307794 -7654 308414 -4742
rect 312294 205954 312914 228484
rect 312294 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 312914 205954
rect 312294 205634 312914 205718
rect 312294 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 312914 205634
rect 312294 169954 312914 205398
rect 312294 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 312914 169954
rect 312294 169634 312914 169718
rect 312294 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 312914 169634
rect 312294 133954 312914 169398
rect 312294 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 312914 133954
rect 312294 133634 312914 133718
rect 312294 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 312914 133634
rect 312294 97954 312914 133398
rect 312294 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 312914 97954
rect 312294 97634 312914 97718
rect 312294 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 312914 97634
rect 312294 61954 312914 97398
rect 312294 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 312914 61954
rect 312294 61634 312914 61718
rect 312294 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 312914 61634
rect 312294 25954 312914 61398
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 312294 -5146 312914 25398
rect 312294 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 312914 -5146
rect 312294 -5466 312914 -5382
rect 312294 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 312914 -5466
rect 312294 -7654 312914 -5702
rect 316794 210454 317414 228484
rect 316794 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 317414 210454
rect 316794 210134 317414 210218
rect 316794 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 317414 210134
rect 316794 174454 317414 209898
rect 316794 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 317414 174454
rect 316794 174134 317414 174218
rect 316794 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 317414 174134
rect 316794 138454 317414 173898
rect 316794 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 317414 138454
rect 316794 138134 317414 138218
rect 316794 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 317414 138134
rect 316794 102454 317414 137898
rect 316794 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 317414 102454
rect 316794 102134 317414 102218
rect 316794 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 317414 102134
rect 316794 66454 317414 101898
rect 316794 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 317414 66454
rect 316794 66134 317414 66218
rect 316794 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 317414 66134
rect 316794 30454 317414 65898
rect 316794 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 317414 30454
rect 316794 30134 317414 30218
rect 316794 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 317414 30134
rect 316794 -6106 317414 29898
rect 316794 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 317414 -6106
rect 316794 -6426 317414 -6342
rect 316794 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 317414 -6426
rect 316794 -7654 317414 -6662
rect 321294 214954 321914 228484
rect 321294 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 321914 214954
rect 321294 214634 321914 214718
rect 321294 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 321914 214634
rect 321294 178954 321914 214398
rect 321294 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 321914 178954
rect 321294 178634 321914 178718
rect 321294 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 321914 178634
rect 321294 142954 321914 178398
rect 321294 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 321914 142954
rect 321294 142634 321914 142718
rect 321294 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 321914 142634
rect 321294 106954 321914 142398
rect 321294 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 321914 106954
rect 321294 106634 321914 106718
rect 321294 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 321914 106634
rect 321294 70954 321914 106398
rect 321294 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 321914 70954
rect 321294 70634 321914 70718
rect 321294 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 321914 70634
rect 321294 34954 321914 70398
rect 321294 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 321914 34954
rect 321294 34634 321914 34718
rect 321294 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 321914 34634
rect 321294 -7066 321914 34398
rect 321294 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 321914 -7066
rect 321294 -7386 321914 -7302
rect 321294 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 321914 -7386
rect 321294 -7654 321914 -7622
rect 325794 219454 326414 228484
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 330294 223954 330914 228484
rect 330294 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 330914 223954
rect 330294 223634 330914 223718
rect 330294 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 330914 223634
rect 330294 187954 330914 223398
rect 330294 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 330914 187954
rect 330294 187634 330914 187718
rect 330294 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 330914 187634
rect 330294 151954 330914 187398
rect 330294 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 330914 151954
rect 330294 151634 330914 151718
rect 330294 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 330914 151634
rect 330294 115954 330914 151398
rect 330294 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 330914 115954
rect 330294 115634 330914 115718
rect 330294 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 330914 115634
rect 330294 79954 330914 115398
rect 330294 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 330914 79954
rect 330294 79634 330914 79718
rect 330294 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 330914 79634
rect 330294 43954 330914 79398
rect 330294 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 330914 43954
rect 330294 43634 330914 43718
rect 330294 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 330914 43634
rect 330294 7954 330914 43398
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1306 330914 7398
rect 330294 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 330914 -1306
rect 330294 -1626 330914 -1542
rect 330294 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 330914 -1626
rect 330294 -7654 330914 -1862
rect 334794 228453 335414 228484
rect 334794 228217 334826 228453
rect 335062 228217 335146 228453
rect 335382 228217 335414 228453
rect 334794 228133 335414 228217
rect 334794 227897 334826 228133
rect 335062 227897 335146 228133
rect 335382 227897 335414 228133
rect 334794 192454 335414 227897
rect 334794 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 335414 192454
rect 334794 192134 335414 192218
rect 334794 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 335414 192134
rect 334794 156454 335414 191898
rect 334794 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 335414 156454
rect 334794 156134 335414 156218
rect 334794 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 335414 156134
rect 334794 120454 335414 155898
rect 334794 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 335414 120454
rect 334794 120134 335414 120218
rect 334794 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 335414 120134
rect 334794 84454 335414 119898
rect 334794 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 335414 84454
rect 334794 84134 335414 84218
rect 334794 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 335414 84134
rect 334794 48454 335414 83898
rect 334794 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 335414 48454
rect 334794 48134 335414 48218
rect 334794 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 335414 48134
rect 334794 12454 335414 47898
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2266 335414 11898
rect 334794 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 335414 -2266
rect 334794 -2586 335414 -2502
rect 334794 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 335414 -2586
rect 334794 -7654 335414 -2822
rect 339294 196954 339914 228484
rect 339294 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 339914 196954
rect 339294 196634 339914 196718
rect 339294 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 339914 196634
rect 339294 160954 339914 196398
rect 339294 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 339914 160954
rect 339294 160634 339914 160718
rect 339294 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 339914 160634
rect 339294 124954 339914 160398
rect 339294 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 339914 124954
rect 339294 124634 339914 124718
rect 339294 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 339914 124634
rect 339294 88954 339914 124398
rect 339294 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 339914 88954
rect 339294 88634 339914 88718
rect 339294 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 339914 88634
rect 339294 52954 339914 88398
rect 339294 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 339914 52954
rect 339294 52634 339914 52718
rect 339294 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 339914 52634
rect 339294 16954 339914 52398
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3226 339914 16398
rect 339294 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 339914 -3226
rect 339294 -3546 339914 -3462
rect 339294 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 339914 -3546
rect 339294 -7654 339914 -3782
rect 343794 201454 344414 228484
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -4186 344414 20898
rect 343794 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 344414 -4186
rect 343794 -4506 344414 -4422
rect 343794 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 344414 -4506
rect 343794 -7654 344414 -4742
rect 348294 205954 348914 228484
rect 348294 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 348914 205954
rect 348294 205634 348914 205718
rect 348294 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 348914 205634
rect 348294 169954 348914 205398
rect 348294 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 348914 169954
rect 348294 169634 348914 169718
rect 348294 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 348914 169634
rect 348294 133954 348914 169398
rect 348294 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 348914 133954
rect 348294 133634 348914 133718
rect 348294 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 348914 133634
rect 348294 97954 348914 133398
rect 348294 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 348914 97954
rect 348294 97634 348914 97718
rect 348294 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 348914 97634
rect 348294 61954 348914 97398
rect 348294 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 348914 61954
rect 348294 61634 348914 61718
rect 348294 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 348914 61634
rect 348294 25954 348914 61398
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 348294 -5146 348914 25398
rect 348294 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 348914 -5146
rect 348294 -5466 348914 -5382
rect 348294 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 348914 -5466
rect 348294 -7654 348914 -5702
rect 352794 210454 353414 228484
rect 352794 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 353414 210454
rect 352794 210134 353414 210218
rect 352794 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 353414 210134
rect 352794 174454 353414 209898
rect 352794 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 353414 174454
rect 352794 174134 353414 174218
rect 352794 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 353414 174134
rect 352794 138454 353414 173898
rect 352794 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 353414 138454
rect 352794 138134 353414 138218
rect 352794 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 353414 138134
rect 352794 102454 353414 137898
rect 352794 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 353414 102454
rect 352794 102134 353414 102218
rect 352794 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 353414 102134
rect 352794 66454 353414 101898
rect 352794 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 353414 66454
rect 352794 66134 353414 66218
rect 352794 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 353414 66134
rect 352794 30454 353414 65898
rect 352794 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 353414 30454
rect 352794 30134 353414 30218
rect 352794 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 353414 30134
rect 352794 -6106 353414 29898
rect 352794 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 353414 -6106
rect 352794 -6426 353414 -6342
rect 352794 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 353414 -6426
rect 352794 -7654 353414 -6662
rect 357294 214954 357914 228484
rect 357294 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 357914 214954
rect 357294 214634 357914 214718
rect 357294 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 357914 214634
rect 357294 178954 357914 214398
rect 357294 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 357914 178954
rect 357294 178634 357914 178718
rect 357294 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 357914 178634
rect 357294 142954 357914 178398
rect 357294 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 357914 142954
rect 357294 142634 357914 142718
rect 357294 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 357914 142634
rect 357294 106954 357914 142398
rect 357294 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 357914 106954
rect 357294 106634 357914 106718
rect 357294 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 357914 106634
rect 357294 70954 357914 106398
rect 357294 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 357914 70954
rect 357294 70634 357914 70718
rect 357294 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 357914 70634
rect 357294 34954 357914 70398
rect 357294 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 357914 34954
rect 357294 34634 357914 34718
rect 357294 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 357914 34634
rect 357294 -7066 357914 34398
rect 357294 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 357914 -7066
rect 357294 -7386 357914 -7302
rect 357294 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 357914 -7386
rect 357294 -7654 357914 -7622
rect 361794 219454 362414 228484
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 366294 223954 366914 228484
rect 366294 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 366914 223954
rect 366294 223634 366914 223718
rect 366294 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 366914 223634
rect 366294 187954 366914 223398
rect 366294 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 366914 187954
rect 366294 187634 366914 187718
rect 366294 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 366914 187634
rect 366294 151954 366914 187398
rect 366294 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 366914 151954
rect 366294 151634 366914 151718
rect 366294 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 366914 151634
rect 366294 115954 366914 151398
rect 366294 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 366914 115954
rect 366294 115634 366914 115718
rect 366294 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 366914 115634
rect 366294 79954 366914 115398
rect 366294 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 366914 79954
rect 366294 79634 366914 79718
rect 366294 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 366914 79634
rect 366294 43954 366914 79398
rect 366294 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 366914 43954
rect 366294 43634 366914 43718
rect 366294 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 366914 43634
rect 366294 7954 366914 43398
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 366294 -1306 366914 7398
rect 366294 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 366914 -1306
rect 366294 -1626 366914 -1542
rect 366294 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 366914 -1626
rect 366294 -7654 366914 -1862
rect 370794 228453 371414 228484
rect 370794 228217 370826 228453
rect 371062 228217 371146 228453
rect 371382 228217 371414 228453
rect 370794 228133 371414 228217
rect 370794 227897 370826 228133
rect 371062 227897 371146 228133
rect 371382 227897 371414 228133
rect 370794 192454 371414 227897
rect 370794 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 371414 192454
rect 370794 192134 371414 192218
rect 370794 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 371414 192134
rect 370794 156454 371414 191898
rect 370794 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 371414 156454
rect 370794 156134 371414 156218
rect 370794 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 371414 156134
rect 370794 120454 371414 155898
rect 370794 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 371414 120454
rect 370794 120134 371414 120218
rect 370794 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 371414 120134
rect 370794 84454 371414 119898
rect 370794 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 371414 84454
rect 370794 84134 371414 84218
rect 370794 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 371414 84134
rect 370794 48454 371414 83898
rect 370794 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 371414 48454
rect 370794 48134 371414 48218
rect 370794 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 371414 48134
rect 370794 12454 371414 47898
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -2266 371414 11898
rect 370794 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 371414 -2266
rect 370794 -2586 371414 -2502
rect 370794 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 371414 -2586
rect 370794 -7654 371414 -2822
rect 375294 196954 375914 228484
rect 375294 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 375914 196954
rect 375294 196634 375914 196718
rect 375294 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 375914 196634
rect 375294 160954 375914 196398
rect 375294 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 375914 160954
rect 375294 160634 375914 160718
rect 375294 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 375914 160634
rect 375294 124954 375914 160398
rect 375294 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 375914 124954
rect 375294 124634 375914 124718
rect 375294 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 375914 124634
rect 375294 88954 375914 124398
rect 375294 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 375914 88954
rect 375294 88634 375914 88718
rect 375294 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 375914 88634
rect 375294 52954 375914 88398
rect 375294 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 375914 52954
rect 375294 52634 375914 52718
rect 375294 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 375914 52634
rect 375294 16954 375914 52398
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3226 375914 16398
rect 375294 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 375914 -3226
rect 375294 -3546 375914 -3462
rect 375294 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 375914 -3546
rect 375294 -7654 375914 -3782
rect 379794 201454 380414 228484
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4186 380414 20898
rect 379794 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 380414 -4186
rect 379794 -4506 380414 -4422
rect 379794 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 380414 -4506
rect 379794 -7654 380414 -4742
rect 384294 205954 384914 228484
rect 384294 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 384914 205954
rect 384294 205634 384914 205718
rect 384294 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 384914 205634
rect 384294 169954 384914 205398
rect 384294 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 384914 169954
rect 384294 169634 384914 169718
rect 384294 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 384914 169634
rect 384294 133954 384914 169398
rect 384294 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 384914 133954
rect 384294 133634 384914 133718
rect 384294 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 384914 133634
rect 384294 97954 384914 133398
rect 384294 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 384914 97954
rect 384294 97634 384914 97718
rect 384294 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 384914 97634
rect 384294 61954 384914 97398
rect 384294 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 384914 61954
rect 384294 61634 384914 61718
rect 384294 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 384914 61634
rect 384294 25954 384914 61398
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5146 384914 25398
rect 384294 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 384914 -5146
rect 384294 -5466 384914 -5382
rect 384294 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 384914 -5466
rect 384294 -7654 384914 -5702
rect 388794 210454 389414 228484
rect 388794 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 389414 210454
rect 388794 210134 389414 210218
rect 388794 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 389414 210134
rect 388794 174454 389414 209898
rect 388794 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 389414 174454
rect 388794 174134 389414 174218
rect 388794 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 389414 174134
rect 388794 138454 389414 173898
rect 388794 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 389414 138454
rect 388794 138134 389414 138218
rect 388794 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 389414 138134
rect 388794 102454 389414 137898
rect 388794 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 389414 102454
rect 388794 102134 389414 102218
rect 388794 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 389414 102134
rect 388794 66454 389414 101898
rect 388794 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 389414 66454
rect 388794 66134 389414 66218
rect 388794 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 389414 66134
rect 388794 30454 389414 65898
rect 388794 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 389414 30454
rect 388794 30134 389414 30218
rect 388794 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 389414 30134
rect 388794 -6106 389414 29898
rect 388794 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 389414 -6106
rect 388794 -6426 389414 -6342
rect 388794 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 389414 -6426
rect 388794 -7654 389414 -6662
rect 393294 214954 393914 228484
rect 393294 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 393914 214954
rect 393294 214634 393914 214718
rect 393294 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 393914 214634
rect 393294 178954 393914 214398
rect 393294 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 393914 178954
rect 393294 178634 393914 178718
rect 393294 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 393914 178634
rect 393294 142954 393914 178398
rect 393294 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 393914 142954
rect 393294 142634 393914 142718
rect 393294 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 393914 142634
rect 393294 106954 393914 142398
rect 393294 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 393914 106954
rect 393294 106634 393914 106718
rect 393294 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 393914 106634
rect 393294 70954 393914 106398
rect 396582 78165 396642 696899
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 396763 643244 396829 643245
rect 396763 643180 396764 643244
rect 396828 643180 396829 643244
rect 396763 643179 396829 643180
rect 396766 78437 396826 643179
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 248684 398414 254898
rect 402294 705798 402914 711590
rect 402294 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 402914 705798
rect 402294 705478 402914 705562
rect 402294 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 402914 705478
rect 402294 691954 402914 705242
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 402294 655954 402914 691398
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402294 619954 402914 655398
rect 402294 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 402914 619954
rect 402294 619634 402914 619718
rect 402294 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 402914 619634
rect 402294 583954 402914 619398
rect 402294 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 402914 583954
rect 402294 583634 402914 583718
rect 402294 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 402914 583634
rect 402294 547954 402914 583398
rect 402294 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 402914 547954
rect 402294 547634 402914 547718
rect 402294 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 402914 547634
rect 402294 511954 402914 547398
rect 402294 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 402914 511954
rect 402294 511634 402914 511718
rect 402294 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 402914 511634
rect 402294 475954 402914 511398
rect 402294 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 402914 475954
rect 402294 475634 402914 475718
rect 402294 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 402914 475634
rect 402294 439954 402914 475398
rect 402294 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 402914 439954
rect 402294 439634 402914 439718
rect 402294 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 402914 439634
rect 402294 403954 402914 439398
rect 402294 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 402914 403954
rect 402294 403634 402914 403718
rect 402294 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 402914 403634
rect 402294 367954 402914 403398
rect 402294 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 402914 367954
rect 402294 367634 402914 367718
rect 402294 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 402914 367634
rect 402294 331954 402914 367398
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 295954 402914 331398
rect 402294 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 402914 295954
rect 402294 295634 402914 295718
rect 402294 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 402914 295634
rect 402294 259954 402914 295398
rect 402294 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 402914 259954
rect 402294 259634 402914 259718
rect 402294 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 402914 259634
rect 397794 219454 398414 228484
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 396763 78436 396829 78437
rect 396763 78372 396764 78436
rect 396828 78372 396829 78436
rect 396763 78371 396829 78372
rect 396579 78164 396645 78165
rect 396579 78100 396580 78164
rect 396644 78100 396645 78164
rect 396579 78099 396645 78100
rect 393294 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 393914 70954
rect 393294 70634 393914 70718
rect 393294 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 393914 70634
rect 393294 34954 393914 70398
rect 393294 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 393914 34954
rect 393294 34634 393914 34718
rect 393294 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 393914 34634
rect 393294 -7066 393914 34398
rect 393294 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 393914 -7066
rect 393294 -7386 393914 -7302
rect 393294 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 393914 -7386
rect 393294 -7654 393914 -7622
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 402294 223954 402914 259398
rect 402294 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 402914 223954
rect 402294 223634 402914 223718
rect 402294 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 402914 223634
rect 402294 187954 402914 223398
rect 402294 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 402914 187954
rect 402294 187634 402914 187718
rect 402294 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 402914 187634
rect 402294 151954 402914 187398
rect 402294 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 402914 151954
rect 402294 151634 402914 151718
rect 402294 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 402914 151634
rect 402294 115954 402914 151398
rect 402294 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 402914 115954
rect 402294 115634 402914 115718
rect 402294 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 402914 115634
rect 402294 79954 402914 115398
rect 402294 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 402914 79954
rect 402294 79634 402914 79718
rect 402294 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 402914 79634
rect 402294 43954 402914 79398
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1306 402914 7398
rect 402294 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 402914 -1306
rect 402294 -1626 402914 -1542
rect 402294 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 402914 -1626
rect 402294 -7654 402914 -1862
rect 406794 706758 407414 711590
rect 406794 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 407414 706758
rect 406794 706438 407414 706522
rect 406794 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 407414 706438
rect 406794 696454 407414 706202
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 406794 660454 407414 695898
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 624454 407414 659898
rect 406794 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 407414 624454
rect 406794 624134 407414 624218
rect 406794 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 407414 624134
rect 406794 588454 407414 623898
rect 406794 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 407414 588454
rect 406794 588134 407414 588218
rect 406794 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 407414 588134
rect 406794 552454 407414 587898
rect 406794 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 407414 552454
rect 406794 552134 407414 552218
rect 406794 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 407414 552134
rect 406794 516454 407414 551898
rect 406794 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 407414 516454
rect 406794 516134 407414 516218
rect 406794 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 407414 516134
rect 406794 480454 407414 515898
rect 406794 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 407414 480454
rect 406794 480134 407414 480218
rect 406794 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 407414 480134
rect 406794 444454 407414 479898
rect 406794 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 407414 444454
rect 406794 444134 407414 444218
rect 406794 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 407414 444134
rect 406794 408454 407414 443898
rect 406794 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 407414 408454
rect 406794 408134 407414 408218
rect 406794 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 407414 408134
rect 406794 372454 407414 407898
rect 406794 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 407414 372454
rect 406794 372134 407414 372218
rect 406794 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 407414 372134
rect 406794 336454 407414 371898
rect 406794 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 407414 336454
rect 406794 336134 407414 336218
rect 406794 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 407414 336134
rect 406794 300454 407414 335898
rect 406794 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 407414 300454
rect 406794 300134 407414 300218
rect 406794 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 407414 300134
rect 406794 264454 407414 299898
rect 406794 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 407414 264454
rect 406794 264134 407414 264218
rect 406794 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 407414 264134
rect 406794 228454 407414 263898
rect 406794 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 407414 228454
rect 406794 228134 407414 228218
rect 406794 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 407414 228134
rect 406794 192454 407414 227898
rect 406794 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 407414 192454
rect 406794 192134 407414 192218
rect 406794 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 407414 192134
rect 406794 156454 407414 191898
rect 406794 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 407414 156454
rect 406794 156134 407414 156218
rect 406794 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 407414 156134
rect 406794 120454 407414 155898
rect 406794 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 407414 120454
rect 406794 120134 407414 120218
rect 406794 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 407414 120134
rect 406794 84454 407414 119898
rect 406794 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 407414 84454
rect 406794 84134 407414 84218
rect 406794 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 407414 84134
rect 406794 48454 407414 83898
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2266 407414 11898
rect 406794 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 407414 -2266
rect 406794 -2586 407414 -2502
rect 406794 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 407414 -2586
rect 406794 -7654 407414 -2822
rect 411294 707718 411914 711590
rect 411294 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 411914 707718
rect 411294 707398 411914 707482
rect 411294 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 411914 707398
rect 411294 700954 411914 707162
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 664954 411914 700398
rect 411294 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 411914 664954
rect 411294 664634 411914 664718
rect 411294 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 411914 664634
rect 411294 628954 411914 664398
rect 411294 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 411914 628954
rect 411294 628634 411914 628718
rect 411294 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 411914 628634
rect 411294 592954 411914 628398
rect 411294 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 411914 592954
rect 411294 592634 411914 592718
rect 411294 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 411914 592634
rect 411294 556954 411914 592398
rect 411294 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 411914 556954
rect 411294 556634 411914 556718
rect 411294 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 411914 556634
rect 411294 520954 411914 556398
rect 411294 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 411914 520954
rect 411294 520634 411914 520718
rect 411294 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 411914 520634
rect 411294 484954 411914 520398
rect 411294 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 411914 484954
rect 411294 484634 411914 484718
rect 411294 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 411914 484634
rect 411294 448954 411914 484398
rect 411294 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 411914 448954
rect 411294 448634 411914 448718
rect 411294 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 411914 448634
rect 411294 412954 411914 448398
rect 411294 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 411914 412954
rect 411294 412634 411914 412718
rect 411294 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 411914 412634
rect 411294 376954 411914 412398
rect 411294 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 411914 376954
rect 411294 376634 411914 376718
rect 411294 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 411914 376634
rect 411294 340954 411914 376398
rect 411294 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 411914 340954
rect 411294 340634 411914 340718
rect 411294 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 411914 340634
rect 411294 304954 411914 340398
rect 411294 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 411914 304954
rect 411294 304634 411914 304718
rect 411294 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 411914 304634
rect 411294 268954 411914 304398
rect 411294 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 411914 268954
rect 411294 268634 411914 268718
rect 411294 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 411914 268634
rect 411294 232954 411914 268398
rect 411294 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 411914 232954
rect 411294 232634 411914 232718
rect 411294 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 411914 232634
rect 411294 196954 411914 232398
rect 411294 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 411914 196954
rect 411294 196634 411914 196718
rect 411294 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 411914 196634
rect 411294 160954 411914 196398
rect 411294 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 411914 160954
rect 411294 160634 411914 160718
rect 411294 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 411914 160634
rect 411294 124954 411914 160398
rect 411294 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 411914 124954
rect 411294 124634 411914 124718
rect 411294 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 411914 124634
rect 411294 88954 411914 124398
rect 411294 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 411914 88954
rect 411294 88634 411914 88718
rect 411294 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 411914 88634
rect 411294 52954 411914 88398
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3226 411914 16398
rect 411294 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 411914 -3226
rect 411294 -3546 411914 -3462
rect 411294 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 411914 -3546
rect 411294 -7654 411914 -3782
rect 415794 708678 416414 711590
rect 415794 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 416414 708678
rect 415794 708358 416414 708442
rect 415794 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 416414 708358
rect 415794 669454 416414 708122
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4186 416414 20898
rect 415794 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 416414 -4186
rect 415794 -4506 416414 -4422
rect 415794 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 416414 -4506
rect 415794 -7654 416414 -4742
rect 420294 709638 420914 711590
rect 420294 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 420914 709638
rect 420294 709318 420914 709402
rect 420294 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 420914 709318
rect 420294 673954 420914 709082
rect 420294 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 420914 673954
rect 420294 673634 420914 673718
rect 420294 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 420914 673634
rect 420294 637954 420914 673398
rect 420294 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 420914 637954
rect 420294 637634 420914 637718
rect 420294 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 420914 637634
rect 420294 601954 420914 637398
rect 420294 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 420914 601954
rect 420294 601634 420914 601718
rect 420294 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 420914 601634
rect 420294 565954 420914 601398
rect 420294 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 420914 565954
rect 420294 565634 420914 565718
rect 420294 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 420914 565634
rect 420294 529954 420914 565398
rect 420294 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 420914 529954
rect 420294 529634 420914 529718
rect 420294 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 420914 529634
rect 420294 493954 420914 529398
rect 420294 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 420914 493954
rect 420294 493634 420914 493718
rect 420294 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 420914 493634
rect 420294 457954 420914 493398
rect 420294 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 420914 457954
rect 420294 457634 420914 457718
rect 420294 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 420914 457634
rect 420294 421954 420914 457398
rect 420294 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 420914 421954
rect 420294 421634 420914 421718
rect 420294 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 420914 421634
rect 420294 385954 420914 421398
rect 420294 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 420914 385954
rect 420294 385634 420914 385718
rect 420294 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 420914 385634
rect 420294 349954 420914 385398
rect 420294 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 420914 349954
rect 420294 349634 420914 349718
rect 420294 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 420914 349634
rect 420294 313954 420914 349398
rect 420294 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 420914 313954
rect 420294 313634 420914 313718
rect 420294 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 420914 313634
rect 420294 277954 420914 313398
rect 420294 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 420914 277954
rect 420294 277634 420914 277718
rect 420294 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 420914 277634
rect 420294 241954 420914 277398
rect 420294 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 420914 241954
rect 420294 241634 420914 241718
rect 420294 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 420914 241634
rect 420294 205954 420914 241398
rect 420294 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 420914 205954
rect 420294 205634 420914 205718
rect 420294 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 420914 205634
rect 420294 169954 420914 205398
rect 420294 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 420914 169954
rect 420294 169634 420914 169718
rect 420294 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 420914 169634
rect 420294 133954 420914 169398
rect 420294 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 420914 133954
rect 420294 133634 420914 133718
rect 420294 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 420914 133634
rect 420294 97954 420914 133398
rect 420294 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 420914 97954
rect 420294 97634 420914 97718
rect 420294 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 420914 97634
rect 420294 61954 420914 97398
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5146 420914 25398
rect 420294 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 420914 -5146
rect 420294 -5466 420914 -5382
rect 420294 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 420914 -5466
rect 420294 -7654 420914 -5702
rect 424794 710598 425414 711590
rect 424794 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 425414 710598
rect 424794 710278 425414 710362
rect 424794 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 425414 710278
rect 424794 678454 425414 710042
rect 424794 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 425414 678454
rect 424794 678134 425414 678218
rect 424794 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 425414 678134
rect 424794 642454 425414 677898
rect 424794 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 425414 642454
rect 424794 642134 425414 642218
rect 424794 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 425414 642134
rect 424794 606454 425414 641898
rect 424794 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 425414 606454
rect 424794 606134 425414 606218
rect 424794 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 425414 606134
rect 424794 570454 425414 605898
rect 424794 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 425414 570454
rect 424794 570134 425414 570218
rect 424794 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 425414 570134
rect 424794 534454 425414 569898
rect 424794 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 425414 534454
rect 424794 534134 425414 534218
rect 424794 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 425414 534134
rect 424794 498454 425414 533898
rect 424794 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 425414 498454
rect 424794 498134 425414 498218
rect 424794 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 425414 498134
rect 424794 462454 425414 497898
rect 424794 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 425414 462454
rect 424794 462134 425414 462218
rect 424794 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 425414 462134
rect 424794 426454 425414 461898
rect 424794 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 425414 426454
rect 424794 426134 425414 426218
rect 424794 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 425414 426134
rect 424794 390454 425414 425898
rect 424794 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 425414 390454
rect 424794 390134 425414 390218
rect 424794 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 425414 390134
rect 424794 354454 425414 389898
rect 424794 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 425414 354454
rect 424794 354134 425414 354218
rect 424794 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 425414 354134
rect 424794 318454 425414 353898
rect 424794 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 425414 318454
rect 424794 318134 425414 318218
rect 424794 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 425414 318134
rect 424794 282454 425414 317898
rect 424794 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 425414 282454
rect 424794 282134 425414 282218
rect 424794 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 425414 282134
rect 424794 246454 425414 281898
rect 424794 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 425414 246454
rect 424794 246134 425414 246218
rect 424794 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 425414 246134
rect 424794 210454 425414 245898
rect 424794 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 425414 210454
rect 424794 210134 425414 210218
rect 424794 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 425414 210134
rect 424794 174454 425414 209898
rect 424794 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 425414 174454
rect 424794 174134 425414 174218
rect 424794 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 425414 174134
rect 424794 138454 425414 173898
rect 424794 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 425414 138454
rect 424794 138134 425414 138218
rect 424794 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 425414 138134
rect 424794 102454 425414 137898
rect 424794 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 425414 102454
rect 424794 102134 425414 102218
rect 424794 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 425414 102134
rect 424794 66454 425414 101898
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6106 425414 29898
rect 424794 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 425414 -6106
rect 424794 -6426 425414 -6342
rect 424794 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 425414 -6426
rect 424794 -7654 425414 -6662
rect 429294 711558 429914 711590
rect 429294 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 429914 711558
rect 429294 711238 429914 711322
rect 429294 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 429914 711238
rect 429294 682954 429914 711002
rect 429294 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 429914 682954
rect 429294 682634 429914 682718
rect 429294 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 429914 682634
rect 429294 646954 429914 682398
rect 429294 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 429914 646954
rect 429294 646634 429914 646718
rect 429294 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 429914 646634
rect 429294 610954 429914 646398
rect 429294 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 429914 610954
rect 429294 610634 429914 610718
rect 429294 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 429914 610634
rect 429294 574954 429914 610398
rect 429294 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 429914 574954
rect 429294 574634 429914 574718
rect 429294 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 429914 574634
rect 429294 538954 429914 574398
rect 429294 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 429914 538954
rect 429294 538634 429914 538718
rect 429294 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 429914 538634
rect 429294 502954 429914 538398
rect 429294 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 429914 502954
rect 429294 502634 429914 502718
rect 429294 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 429914 502634
rect 429294 466954 429914 502398
rect 429294 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 429914 466954
rect 429294 466634 429914 466718
rect 429294 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 429914 466634
rect 429294 430954 429914 466398
rect 429294 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 429914 430954
rect 429294 430634 429914 430718
rect 429294 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 429914 430634
rect 429294 394954 429914 430398
rect 429294 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 429914 394954
rect 429294 394634 429914 394718
rect 429294 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 429914 394634
rect 429294 358954 429914 394398
rect 429294 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 429914 358954
rect 429294 358634 429914 358718
rect 429294 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 429914 358634
rect 429294 322954 429914 358398
rect 429294 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 429914 322954
rect 429294 322634 429914 322718
rect 429294 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 429914 322634
rect 429294 286954 429914 322398
rect 429294 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 429914 286954
rect 429294 286634 429914 286718
rect 429294 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 429914 286634
rect 429294 250954 429914 286398
rect 429294 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 429914 250954
rect 429294 250634 429914 250718
rect 429294 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 429914 250634
rect 429294 214954 429914 250398
rect 429294 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 429914 214954
rect 429294 214634 429914 214718
rect 429294 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 429914 214634
rect 429294 178954 429914 214398
rect 429294 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 429914 178954
rect 429294 178634 429914 178718
rect 429294 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 429914 178634
rect 429294 142954 429914 178398
rect 429294 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 429914 142954
rect 429294 142634 429914 142718
rect 429294 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 429914 142634
rect 429294 106954 429914 142398
rect 429294 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 429914 106954
rect 429294 106634 429914 106718
rect 429294 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 429914 106634
rect 429294 70954 429914 106398
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7066 429914 34398
rect 429294 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 429914 -7066
rect 429294 -7386 429914 -7302
rect 429294 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 429914 -7386
rect 429294 -7654 429914 -7622
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 438294 705798 438914 711590
rect 438294 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 438914 705798
rect 438294 705478 438914 705562
rect 438294 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 438914 705478
rect 438294 691954 438914 705242
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 655954 438914 691398
rect 438294 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 438914 655954
rect 438294 655634 438914 655718
rect 438294 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 438914 655634
rect 438294 619954 438914 655398
rect 438294 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 438914 619954
rect 438294 619634 438914 619718
rect 438294 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 438914 619634
rect 438294 583954 438914 619398
rect 438294 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 438914 583954
rect 438294 583634 438914 583718
rect 438294 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 438914 583634
rect 438294 547954 438914 583398
rect 438294 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 438914 547954
rect 438294 547634 438914 547718
rect 438294 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 438914 547634
rect 438294 511954 438914 547398
rect 438294 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 438914 511954
rect 438294 511634 438914 511718
rect 438294 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 438914 511634
rect 438294 475954 438914 511398
rect 438294 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 438914 475954
rect 438294 475634 438914 475718
rect 438294 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 438914 475634
rect 438294 439954 438914 475398
rect 438294 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 438914 439954
rect 438294 439634 438914 439718
rect 438294 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 438914 439634
rect 438294 403954 438914 439398
rect 438294 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 438914 403954
rect 438294 403634 438914 403718
rect 438294 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 438914 403634
rect 438294 367954 438914 403398
rect 438294 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 438914 367954
rect 438294 367634 438914 367718
rect 438294 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 438914 367634
rect 438294 331954 438914 367398
rect 438294 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 438914 331954
rect 438294 331634 438914 331718
rect 438294 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 438914 331634
rect 438294 295954 438914 331398
rect 438294 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 438914 295954
rect 438294 295634 438914 295718
rect 438294 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 438914 295634
rect 438294 259954 438914 295398
rect 438294 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 438914 259954
rect 438294 259634 438914 259718
rect 438294 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 438914 259634
rect 438294 223954 438914 259398
rect 438294 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 438914 223954
rect 438294 223634 438914 223718
rect 438294 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 438914 223634
rect 438294 187954 438914 223398
rect 438294 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 438914 187954
rect 438294 187634 438914 187718
rect 438294 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 438914 187634
rect 438294 151954 438914 187398
rect 438294 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 438914 151954
rect 438294 151634 438914 151718
rect 438294 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 438914 151634
rect 438294 115954 438914 151398
rect 438294 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 438914 115954
rect 438294 115634 438914 115718
rect 438294 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 438914 115634
rect 438294 79954 438914 115398
rect 438294 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 438914 79954
rect 438294 79634 438914 79718
rect 438294 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 438914 79634
rect 438294 43954 438914 79398
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1306 438914 7398
rect 438294 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 438914 -1306
rect 438294 -1626 438914 -1542
rect 438294 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 438914 -1626
rect 438294 -7654 438914 -1862
rect 442794 706758 443414 711590
rect 442794 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 443414 706758
rect 442794 706438 443414 706522
rect 442794 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 443414 706438
rect 442794 696454 443414 706202
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 660454 443414 695898
rect 442794 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 443414 660454
rect 442794 660134 443414 660218
rect 442794 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 443414 660134
rect 442794 624454 443414 659898
rect 442794 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 443414 624454
rect 442794 624134 443414 624218
rect 442794 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 443414 624134
rect 442794 588454 443414 623898
rect 442794 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 443414 588454
rect 442794 588134 443414 588218
rect 442794 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 443414 588134
rect 442794 552454 443414 587898
rect 442794 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 443414 552454
rect 442794 552134 443414 552218
rect 442794 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 443414 552134
rect 442794 516454 443414 551898
rect 442794 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 443414 516454
rect 442794 516134 443414 516218
rect 442794 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 443414 516134
rect 442794 480454 443414 515898
rect 442794 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 443414 480454
rect 442794 480134 443414 480218
rect 442794 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 443414 480134
rect 442794 444454 443414 479898
rect 442794 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 443414 444454
rect 442794 444134 443414 444218
rect 442794 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 443414 444134
rect 442794 408454 443414 443898
rect 442794 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 443414 408454
rect 442794 408134 443414 408218
rect 442794 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 443414 408134
rect 442794 372454 443414 407898
rect 442794 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 443414 372454
rect 442794 372134 443414 372218
rect 442794 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 443414 372134
rect 442794 336454 443414 371898
rect 442794 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 443414 336454
rect 442794 336134 443414 336218
rect 442794 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 443414 336134
rect 442794 300454 443414 335898
rect 442794 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 443414 300454
rect 442794 300134 443414 300218
rect 442794 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 443414 300134
rect 442794 264454 443414 299898
rect 442794 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 443414 264454
rect 442794 264134 443414 264218
rect 442794 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 443414 264134
rect 442794 228454 443414 263898
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 192454 443414 227898
rect 442794 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 443414 192454
rect 442794 192134 443414 192218
rect 442794 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 443414 192134
rect 442794 156454 443414 191898
rect 442794 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 443414 156454
rect 442794 156134 443414 156218
rect 442794 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 443414 156134
rect 442794 120454 443414 155898
rect 442794 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 443414 120454
rect 442794 120134 443414 120218
rect 442794 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 443414 120134
rect 442794 84454 443414 119898
rect 442794 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 443414 84454
rect 442794 84134 443414 84218
rect 442794 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 443414 84134
rect 442794 48454 443414 83898
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2266 443414 11898
rect 442794 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 443414 -2266
rect 442794 -2586 443414 -2502
rect 442794 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 443414 -2586
rect 442794 -7654 443414 -2822
rect 447294 707718 447914 711590
rect 447294 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 447914 707718
rect 447294 707398 447914 707482
rect 447294 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 447914 707398
rect 447294 700954 447914 707162
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 664954 447914 700398
rect 447294 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 447914 664954
rect 447294 664634 447914 664718
rect 447294 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 447914 664634
rect 447294 628954 447914 664398
rect 447294 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 447914 628954
rect 447294 628634 447914 628718
rect 447294 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 447914 628634
rect 447294 592954 447914 628398
rect 447294 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 447914 592954
rect 447294 592634 447914 592718
rect 447294 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 447914 592634
rect 447294 556954 447914 592398
rect 447294 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 447914 556954
rect 447294 556634 447914 556718
rect 447294 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 447914 556634
rect 447294 520954 447914 556398
rect 447294 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 447914 520954
rect 447294 520634 447914 520718
rect 447294 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 447914 520634
rect 447294 484954 447914 520398
rect 447294 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 447914 484954
rect 447294 484634 447914 484718
rect 447294 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 447914 484634
rect 447294 448954 447914 484398
rect 447294 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 447914 448954
rect 447294 448634 447914 448718
rect 447294 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 447914 448634
rect 447294 412954 447914 448398
rect 447294 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 447914 412954
rect 447294 412634 447914 412718
rect 447294 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 447914 412634
rect 447294 376954 447914 412398
rect 447294 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 447914 376954
rect 447294 376634 447914 376718
rect 447294 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 447914 376634
rect 447294 340954 447914 376398
rect 447294 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 447914 340954
rect 447294 340634 447914 340718
rect 447294 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 447914 340634
rect 447294 304954 447914 340398
rect 447294 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 447914 304954
rect 447294 304634 447914 304718
rect 447294 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 447914 304634
rect 447294 268954 447914 304398
rect 447294 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 447914 268954
rect 447294 268634 447914 268718
rect 447294 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 447914 268634
rect 447294 232954 447914 268398
rect 447294 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 447914 232954
rect 447294 232634 447914 232718
rect 447294 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 447914 232634
rect 447294 196954 447914 232398
rect 447294 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 447914 196954
rect 447294 196634 447914 196718
rect 447294 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 447914 196634
rect 447294 160954 447914 196398
rect 447294 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 447914 160954
rect 447294 160634 447914 160718
rect 447294 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 447914 160634
rect 447294 124954 447914 160398
rect 447294 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 447914 124954
rect 447294 124634 447914 124718
rect 447294 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 447914 124634
rect 447294 88954 447914 124398
rect 447294 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 447914 88954
rect 447294 88634 447914 88718
rect 447294 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 447914 88634
rect 447294 52954 447914 88398
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3226 447914 16398
rect 447294 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 447914 -3226
rect 447294 -3546 447914 -3462
rect 447294 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 447914 -3546
rect 447294 -7654 447914 -3782
rect 451794 708678 452414 711590
rect 451794 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 452414 708678
rect 451794 708358 452414 708442
rect 451794 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 452414 708358
rect 451794 669454 452414 708122
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4186 452414 20898
rect 451794 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 452414 -4186
rect 451794 -4506 452414 -4422
rect 451794 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 452414 -4506
rect 451794 -7654 452414 -4742
rect 456294 709638 456914 711590
rect 456294 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 456914 709638
rect 456294 709318 456914 709402
rect 456294 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 456914 709318
rect 456294 673954 456914 709082
rect 456294 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 456914 673954
rect 456294 673634 456914 673718
rect 456294 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 456914 673634
rect 456294 637954 456914 673398
rect 456294 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 456914 637954
rect 456294 637634 456914 637718
rect 456294 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 456914 637634
rect 456294 601954 456914 637398
rect 456294 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 456914 601954
rect 456294 601634 456914 601718
rect 456294 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 456914 601634
rect 456294 565954 456914 601398
rect 456294 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 456914 565954
rect 456294 565634 456914 565718
rect 456294 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 456914 565634
rect 456294 529954 456914 565398
rect 456294 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 456914 529954
rect 456294 529634 456914 529718
rect 456294 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 456914 529634
rect 456294 493954 456914 529398
rect 456294 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 456914 493954
rect 456294 493634 456914 493718
rect 456294 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 456914 493634
rect 456294 457954 456914 493398
rect 456294 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 456914 457954
rect 456294 457634 456914 457718
rect 456294 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 456914 457634
rect 456294 421954 456914 457398
rect 456294 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 456914 421954
rect 456294 421634 456914 421718
rect 456294 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 456914 421634
rect 456294 385954 456914 421398
rect 456294 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 456914 385954
rect 456294 385634 456914 385718
rect 456294 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 456914 385634
rect 456294 349954 456914 385398
rect 456294 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 456914 349954
rect 456294 349634 456914 349718
rect 456294 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 456914 349634
rect 456294 313954 456914 349398
rect 456294 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 456914 313954
rect 456294 313634 456914 313718
rect 456294 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 456914 313634
rect 456294 277954 456914 313398
rect 456294 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 456914 277954
rect 456294 277634 456914 277718
rect 456294 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 456914 277634
rect 456294 241954 456914 277398
rect 456294 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 456914 241954
rect 456294 241634 456914 241718
rect 456294 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 456914 241634
rect 456294 205954 456914 241398
rect 456294 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 456914 205954
rect 456294 205634 456914 205718
rect 456294 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 456914 205634
rect 456294 169954 456914 205398
rect 456294 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 456914 169954
rect 456294 169634 456914 169718
rect 456294 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 456914 169634
rect 456294 133954 456914 169398
rect 456294 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 456914 133954
rect 456294 133634 456914 133718
rect 456294 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 456914 133634
rect 456294 97954 456914 133398
rect 456294 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 456914 97954
rect 456294 97634 456914 97718
rect 456294 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 456914 97634
rect 456294 61954 456914 97398
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5146 456914 25398
rect 456294 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 456914 -5146
rect 456294 -5466 456914 -5382
rect 456294 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 456914 -5466
rect 456294 -7654 456914 -5702
rect 460794 710598 461414 711590
rect 460794 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 461414 710598
rect 460794 710278 461414 710362
rect 460794 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 461414 710278
rect 460794 678454 461414 710042
rect 460794 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 461414 678454
rect 460794 678134 461414 678218
rect 460794 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 461414 678134
rect 460794 642454 461414 677898
rect 460794 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 461414 642454
rect 460794 642134 461414 642218
rect 460794 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 461414 642134
rect 460794 606454 461414 641898
rect 460794 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 461414 606454
rect 460794 606134 461414 606218
rect 460794 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 461414 606134
rect 460794 570454 461414 605898
rect 460794 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 461414 570454
rect 460794 570134 461414 570218
rect 460794 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 461414 570134
rect 460794 534454 461414 569898
rect 460794 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 461414 534454
rect 460794 534134 461414 534218
rect 460794 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 461414 534134
rect 460794 498454 461414 533898
rect 460794 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 461414 498454
rect 460794 498134 461414 498218
rect 460794 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 461414 498134
rect 460794 462454 461414 497898
rect 460794 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 461414 462454
rect 460794 462134 461414 462218
rect 460794 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 461414 462134
rect 460794 426454 461414 461898
rect 460794 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 461414 426454
rect 460794 426134 461414 426218
rect 460794 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 461414 426134
rect 460794 390454 461414 425898
rect 460794 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 461414 390454
rect 460794 390134 461414 390218
rect 460794 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 461414 390134
rect 460794 354454 461414 389898
rect 460794 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 461414 354454
rect 460794 354134 461414 354218
rect 460794 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 461414 354134
rect 460794 318454 461414 353898
rect 460794 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 461414 318454
rect 460794 318134 461414 318218
rect 460794 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 461414 318134
rect 460794 282454 461414 317898
rect 460794 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 461414 282454
rect 460794 282134 461414 282218
rect 460794 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 461414 282134
rect 460794 246454 461414 281898
rect 460794 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 461414 246454
rect 460794 246134 461414 246218
rect 460794 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 461414 246134
rect 460794 210454 461414 245898
rect 460794 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 461414 210454
rect 460794 210134 461414 210218
rect 460794 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 461414 210134
rect 460794 174454 461414 209898
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 460794 138454 461414 173898
rect 460794 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 461414 138454
rect 460794 138134 461414 138218
rect 460794 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 461414 138134
rect 460794 102454 461414 137898
rect 460794 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 461414 102454
rect 460794 102134 461414 102218
rect 460794 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 461414 102134
rect 460794 66454 461414 101898
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6106 461414 29898
rect 460794 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 461414 -6106
rect 460794 -6426 461414 -6342
rect 460794 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 461414 -6426
rect 460794 -7654 461414 -6662
rect 465294 711558 465914 711590
rect 465294 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 465914 711558
rect 465294 711238 465914 711322
rect 465294 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 465914 711238
rect 465294 682954 465914 711002
rect 465294 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 465914 682954
rect 465294 682634 465914 682718
rect 465294 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 465914 682634
rect 465294 646954 465914 682398
rect 465294 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 465914 646954
rect 465294 646634 465914 646718
rect 465294 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 465914 646634
rect 465294 610954 465914 646398
rect 465294 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 465914 610954
rect 465294 610634 465914 610718
rect 465294 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 465914 610634
rect 465294 574954 465914 610398
rect 465294 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 465914 574954
rect 465294 574634 465914 574718
rect 465294 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 465914 574634
rect 465294 538954 465914 574398
rect 465294 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 465914 538954
rect 465294 538634 465914 538718
rect 465294 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 465914 538634
rect 465294 502954 465914 538398
rect 465294 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 465914 502954
rect 465294 502634 465914 502718
rect 465294 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 465914 502634
rect 465294 466954 465914 502398
rect 465294 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 465914 466954
rect 465294 466634 465914 466718
rect 465294 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 465914 466634
rect 465294 430954 465914 466398
rect 465294 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 465914 430954
rect 465294 430634 465914 430718
rect 465294 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 465914 430634
rect 465294 394954 465914 430398
rect 465294 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 465914 394954
rect 465294 394634 465914 394718
rect 465294 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 465914 394634
rect 465294 358954 465914 394398
rect 465294 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 465914 358954
rect 465294 358634 465914 358718
rect 465294 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 465914 358634
rect 465294 322954 465914 358398
rect 465294 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 465914 322954
rect 465294 322634 465914 322718
rect 465294 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 465914 322634
rect 465294 286954 465914 322398
rect 465294 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 465914 286954
rect 465294 286634 465914 286718
rect 465294 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 465914 286634
rect 465294 250954 465914 286398
rect 465294 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 465914 250954
rect 465294 250634 465914 250718
rect 465294 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 465914 250634
rect 465294 214954 465914 250398
rect 465294 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 465914 214954
rect 465294 214634 465914 214718
rect 465294 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 465914 214634
rect 465294 178954 465914 214398
rect 465294 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 465914 178954
rect 465294 178634 465914 178718
rect 465294 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 465914 178634
rect 465294 142954 465914 178398
rect 465294 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 465914 142954
rect 465294 142634 465914 142718
rect 465294 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 465914 142634
rect 465294 106954 465914 142398
rect 465294 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 465914 106954
rect 465294 106634 465914 106718
rect 465294 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 465914 106634
rect 465294 70954 465914 106398
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7066 465914 34398
rect 465294 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 465914 -7066
rect 465294 -7386 465914 -7302
rect 465294 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 465914 -7386
rect 465294 -7654 465914 -7622
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 474294 705798 474914 711590
rect 474294 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 474914 705798
rect 474294 705478 474914 705562
rect 474294 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 474914 705478
rect 474294 691954 474914 705242
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 655954 474914 691398
rect 474294 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 474914 655954
rect 474294 655634 474914 655718
rect 474294 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 474914 655634
rect 474294 619954 474914 655398
rect 474294 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 474914 619954
rect 474294 619634 474914 619718
rect 474294 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 474914 619634
rect 474294 583954 474914 619398
rect 474294 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 474914 583954
rect 474294 583634 474914 583718
rect 474294 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 474914 583634
rect 474294 547954 474914 583398
rect 474294 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 474914 547954
rect 474294 547634 474914 547718
rect 474294 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 474914 547634
rect 474294 511954 474914 547398
rect 474294 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 474914 511954
rect 474294 511634 474914 511718
rect 474294 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 474914 511634
rect 474294 475954 474914 511398
rect 474294 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 474914 475954
rect 474294 475634 474914 475718
rect 474294 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 474914 475634
rect 474294 439954 474914 475398
rect 474294 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 474914 439954
rect 474294 439634 474914 439718
rect 474294 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 474914 439634
rect 474294 403954 474914 439398
rect 474294 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 474914 403954
rect 474294 403634 474914 403718
rect 474294 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 474914 403634
rect 474294 367954 474914 403398
rect 474294 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 474914 367954
rect 474294 367634 474914 367718
rect 474294 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 474914 367634
rect 474294 331954 474914 367398
rect 474294 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 474914 331954
rect 474294 331634 474914 331718
rect 474294 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 474914 331634
rect 474294 295954 474914 331398
rect 474294 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 474914 295954
rect 474294 295634 474914 295718
rect 474294 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 474914 295634
rect 474294 259954 474914 295398
rect 474294 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 474914 259954
rect 474294 259634 474914 259718
rect 474294 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 474914 259634
rect 474294 223954 474914 259398
rect 474294 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 474914 223954
rect 474294 223634 474914 223718
rect 474294 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 474914 223634
rect 474294 187954 474914 223398
rect 474294 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 474914 187954
rect 474294 187634 474914 187718
rect 474294 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 474914 187634
rect 474294 151954 474914 187398
rect 474294 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 474914 151954
rect 474294 151634 474914 151718
rect 474294 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 474914 151634
rect 474294 115954 474914 151398
rect 474294 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 474914 115954
rect 474294 115634 474914 115718
rect 474294 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 474914 115634
rect 474294 79954 474914 115398
rect 474294 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 474914 79954
rect 474294 79634 474914 79718
rect 474294 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 474914 79634
rect 474294 43954 474914 79398
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1306 474914 7398
rect 474294 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 474914 -1306
rect 474294 -1626 474914 -1542
rect 474294 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 474914 -1626
rect 474294 -7654 474914 -1862
rect 478794 706758 479414 711590
rect 478794 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 479414 706758
rect 478794 706438 479414 706522
rect 478794 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 479414 706438
rect 478794 696454 479414 706202
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 660454 479414 695898
rect 478794 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 479414 660454
rect 478794 660134 479414 660218
rect 478794 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 479414 660134
rect 478794 624454 479414 659898
rect 478794 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 479414 624454
rect 478794 624134 479414 624218
rect 478794 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 479414 624134
rect 478794 588454 479414 623898
rect 478794 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 479414 588454
rect 478794 588134 479414 588218
rect 478794 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 479414 588134
rect 478794 552454 479414 587898
rect 478794 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 479414 552454
rect 478794 552134 479414 552218
rect 478794 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 479414 552134
rect 478794 516454 479414 551898
rect 478794 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 479414 516454
rect 478794 516134 479414 516218
rect 478794 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 479414 516134
rect 478794 480454 479414 515898
rect 478794 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 479414 480454
rect 478794 480134 479414 480218
rect 478794 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 479414 480134
rect 478794 444454 479414 479898
rect 478794 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 479414 444454
rect 478794 444134 479414 444218
rect 478794 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 479414 444134
rect 478794 408454 479414 443898
rect 478794 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 479414 408454
rect 478794 408134 479414 408218
rect 478794 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 479414 408134
rect 478794 372454 479414 407898
rect 478794 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 479414 372454
rect 478794 372134 479414 372218
rect 478794 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 479414 372134
rect 478794 336454 479414 371898
rect 478794 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 479414 336454
rect 478794 336134 479414 336218
rect 478794 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 479414 336134
rect 478794 300454 479414 335898
rect 478794 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 479414 300454
rect 478794 300134 479414 300218
rect 478794 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 479414 300134
rect 478794 264454 479414 299898
rect 478794 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 479414 264454
rect 478794 264134 479414 264218
rect 478794 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 479414 264134
rect 478794 228454 479414 263898
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 192454 479414 227898
rect 478794 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 479414 192454
rect 478794 192134 479414 192218
rect 478794 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 479414 192134
rect 478794 156454 479414 191898
rect 478794 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 479414 156454
rect 478794 156134 479414 156218
rect 478794 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 479414 156134
rect 478794 120454 479414 155898
rect 478794 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 479414 120454
rect 478794 120134 479414 120218
rect 478794 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 479414 120134
rect 478794 84454 479414 119898
rect 478794 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 479414 84454
rect 478794 84134 479414 84218
rect 478794 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 479414 84134
rect 478794 48454 479414 83898
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2266 479414 11898
rect 478794 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 479414 -2266
rect 478794 -2586 479414 -2502
rect 478794 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 479414 -2586
rect 478794 -7654 479414 -2822
rect 483294 707718 483914 711590
rect 483294 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 483914 707718
rect 483294 707398 483914 707482
rect 483294 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 483914 707398
rect 483294 700954 483914 707162
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 664954 483914 700398
rect 483294 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 483914 664954
rect 483294 664634 483914 664718
rect 483294 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 483914 664634
rect 483294 628954 483914 664398
rect 483294 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 483914 628954
rect 483294 628634 483914 628718
rect 483294 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 483914 628634
rect 483294 592954 483914 628398
rect 483294 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 483914 592954
rect 483294 592634 483914 592718
rect 483294 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 483914 592634
rect 483294 556954 483914 592398
rect 483294 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 483914 556954
rect 483294 556634 483914 556718
rect 483294 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 483914 556634
rect 483294 520954 483914 556398
rect 483294 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 483914 520954
rect 483294 520634 483914 520718
rect 483294 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 483914 520634
rect 483294 484954 483914 520398
rect 483294 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 483914 484954
rect 483294 484634 483914 484718
rect 483294 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 483914 484634
rect 483294 448954 483914 484398
rect 483294 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 483914 448954
rect 483294 448634 483914 448718
rect 483294 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 483914 448634
rect 483294 412954 483914 448398
rect 483294 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 483914 412954
rect 483294 412634 483914 412718
rect 483294 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 483914 412634
rect 483294 376954 483914 412398
rect 483294 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 483914 376954
rect 483294 376634 483914 376718
rect 483294 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 483914 376634
rect 483294 340954 483914 376398
rect 483294 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 483914 340954
rect 483294 340634 483914 340718
rect 483294 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 483914 340634
rect 483294 304954 483914 340398
rect 483294 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 483914 304954
rect 483294 304634 483914 304718
rect 483294 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 483914 304634
rect 483294 268954 483914 304398
rect 483294 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 483914 268954
rect 483294 268634 483914 268718
rect 483294 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 483914 268634
rect 483294 232954 483914 268398
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 124954 483914 160398
rect 483294 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 483914 124954
rect 483294 124634 483914 124718
rect 483294 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 483914 124634
rect 483294 88954 483914 124398
rect 483294 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 483914 88954
rect 483294 88634 483914 88718
rect 483294 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 483914 88634
rect 483294 52954 483914 88398
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3226 483914 16398
rect 483294 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 483914 -3226
rect 483294 -3546 483914 -3462
rect 483294 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 483914 -3546
rect 483294 -7654 483914 -3782
rect 487794 708678 488414 711590
rect 487794 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 488414 708678
rect 487794 708358 488414 708442
rect 487794 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 488414 708358
rect 487794 669454 488414 708122
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4186 488414 20898
rect 487794 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 488414 -4186
rect 487794 -4506 488414 -4422
rect 487794 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 488414 -4506
rect 487794 -7654 488414 -4742
rect 492294 709638 492914 711590
rect 492294 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 492914 709638
rect 492294 709318 492914 709402
rect 492294 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 492914 709318
rect 492294 673954 492914 709082
rect 492294 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 492914 673954
rect 492294 673634 492914 673718
rect 492294 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 492914 673634
rect 492294 637954 492914 673398
rect 492294 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 492914 637954
rect 492294 637634 492914 637718
rect 492294 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 492914 637634
rect 492294 601954 492914 637398
rect 492294 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 492914 601954
rect 492294 601634 492914 601718
rect 492294 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 492914 601634
rect 492294 565954 492914 601398
rect 492294 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 492914 565954
rect 492294 565634 492914 565718
rect 492294 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 492914 565634
rect 492294 529954 492914 565398
rect 492294 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 492914 529954
rect 492294 529634 492914 529718
rect 492294 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 492914 529634
rect 492294 493954 492914 529398
rect 492294 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 492914 493954
rect 492294 493634 492914 493718
rect 492294 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 492914 493634
rect 492294 457954 492914 493398
rect 492294 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 492914 457954
rect 492294 457634 492914 457718
rect 492294 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 492914 457634
rect 492294 421954 492914 457398
rect 492294 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 492914 421954
rect 492294 421634 492914 421718
rect 492294 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 492914 421634
rect 492294 385954 492914 421398
rect 492294 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 492914 385954
rect 492294 385634 492914 385718
rect 492294 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 492914 385634
rect 492294 349954 492914 385398
rect 492294 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 492914 349954
rect 492294 349634 492914 349718
rect 492294 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 492914 349634
rect 492294 313954 492914 349398
rect 492294 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 492914 313954
rect 492294 313634 492914 313718
rect 492294 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 492914 313634
rect 492294 277954 492914 313398
rect 492294 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 492914 277954
rect 492294 277634 492914 277718
rect 492294 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 492914 277634
rect 492294 241954 492914 277398
rect 492294 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 492914 241954
rect 492294 241634 492914 241718
rect 492294 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 492914 241634
rect 492294 205954 492914 241398
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 133954 492914 169398
rect 492294 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 492914 133954
rect 492294 133634 492914 133718
rect 492294 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 492914 133634
rect 492294 97954 492914 133398
rect 492294 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 492914 97954
rect 492294 97634 492914 97718
rect 492294 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 492914 97634
rect 492294 61954 492914 97398
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5146 492914 25398
rect 492294 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 492914 -5146
rect 492294 -5466 492914 -5382
rect 492294 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 492914 -5466
rect 492294 -7654 492914 -5702
rect 496794 710598 497414 711590
rect 496794 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 497414 710598
rect 496794 710278 497414 710362
rect 496794 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 497414 710278
rect 496794 678454 497414 710042
rect 496794 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 497414 678454
rect 496794 678134 497414 678218
rect 496794 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 497414 678134
rect 496794 642454 497414 677898
rect 496794 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 497414 642454
rect 496794 642134 497414 642218
rect 496794 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 497414 642134
rect 496794 606454 497414 641898
rect 496794 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 497414 606454
rect 496794 606134 497414 606218
rect 496794 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 497414 606134
rect 496794 570454 497414 605898
rect 496794 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 497414 570454
rect 496794 570134 497414 570218
rect 496794 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 497414 570134
rect 496794 534454 497414 569898
rect 496794 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 497414 534454
rect 496794 534134 497414 534218
rect 496794 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 497414 534134
rect 496794 498454 497414 533898
rect 496794 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 497414 498454
rect 496794 498134 497414 498218
rect 496794 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 497414 498134
rect 496794 462454 497414 497898
rect 496794 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 497414 462454
rect 496794 462134 497414 462218
rect 496794 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 497414 462134
rect 496794 426454 497414 461898
rect 496794 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 497414 426454
rect 496794 426134 497414 426218
rect 496794 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 497414 426134
rect 496794 390454 497414 425898
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 354454 497414 389898
rect 496794 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 497414 354454
rect 496794 354134 497414 354218
rect 496794 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 497414 354134
rect 496794 318454 497414 353898
rect 496794 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 497414 318454
rect 496794 318134 497414 318218
rect 496794 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 497414 318134
rect 496794 282454 497414 317898
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 246454 497414 281898
rect 496794 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 497414 246454
rect 496794 246134 497414 246218
rect 496794 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 497414 246134
rect 496794 210454 497414 245898
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 138454 497414 173898
rect 496794 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 497414 138454
rect 496794 138134 497414 138218
rect 496794 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 497414 138134
rect 496794 102454 497414 137898
rect 496794 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 497414 102454
rect 496794 102134 497414 102218
rect 496794 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 497414 102134
rect 496794 66454 497414 101898
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6106 497414 29898
rect 496794 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 497414 -6106
rect 496794 -6426 497414 -6342
rect 496794 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 497414 -6426
rect 496794 -7654 497414 -6662
rect 501294 711558 501914 711590
rect 501294 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 501914 711558
rect 501294 711238 501914 711322
rect 501294 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 501914 711238
rect 501294 682954 501914 711002
rect 501294 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 501914 682954
rect 501294 682634 501914 682718
rect 501294 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 501914 682634
rect 501294 646954 501914 682398
rect 501294 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 501914 646954
rect 501294 646634 501914 646718
rect 501294 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 501914 646634
rect 501294 610954 501914 646398
rect 501294 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 501914 610954
rect 501294 610634 501914 610718
rect 501294 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 501914 610634
rect 501294 574954 501914 610398
rect 501294 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 501914 574954
rect 501294 574634 501914 574718
rect 501294 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 501914 574634
rect 501294 538954 501914 574398
rect 501294 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 501914 538954
rect 501294 538634 501914 538718
rect 501294 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 501914 538634
rect 501294 502954 501914 538398
rect 501294 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 501914 502954
rect 501294 502634 501914 502718
rect 501294 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 501914 502634
rect 501294 466954 501914 502398
rect 501294 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 501914 466954
rect 501294 466634 501914 466718
rect 501294 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 501914 466634
rect 501294 430954 501914 466398
rect 501294 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 501914 430954
rect 501294 430634 501914 430718
rect 501294 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 501914 430634
rect 501294 394954 501914 430398
rect 501294 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 501914 394954
rect 501294 394634 501914 394718
rect 501294 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 501914 394634
rect 501294 358954 501914 394398
rect 501294 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 501914 358954
rect 501294 358634 501914 358718
rect 501294 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 501914 358634
rect 501294 322954 501914 358398
rect 501294 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 501914 322954
rect 501294 322634 501914 322718
rect 501294 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 501914 322634
rect 501294 286954 501914 322398
rect 501294 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 501914 286954
rect 501294 286634 501914 286718
rect 501294 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 501914 286634
rect 501294 250954 501914 286398
rect 501294 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 501914 250954
rect 501294 250634 501914 250718
rect 501294 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 501914 250634
rect 501294 214954 501914 250398
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 142954 501914 178398
rect 501294 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 501914 142954
rect 501294 142634 501914 142718
rect 501294 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 501914 142634
rect 501294 106954 501914 142398
rect 501294 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 501914 106954
rect 501294 106634 501914 106718
rect 501294 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 501914 106634
rect 501294 70954 501914 106398
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7066 501914 34398
rect 501294 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 501914 -7066
rect 501294 -7386 501914 -7302
rect 501294 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 501914 -7386
rect 501294 -7654 501914 -7622
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 510294 705798 510914 711590
rect 510294 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 510914 705798
rect 510294 705478 510914 705562
rect 510294 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 510914 705478
rect 510294 691954 510914 705242
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 655954 510914 691398
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 619954 510914 655398
rect 510294 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 510914 619954
rect 510294 619634 510914 619718
rect 510294 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 510914 619634
rect 510294 583954 510914 619398
rect 510294 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 510914 583954
rect 510294 583634 510914 583718
rect 510294 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 510914 583634
rect 510294 547954 510914 583398
rect 510294 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 510914 547954
rect 510294 547634 510914 547718
rect 510294 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 510914 547634
rect 510294 511954 510914 547398
rect 510294 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 510914 511954
rect 510294 511634 510914 511718
rect 510294 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 510914 511634
rect 510294 475954 510914 511398
rect 510294 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 510914 475954
rect 510294 475634 510914 475718
rect 510294 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 510914 475634
rect 510294 439954 510914 475398
rect 510294 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 510914 439954
rect 510294 439634 510914 439718
rect 510294 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 510914 439634
rect 510294 403954 510914 439398
rect 510294 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 510914 403954
rect 510294 403634 510914 403718
rect 510294 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 510914 403634
rect 510294 367954 510914 403398
rect 510294 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 510914 367954
rect 510294 367634 510914 367718
rect 510294 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 510914 367634
rect 510294 331954 510914 367398
rect 510294 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 510914 331954
rect 510294 331634 510914 331718
rect 510294 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 510914 331634
rect 510294 295954 510914 331398
rect 510294 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 510914 295954
rect 510294 295634 510914 295718
rect 510294 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 510914 295634
rect 510294 259954 510914 295398
rect 510294 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 510914 259954
rect 510294 259634 510914 259718
rect 510294 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 510914 259634
rect 510294 223954 510914 259398
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 151954 510914 187398
rect 510294 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 510914 151954
rect 510294 151634 510914 151718
rect 510294 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 510914 151634
rect 510294 115954 510914 151398
rect 510294 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 510914 115954
rect 510294 115634 510914 115718
rect 510294 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 510914 115634
rect 510294 79954 510914 115398
rect 510294 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 510914 79954
rect 510294 79634 510914 79718
rect 510294 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 510914 79634
rect 510294 43954 510914 79398
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1306 510914 7398
rect 510294 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 510914 -1306
rect 510294 -1626 510914 -1542
rect 510294 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 510914 -1626
rect 510294 -7654 510914 -1862
rect 514794 706758 515414 711590
rect 514794 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 515414 706758
rect 514794 706438 515414 706522
rect 514794 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 515414 706438
rect 514794 696454 515414 706202
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 624454 515414 659898
rect 514794 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 515414 624454
rect 514794 624134 515414 624218
rect 514794 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 515414 624134
rect 514794 588454 515414 623898
rect 514794 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 515414 588454
rect 514794 588134 515414 588218
rect 514794 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 515414 588134
rect 514794 552454 515414 587898
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 514794 516454 515414 551898
rect 514794 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 515414 516454
rect 514794 516134 515414 516218
rect 514794 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 515414 516134
rect 514794 480454 515414 515898
rect 514794 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 515414 480454
rect 514794 480134 515414 480218
rect 514794 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 515414 480134
rect 514794 444454 515414 479898
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 514794 408454 515414 443898
rect 514794 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 515414 408454
rect 514794 408134 515414 408218
rect 514794 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 515414 408134
rect 514794 372454 515414 407898
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 514794 264454 515414 299898
rect 514794 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 515414 264454
rect 514794 264134 515414 264218
rect 514794 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 515414 264134
rect 514794 228454 515414 263898
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 120454 515414 155898
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 514794 84454 515414 119898
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2266 515414 11898
rect 514794 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 515414 -2266
rect 514794 -2586 515414 -2502
rect 514794 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 515414 -2586
rect 514794 -7654 515414 -2822
rect 519294 707718 519914 711590
rect 519294 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 519914 707718
rect 519294 707398 519914 707482
rect 519294 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 519914 707398
rect 519294 700954 519914 707162
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 628954 519914 664398
rect 519294 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 519914 628954
rect 519294 628634 519914 628718
rect 519294 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 519914 628634
rect 519294 592954 519914 628398
rect 519294 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 519914 592954
rect 519294 592634 519914 592718
rect 519294 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 519914 592634
rect 519294 556954 519914 592398
rect 519294 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 519914 556954
rect 519294 556634 519914 556718
rect 519294 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 519914 556634
rect 519294 520954 519914 556398
rect 519294 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 519914 520954
rect 519294 520634 519914 520718
rect 519294 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 519914 520634
rect 519294 484954 519914 520398
rect 519294 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 519914 484954
rect 519294 484634 519914 484718
rect 519294 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 519914 484634
rect 519294 448954 519914 484398
rect 519294 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 519914 448954
rect 519294 448634 519914 448718
rect 519294 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 519914 448634
rect 519294 412954 519914 448398
rect 519294 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 519914 412954
rect 519294 412634 519914 412718
rect 519294 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 519914 412634
rect 519294 376954 519914 412398
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 268954 519914 304398
rect 519294 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 519914 268954
rect 519294 268634 519914 268718
rect 519294 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 519914 268634
rect 519294 232954 519914 268398
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 124954 519914 160398
rect 519294 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 519914 124954
rect 519294 124634 519914 124718
rect 519294 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 519914 124634
rect 519294 88954 519914 124398
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3226 519914 16398
rect 519294 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 519914 -3226
rect 519294 -3546 519914 -3462
rect 519294 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 519914 -3546
rect 519294 -7654 519914 -3782
rect 523794 708678 524414 711590
rect 523794 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 524414 708678
rect 523794 708358 524414 708442
rect 523794 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 524414 708358
rect 523794 669454 524414 708122
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4186 524414 20898
rect 523794 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 524414 -4186
rect 523794 -4506 524414 -4422
rect 523794 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 524414 -4506
rect 523794 -7654 524414 -4742
rect 528294 709638 528914 711590
rect 528294 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 528914 709638
rect 528294 709318 528914 709402
rect 528294 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 528914 709318
rect 528294 673954 528914 709082
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 528294 565954 528914 601398
rect 528294 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 528914 565954
rect 528294 565634 528914 565718
rect 528294 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 528914 565634
rect 528294 529954 528914 565398
rect 528294 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 528914 529954
rect 528294 529634 528914 529718
rect 528294 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 528914 529634
rect 528294 493954 528914 529398
rect 528294 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 528914 493954
rect 528294 493634 528914 493718
rect 528294 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 528914 493634
rect 528294 457954 528914 493398
rect 528294 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 528914 457954
rect 528294 457634 528914 457718
rect 528294 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 528914 457634
rect 528294 421954 528914 457398
rect 528294 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 528914 421954
rect 528294 421634 528914 421718
rect 528294 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 528914 421634
rect 528294 385954 528914 421398
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 277954 528914 313398
rect 528294 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 528914 277954
rect 528294 277634 528914 277718
rect 528294 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 528914 277634
rect 528294 241954 528914 277398
rect 528294 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 528914 241954
rect 528294 241634 528914 241718
rect 528294 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 528914 241634
rect 528294 205954 528914 241398
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 133954 528914 169398
rect 528294 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 528914 133954
rect 528294 133634 528914 133718
rect 528294 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 528914 133634
rect 528294 97954 528914 133398
rect 528294 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 528914 97954
rect 528294 97634 528914 97718
rect 528294 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 528914 97634
rect 528294 61954 528914 97398
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5146 528914 25398
rect 528294 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 528914 -5146
rect 528294 -5466 528914 -5382
rect 528294 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 528914 -5466
rect 528294 -7654 528914 -5702
rect 532794 710598 533414 711590
rect 532794 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 533414 710598
rect 532794 710278 533414 710362
rect 532794 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 533414 710278
rect 532794 678454 533414 710042
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 570454 533414 605898
rect 532794 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 533414 570454
rect 532794 570134 533414 570218
rect 532794 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 533414 570134
rect 532794 534454 533414 569898
rect 532794 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 533414 534454
rect 532794 534134 533414 534218
rect 532794 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 533414 534134
rect 532794 498454 533414 533898
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 462454 533414 497898
rect 532794 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 533414 462454
rect 532794 462134 533414 462218
rect 532794 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 533414 462134
rect 532794 426454 533414 461898
rect 532794 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 533414 426454
rect 532794 426134 533414 426218
rect 532794 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 533414 426134
rect 532794 390454 533414 425898
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 246454 533414 281898
rect 532794 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 533414 246454
rect 532794 246134 533414 246218
rect 532794 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 533414 246134
rect 532794 210454 533414 245898
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 138454 533414 173898
rect 532794 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 533414 138454
rect 532794 138134 533414 138218
rect 532794 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 533414 138134
rect 532794 102454 533414 137898
rect 532794 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 533414 102454
rect 532794 102134 533414 102218
rect 532794 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 533414 102134
rect 532794 66454 533414 101898
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6106 533414 29898
rect 532794 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 533414 -6106
rect 532794 -6426 533414 -6342
rect 532794 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 533414 -6426
rect 532794 -7654 533414 -6662
rect 537294 711558 537914 711590
rect 537294 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 537914 711558
rect 537294 711238 537914 711322
rect 537294 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 537914 711238
rect 537294 682954 537914 711002
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 537294 574954 537914 610398
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 250954 537914 286398
rect 537294 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 537914 250954
rect 537294 250634 537914 250718
rect 537294 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 537914 250634
rect 537294 214954 537914 250398
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 142954 537914 178398
rect 537294 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 537914 142954
rect 537294 142634 537914 142718
rect 537294 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 537914 142634
rect 537294 106954 537914 142398
rect 537294 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 537914 106954
rect 537294 106634 537914 106718
rect 537294 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 537914 106634
rect 537294 70954 537914 106398
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7066 537914 34398
rect 537294 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 537914 -7066
rect 537294 -7386 537914 -7302
rect 537294 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 537914 -7386
rect 537294 -7654 537914 -7622
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 546294 705798 546914 711590
rect 546294 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 546914 705798
rect 546294 705478 546914 705562
rect 546294 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 546914 705478
rect 546294 691954 546914 705242
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 295954 546914 331398
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 259954 546914 295398
rect 546294 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 546914 259954
rect 546294 259634 546914 259718
rect 546294 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 546914 259634
rect 546294 223954 546914 259398
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1306 546914 7398
rect 546294 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 546914 -1306
rect 546294 -1626 546914 -1542
rect 546294 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 546914 -1626
rect 546294 -7654 546914 -1862
rect 550794 706758 551414 711590
rect 550794 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 551414 706758
rect 550794 706438 551414 706522
rect 550794 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 551414 706438
rect 550794 696454 551414 706202
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 300454 551414 335898
rect 550794 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 551414 300454
rect 550794 300134 551414 300218
rect 550794 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 551414 300134
rect 550794 264454 551414 299898
rect 550794 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 551414 264454
rect 550794 264134 551414 264218
rect 550794 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 551414 264134
rect 550794 228454 551414 263898
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2266 551414 11898
rect 550794 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 551414 -2266
rect 550794 -2586 551414 -2502
rect 550794 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 551414 -2586
rect 550794 -7654 551414 -2822
rect 555294 707718 555914 711590
rect 555294 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 555914 707718
rect 555294 707398 555914 707482
rect 555294 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 555914 707398
rect 555294 700954 555914 707162
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3226 555914 16398
rect 555294 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 555914 -3226
rect 555294 -3546 555914 -3462
rect 555294 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 555914 -3546
rect 555294 -7654 555914 -3782
rect 559794 708678 560414 711590
rect 559794 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 560414 708678
rect 559794 708358 560414 708442
rect 559794 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 560414 708358
rect 559794 669454 560414 708122
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4186 560414 20898
rect 559794 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 560414 -4186
rect 559794 -4506 560414 -4422
rect 559794 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 560414 -4506
rect 559794 -7654 560414 -4742
rect 564294 709638 564914 711590
rect 564294 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 564914 709638
rect 564294 709318 564914 709402
rect 564294 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 564914 709318
rect 564294 673954 564914 709082
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5146 564914 25398
rect 564294 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 564914 -5146
rect 564294 -5466 564914 -5382
rect 564294 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 564914 -5466
rect 564294 -7654 564914 -5702
rect 568794 710598 569414 711590
rect 568794 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 569414 710598
rect 568794 710278 569414 710362
rect 568794 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 569414 710278
rect 568794 678454 569414 710042
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6106 569414 29898
rect 568794 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 569414 -6106
rect 568794 -6426 569414 -6342
rect 568794 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 569414 -6426
rect 568794 -7654 569414 -6662
rect 573294 711558 573914 711590
rect 573294 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 573914 711558
rect 573294 711238 573914 711322
rect 573294 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 573914 711238
rect 573294 682954 573914 711002
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7066 573914 34398
rect 573294 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 573914 -7066
rect 573294 -7386 573914 -7302
rect 573294 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 573914 -7386
rect 573294 -7654 573914 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect 582294 691954 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1306 582914 7398
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691954 586890 705242
rect 586270 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 586890 691954
rect 586270 691634 586890 691718
rect 586270 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 586890 691634
rect 586270 655954 586890 691398
rect 586270 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 586890 655954
rect 586270 655634 586890 655718
rect 586270 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 586890 655634
rect 586270 619954 586890 655398
rect 586270 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 586890 619954
rect 586270 619634 586890 619718
rect 586270 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 586890 619634
rect 586270 583954 586890 619398
rect 586270 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 586890 583954
rect 586270 583634 586890 583718
rect 586270 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 586890 583634
rect 586270 547954 586890 583398
rect 586270 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 586890 547954
rect 586270 547634 586890 547718
rect 586270 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 586890 547634
rect 586270 511954 586890 547398
rect 586270 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 586890 511954
rect 586270 511634 586890 511718
rect 586270 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 586890 511634
rect 586270 475954 586890 511398
rect 586270 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 586890 475954
rect 586270 475634 586890 475718
rect 586270 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 586890 475634
rect 586270 439954 586890 475398
rect 586270 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 586890 439954
rect 586270 439634 586890 439718
rect 586270 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 586890 439634
rect 586270 403954 586890 439398
rect 586270 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 586890 403954
rect 586270 403634 586890 403718
rect 586270 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 586890 403634
rect 586270 367954 586890 403398
rect 586270 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 586890 367954
rect 586270 367634 586890 367718
rect 586270 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 586890 367634
rect 586270 331954 586890 367398
rect 586270 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 586890 331954
rect 586270 331634 586890 331718
rect 586270 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 586890 331634
rect 586270 295954 586890 331398
rect 586270 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 586890 295954
rect 586270 295634 586890 295718
rect 586270 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 586890 295634
rect 586270 259954 586890 295398
rect 586270 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 586890 259954
rect 586270 259634 586890 259718
rect 586270 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 586890 259634
rect 586270 223954 586890 259398
rect 586270 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 586890 223954
rect 586270 223634 586890 223718
rect 586270 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 586890 223634
rect 586270 187954 586890 223398
rect 586270 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 586890 187954
rect 586270 187634 586890 187718
rect 586270 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 586890 187634
rect 586270 151954 586890 187398
rect 586270 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 586890 151954
rect 586270 151634 586890 151718
rect 586270 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 586890 151634
rect 586270 115954 586890 151398
rect 586270 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 586890 115954
rect 586270 115634 586890 115718
rect 586270 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 586890 115634
rect 586270 79954 586890 115398
rect 586270 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 586890 79954
rect 586270 79634 586890 79718
rect 586270 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 586890 79634
rect 586270 43954 586890 79398
rect 586270 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 586890 43954
rect 586270 43634 586890 43718
rect 586270 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 586890 43634
rect 586270 7954 586890 43398
rect 586270 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 586890 7954
rect 586270 7634 586890 7718
rect 586270 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 586890 7634
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 7398
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 696454 587850 706202
rect 587230 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 587850 696454
rect 587230 696134 587850 696218
rect 587230 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 587850 696134
rect 587230 660454 587850 695898
rect 587230 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 587850 660454
rect 587230 660134 587850 660218
rect 587230 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 587850 660134
rect 587230 624454 587850 659898
rect 587230 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 587850 624454
rect 587230 624134 587850 624218
rect 587230 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 587850 624134
rect 587230 588454 587850 623898
rect 587230 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 587850 588454
rect 587230 588134 587850 588218
rect 587230 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 587850 588134
rect 587230 552454 587850 587898
rect 587230 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 587850 552454
rect 587230 552134 587850 552218
rect 587230 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 587850 552134
rect 587230 516454 587850 551898
rect 587230 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 587850 516454
rect 587230 516134 587850 516218
rect 587230 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 587850 516134
rect 587230 480454 587850 515898
rect 587230 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 587850 480454
rect 587230 480134 587850 480218
rect 587230 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 587850 480134
rect 587230 444454 587850 479898
rect 587230 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 587850 444454
rect 587230 444134 587850 444218
rect 587230 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 587850 444134
rect 587230 408454 587850 443898
rect 587230 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 587850 408454
rect 587230 408134 587850 408218
rect 587230 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 587850 408134
rect 587230 372454 587850 407898
rect 587230 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 587850 372454
rect 587230 372134 587850 372218
rect 587230 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 587850 372134
rect 587230 336454 587850 371898
rect 587230 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 587850 336454
rect 587230 336134 587850 336218
rect 587230 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 587850 336134
rect 587230 300454 587850 335898
rect 587230 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 587850 300454
rect 587230 300134 587850 300218
rect 587230 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 587850 300134
rect 587230 264454 587850 299898
rect 587230 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 587850 264454
rect 587230 264134 587850 264218
rect 587230 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 587850 264134
rect 587230 228454 587850 263898
rect 587230 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 587850 228454
rect 587230 228134 587850 228218
rect 587230 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 587850 228134
rect 587230 192454 587850 227898
rect 587230 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 587850 192454
rect 587230 192134 587850 192218
rect 587230 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 587850 192134
rect 587230 156454 587850 191898
rect 587230 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 587850 156454
rect 587230 156134 587850 156218
rect 587230 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 587850 156134
rect 587230 120454 587850 155898
rect 587230 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 587850 120454
rect 587230 120134 587850 120218
rect 587230 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 587850 120134
rect 587230 84454 587850 119898
rect 587230 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 587850 84454
rect 587230 84134 587850 84218
rect 587230 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 587850 84134
rect 587230 48454 587850 83898
rect 587230 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 587850 48454
rect 587230 48134 587850 48218
rect 587230 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 587850 48134
rect 587230 12454 587850 47898
rect 587230 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 587850 12454
rect 587230 12134 587850 12218
rect 587230 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 587850 12134
rect 587230 -2266 587850 11898
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 700954 588810 707162
rect 588190 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 588810 700954
rect 588190 700634 588810 700718
rect 588190 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 588810 700634
rect 588190 664954 588810 700398
rect 588190 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 588810 664954
rect 588190 664634 588810 664718
rect 588190 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 588810 664634
rect 588190 628954 588810 664398
rect 588190 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 588810 628954
rect 588190 628634 588810 628718
rect 588190 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 588810 628634
rect 588190 592954 588810 628398
rect 588190 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 588810 592954
rect 588190 592634 588810 592718
rect 588190 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 588810 592634
rect 588190 556954 588810 592398
rect 588190 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect 588190 556634 588810 556718
rect 588190 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 588810 556634
rect 588190 520954 588810 556398
rect 588190 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 588810 520954
rect 588190 520634 588810 520718
rect 588190 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 588810 520634
rect 588190 484954 588810 520398
rect 588190 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 588810 484954
rect 588190 484634 588810 484718
rect 588190 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 588810 484634
rect 588190 448954 588810 484398
rect 588190 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 588810 448954
rect 588190 448634 588810 448718
rect 588190 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 588810 448634
rect 588190 412954 588810 448398
rect 588190 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 588810 412954
rect 588190 412634 588810 412718
rect 588190 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 588810 412634
rect 588190 376954 588810 412398
rect 588190 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect 588190 376634 588810 376718
rect 588190 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 588810 376634
rect 588190 340954 588810 376398
rect 588190 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 588810 340954
rect 588190 340634 588810 340718
rect 588190 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 588810 340634
rect 588190 304954 588810 340398
rect 588190 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 588810 304954
rect 588190 304634 588810 304718
rect 588190 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 588810 304634
rect 588190 268954 588810 304398
rect 588190 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 588810 268954
rect 588190 268634 588810 268718
rect 588190 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 588810 268634
rect 588190 232954 588810 268398
rect 588190 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 588810 232954
rect 588190 232634 588810 232718
rect 588190 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 588810 232634
rect 588190 196954 588810 232398
rect 588190 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect 588190 196634 588810 196718
rect 588190 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 588810 196634
rect 588190 160954 588810 196398
rect 588190 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 588810 160954
rect 588190 160634 588810 160718
rect 588190 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 588810 160634
rect 588190 124954 588810 160398
rect 588190 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 588810 124954
rect 588190 124634 588810 124718
rect 588190 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 588810 124634
rect 588190 88954 588810 124398
rect 588190 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 588810 88954
rect 588190 88634 588810 88718
rect 588190 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 588810 88634
rect 588190 52954 588810 88398
rect 588190 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 588810 52954
rect 588190 52634 588810 52718
rect 588190 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 588810 52634
rect 588190 16954 588810 52398
rect 588190 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect 588190 16634 588810 16718
rect 588190 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 588810 16634
rect 588190 -3226 588810 16398
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 669454 589770 708122
rect 589150 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 589770 669454
rect 589150 669134 589770 669218
rect 589150 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 589770 669134
rect 589150 633454 589770 668898
rect 589150 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 589770 633454
rect 589150 633134 589770 633218
rect 589150 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 589770 633134
rect 589150 597454 589770 632898
rect 589150 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 589770 597454
rect 589150 597134 589770 597218
rect 589150 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 589770 597134
rect 589150 561454 589770 596898
rect 589150 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 589770 561454
rect 589150 561134 589770 561218
rect 589150 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 589770 561134
rect 589150 525454 589770 560898
rect 589150 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 589770 525454
rect 589150 525134 589770 525218
rect 589150 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 589770 525134
rect 589150 489454 589770 524898
rect 589150 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 589770 489454
rect 589150 489134 589770 489218
rect 589150 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 589770 489134
rect 589150 453454 589770 488898
rect 589150 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 589770 453454
rect 589150 453134 589770 453218
rect 589150 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 589770 453134
rect 589150 417454 589770 452898
rect 589150 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 589770 417454
rect 589150 417134 589770 417218
rect 589150 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 589770 417134
rect 589150 381454 589770 416898
rect 589150 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 589770 381454
rect 589150 381134 589770 381218
rect 589150 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 589770 381134
rect 589150 345454 589770 380898
rect 589150 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 589770 345454
rect 589150 345134 589770 345218
rect 589150 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 589770 345134
rect 589150 309454 589770 344898
rect 589150 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 589770 309454
rect 589150 309134 589770 309218
rect 589150 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 589770 309134
rect 589150 273454 589770 308898
rect 589150 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 589770 273454
rect 589150 273134 589770 273218
rect 589150 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 589770 273134
rect 589150 237454 589770 272898
rect 589150 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 589770 237454
rect 589150 237134 589770 237218
rect 589150 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 589770 237134
rect 589150 201454 589770 236898
rect 589150 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 589770 201454
rect 589150 201134 589770 201218
rect 589150 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 589770 201134
rect 589150 165454 589770 200898
rect 589150 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 589770 165454
rect 589150 165134 589770 165218
rect 589150 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 589770 165134
rect 589150 129454 589770 164898
rect 589150 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 589770 129454
rect 589150 129134 589770 129218
rect 589150 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 589770 129134
rect 589150 93454 589770 128898
rect 589150 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 589770 93454
rect 589150 93134 589770 93218
rect 589150 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 589770 93134
rect 589150 57454 589770 92898
rect 589150 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 589770 57454
rect 589150 57134 589770 57218
rect 589150 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 589770 57134
rect 589150 21454 589770 56898
rect 589150 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 589770 21454
rect 589150 21134 589770 21218
rect 589150 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 589770 21134
rect 589150 -4186 589770 20898
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 673954 590730 709082
rect 590110 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 590730 673954
rect 590110 673634 590730 673718
rect 590110 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 590730 673634
rect 590110 637954 590730 673398
rect 590110 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 590730 637954
rect 590110 637634 590730 637718
rect 590110 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 590730 637634
rect 590110 601954 590730 637398
rect 590110 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 590730 601954
rect 590110 601634 590730 601718
rect 590110 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 590730 601634
rect 590110 565954 590730 601398
rect 590110 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 590730 565954
rect 590110 565634 590730 565718
rect 590110 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 590730 565634
rect 590110 529954 590730 565398
rect 590110 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 590730 529954
rect 590110 529634 590730 529718
rect 590110 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 590730 529634
rect 590110 493954 590730 529398
rect 590110 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 590730 493954
rect 590110 493634 590730 493718
rect 590110 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 590730 493634
rect 590110 457954 590730 493398
rect 590110 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 590730 457954
rect 590110 457634 590730 457718
rect 590110 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 590730 457634
rect 590110 421954 590730 457398
rect 590110 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 590730 421954
rect 590110 421634 590730 421718
rect 590110 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 590730 421634
rect 590110 385954 590730 421398
rect 590110 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 590730 385954
rect 590110 385634 590730 385718
rect 590110 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 590730 385634
rect 590110 349954 590730 385398
rect 590110 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 590730 349954
rect 590110 349634 590730 349718
rect 590110 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 590730 349634
rect 590110 313954 590730 349398
rect 590110 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 590730 313954
rect 590110 313634 590730 313718
rect 590110 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 590730 313634
rect 590110 277954 590730 313398
rect 590110 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 590730 277954
rect 590110 277634 590730 277718
rect 590110 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 590730 277634
rect 590110 241954 590730 277398
rect 590110 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 590730 241954
rect 590110 241634 590730 241718
rect 590110 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 590730 241634
rect 590110 205954 590730 241398
rect 590110 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 590730 205954
rect 590110 205634 590730 205718
rect 590110 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 590730 205634
rect 590110 169954 590730 205398
rect 590110 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 590730 169954
rect 590110 169634 590730 169718
rect 590110 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 590730 169634
rect 590110 133954 590730 169398
rect 590110 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 590730 133954
rect 590110 133634 590730 133718
rect 590110 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 590730 133634
rect 590110 97954 590730 133398
rect 590110 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 590730 97954
rect 590110 97634 590730 97718
rect 590110 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 590730 97634
rect 590110 61954 590730 97398
rect 590110 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 590730 61954
rect 590110 61634 590730 61718
rect 590110 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 590730 61634
rect 590110 25954 590730 61398
rect 590110 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 590730 25954
rect 590110 25634 590730 25718
rect 590110 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 590730 25634
rect 590110 -5146 590730 25398
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 678454 591690 710042
rect 591070 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 591690 678454
rect 591070 678134 591690 678218
rect 591070 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 591690 678134
rect 591070 642454 591690 677898
rect 591070 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 591690 642454
rect 591070 642134 591690 642218
rect 591070 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 591690 642134
rect 591070 606454 591690 641898
rect 591070 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 591690 606454
rect 591070 606134 591690 606218
rect 591070 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 591690 606134
rect 591070 570454 591690 605898
rect 591070 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 591690 570454
rect 591070 570134 591690 570218
rect 591070 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 591690 570134
rect 591070 534454 591690 569898
rect 591070 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 591690 534454
rect 591070 534134 591690 534218
rect 591070 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 591690 534134
rect 591070 498454 591690 533898
rect 591070 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 591690 498454
rect 591070 498134 591690 498218
rect 591070 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 591690 498134
rect 591070 462454 591690 497898
rect 591070 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 591690 462454
rect 591070 462134 591690 462218
rect 591070 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 591690 462134
rect 591070 426454 591690 461898
rect 591070 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 591690 426454
rect 591070 426134 591690 426218
rect 591070 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 591690 426134
rect 591070 390454 591690 425898
rect 591070 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 591690 390454
rect 591070 390134 591690 390218
rect 591070 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 591690 390134
rect 591070 354454 591690 389898
rect 591070 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 591690 354454
rect 591070 354134 591690 354218
rect 591070 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 591690 354134
rect 591070 318454 591690 353898
rect 591070 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 591690 318454
rect 591070 318134 591690 318218
rect 591070 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 591690 318134
rect 591070 282454 591690 317898
rect 591070 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 591690 282454
rect 591070 282134 591690 282218
rect 591070 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 591690 282134
rect 591070 246454 591690 281898
rect 591070 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 591690 246454
rect 591070 246134 591690 246218
rect 591070 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 591690 246134
rect 591070 210454 591690 245898
rect 591070 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 591690 210454
rect 591070 210134 591690 210218
rect 591070 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 591690 210134
rect 591070 174454 591690 209898
rect 591070 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 591690 174454
rect 591070 174134 591690 174218
rect 591070 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 591690 174134
rect 591070 138454 591690 173898
rect 591070 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 591690 138454
rect 591070 138134 591690 138218
rect 591070 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 591690 138134
rect 591070 102454 591690 137898
rect 591070 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 591690 102454
rect 591070 102134 591690 102218
rect 591070 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 591690 102134
rect 591070 66454 591690 101898
rect 591070 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 591690 66454
rect 591070 66134 591690 66218
rect 591070 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 591690 66134
rect 591070 30454 591690 65898
rect 591070 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 591690 30454
rect 591070 30134 591690 30218
rect 591070 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 591690 30134
rect 591070 -6106 591690 29898
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 682954 592650 711002
rect 592030 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect 592030 682634 592650 682718
rect 592030 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect 592030 646954 592650 682398
rect 592030 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect 592030 646634 592650 646718
rect 592030 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect 592030 610954 592650 646398
rect 592030 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect 592030 610634 592650 610718
rect 592030 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect 592030 574954 592650 610398
rect 592030 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect 592030 574634 592650 574718
rect 592030 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect 592030 538954 592650 574398
rect 592030 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect 592030 538634 592650 538718
rect 592030 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect 592030 502954 592650 538398
rect 592030 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect 592030 502634 592650 502718
rect 592030 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect 592030 466954 592650 502398
rect 592030 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect 592030 466634 592650 466718
rect 592030 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect 592030 430954 592650 466398
rect 592030 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect 592030 430634 592650 430718
rect 592030 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect 592030 394954 592650 430398
rect 592030 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect 592030 394634 592650 394718
rect 592030 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect 592030 358954 592650 394398
rect 592030 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect 592030 358634 592650 358718
rect 592030 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect 592030 322954 592650 358398
rect 592030 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect 592030 322634 592650 322718
rect 592030 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect 592030 286954 592650 322398
rect 592030 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect 592030 286634 592650 286718
rect 592030 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect 592030 250954 592650 286398
rect 592030 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect 592030 250634 592650 250718
rect 592030 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect 592030 214954 592650 250398
rect 592030 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect 592030 214634 592650 214718
rect 592030 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect 592030 178954 592650 214398
rect 592030 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect 592030 178634 592650 178718
rect 592030 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect 592030 142954 592650 178398
rect 592030 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect 592030 142634 592650 142718
rect 592030 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect 592030 106954 592650 142398
rect 592030 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect 592030 106634 592650 106718
rect 592030 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect 592030 70954 592650 106398
rect 592030 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect 592030 70634 592650 70718
rect 592030 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect 592030 34954 592650 70398
rect 592030 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect 592030 34634 592650 34718
rect 592030 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect 592030 -7066 592650 34398
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 682718 -8458 682954
rect -8374 682718 -8138 682954
rect -8694 682398 -8458 682634
rect -8374 682398 -8138 682634
rect -8694 646718 -8458 646954
rect -8374 646718 -8138 646954
rect -8694 646398 -8458 646634
rect -8374 646398 -8138 646634
rect -8694 610718 -8458 610954
rect -8374 610718 -8138 610954
rect -8694 610398 -8458 610634
rect -8374 610398 -8138 610634
rect -8694 574718 -8458 574954
rect -8374 574718 -8138 574954
rect -8694 574398 -8458 574634
rect -8374 574398 -8138 574634
rect -8694 538718 -8458 538954
rect -8374 538718 -8138 538954
rect -8694 538398 -8458 538634
rect -8374 538398 -8138 538634
rect -8694 502718 -8458 502954
rect -8374 502718 -8138 502954
rect -8694 502398 -8458 502634
rect -8374 502398 -8138 502634
rect -8694 466718 -8458 466954
rect -8374 466718 -8138 466954
rect -8694 466398 -8458 466634
rect -8374 466398 -8138 466634
rect -8694 430718 -8458 430954
rect -8374 430718 -8138 430954
rect -8694 430398 -8458 430634
rect -8374 430398 -8138 430634
rect -8694 394718 -8458 394954
rect -8374 394718 -8138 394954
rect -8694 394398 -8458 394634
rect -8374 394398 -8138 394634
rect -8694 358718 -8458 358954
rect -8374 358718 -8138 358954
rect -8694 358398 -8458 358634
rect -8374 358398 -8138 358634
rect -8694 322718 -8458 322954
rect -8374 322718 -8138 322954
rect -8694 322398 -8458 322634
rect -8374 322398 -8138 322634
rect -8694 286718 -8458 286954
rect -8374 286718 -8138 286954
rect -8694 286398 -8458 286634
rect -8374 286398 -8138 286634
rect -8694 250718 -8458 250954
rect -8374 250718 -8138 250954
rect -8694 250398 -8458 250634
rect -8374 250398 -8138 250634
rect -8694 214718 -8458 214954
rect -8374 214718 -8138 214954
rect -8694 214398 -8458 214634
rect -8374 214398 -8138 214634
rect -8694 178718 -8458 178954
rect -8374 178718 -8138 178954
rect -8694 178398 -8458 178634
rect -8374 178398 -8138 178634
rect -8694 142718 -8458 142954
rect -8374 142718 -8138 142954
rect -8694 142398 -8458 142634
rect -8374 142398 -8138 142634
rect -8694 106718 -8458 106954
rect -8374 106718 -8138 106954
rect -8694 106398 -8458 106634
rect -8374 106398 -8138 106634
rect -8694 70718 -8458 70954
rect -8374 70718 -8138 70954
rect -8694 70398 -8458 70634
rect -8374 70398 -8138 70634
rect -8694 34718 -8458 34954
rect -8374 34718 -8138 34954
rect -8694 34398 -8458 34634
rect -8374 34398 -8138 34634
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 678218 -7498 678454
rect -7414 678218 -7178 678454
rect -7734 677898 -7498 678134
rect -7414 677898 -7178 678134
rect -7734 642218 -7498 642454
rect -7414 642218 -7178 642454
rect -7734 641898 -7498 642134
rect -7414 641898 -7178 642134
rect -7734 606218 -7498 606454
rect -7414 606218 -7178 606454
rect -7734 605898 -7498 606134
rect -7414 605898 -7178 606134
rect -7734 570218 -7498 570454
rect -7414 570218 -7178 570454
rect -7734 569898 -7498 570134
rect -7414 569898 -7178 570134
rect -7734 534218 -7498 534454
rect -7414 534218 -7178 534454
rect -7734 533898 -7498 534134
rect -7414 533898 -7178 534134
rect -7734 498218 -7498 498454
rect -7414 498218 -7178 498454
rect -7734 497898 -7498 498134
rect -7414 497898 -7178 498134
rect -7734 462218 -7498 462454
rect -7414 462218 -7178 462454
rect -7734 461898 -7498 462134
rect -7414 461898 -7178 462134
rect -7734 426218 -7498 426454
rect -7414 426218 -7178 426454
rect -7734 425898 -7498 426134
rect -7414 425898 -7178 426134
rect -7734 390218 -7498 390454
rect -7414 390218 -7178 390454
rect -7734 389898 -7498 390134
rect -7414 389898 -7178 390134
rect -7734 354218 -7498 354454
rect -7414 354218 -7178 354454
rect -7734 353898 -7498 354134
rect -7414 353898 -7178 354134
rect -7734 318218 -7498 318454
rect -7414 318218 -7178 318454
rect -7734 317898 -7498 318134
rect -7414 317898 -7178 318134
rect -7734 282218 -7498 282454
rect -7414 282218 -7178 282454
rect -7734 281898 -7498 282134
rect -7414 281898 -7178 282134
rect -7734 246218 -7498 246454
rect -7414 246218 -7178 246454
rect -7734 245898 -7498 246134
rect -7414 245898 -7178 246134
rect -7734 210218 -7498 210454
rect -7414 210218 -7178 210454
rect -7734 209898 -7498 210134
rect -7414 209898 -7178 210134
rect -7734 174218 -7498 174454
rect -7414 174218 -7178 174454
rect -7734 173898 -7498 174134
rect -7414 173898 -7178 174134
rect -7734 138218 -7498 138454
rect -7414 138218 -7178 138454
rect -7734 137898 -7498 138134
rect -7414 137898 -7178 138134
rect -7734 102218 -7498 102454
rect -7414 102218 -7178 102454
rect -7734 101898 -7498 102134
rect -7414 101898 -7178 102134
rect -7734 66218 -7498 66454
rect -7414 66218 -7178 66454
rect -7734 65898 -7498 66134
rect -7414 65898 -7178 66134
rect -7734 30218 -7498 30454
rect -7414 30218 -7178 30454
rect -7734 29898 -7498 30134
rect -7414 29898 -7178 30134
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 673718 -6538 673954
rect -6454 673718 -6218 673954
rect -6774 673398 -6538 673634
rect -6454 673398 -6218 673634
rect -6774 637718 -6538 637954
rect -6454 637718 -6218 637954
rect -6774 637398 -6538 637634
rect -6454 637398 -6218 637634
rect -6774 601718 -6538 601954
rect -6454 601718 -6218 601954
rect -6774 601398 -6538 601634
rect -6454 601398 -6218 601634
rect -6774 565718 -6538 565954
rect -6454 565718 -6218 565954
rect -6774 565398 -6538 565634
rect -6454 565398 -6218 565634
rect -6774 529718 -6538 529954
rect -6454 529718 -6218 529954
rect -6774 529398 -6538 529634
rect -6454 529398 -6218 529634
rect -6774 493718 -6538 493954
rect -6454 493718 -6218 493954
rect -6774 493398 -6538 493634
rect -6454 493398 -6218 493634
rect -6774 457718 -6538 457954
rect -6454 457718 -6218 457954
rect -6774 457398 -6538 457634
rect -6454 457398 -6218 457634
rect -6774 421718 -6538 421954
rect -6454 421718 -6218 421954
rect -6774 421398 -6538 421634
rect -6454 421398 -6218 421634
rect -6774 385718 -6538 385954
rect -6454 385718 -6218 385954
rect -6774 385398 -6538 385634
rect -6454 385398 -6218 385634
rect -6774 349718 -6538 349954
rect -6454 349718 -6218 349954
rect -6774 349398 -6538 349634
rect -6454 349398 -6218 349634
rect -6774 313718 -6538 313954
rect -6454 313718 -6218 313954
rect -6774 313398 -6538 313634
rect -6454 313398 -6218 313634
rect -6774 277718 -6538 277954
rect -6454 277718 -6218 277954
rect -6774 277398 -6538 277634
rect -6454 277398 -6218 277634
rect -6774 241718 -6538 241954
rect -6454 241718 -6218 241954
rect -6774 241398 -6538 241634
rect -6454 241398 -6218 241634
rect -6774 205718 -6538 205954
rect -6454 205718 -6218 205954
rect -6774 205398 -6538 205634
rect -6454 205398 -6218 205634
rect -6774 169718 -6538 169954
rect -6454 169718 -6218 169954
rect -6774 169398 -6538 169634
rect -6454 169398 -6218 169634
rect -6774 133718 -6538 133954
rect -6454 133718 -6218 133954
rect -6774 133398 -6538 133634
rect -6454 133398 -6218 133634
rect -6774 97718 -6538 97954
rect -6454 97718 -6218 97954
rect -6774 97398 -6538 97634
rect -6454 97398 -6218 97634
rect -6774 61718 -6538 61954
rect -6454 61718 -6218 61954
rect -6774 61398 -6538 61634
rect -6454 61398 -6218 61634
rect -6774 25718 -6538 25954
rect -6454 25718 -6218 25954
rect -6774 25398 -6538 25634
rect -6454 25398 -6218 25634
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 669218 -5578 669454
rect -5494 669218 -5258 669454
rect -5814 668898 -5578 669134
rect -5494 668898 -5258 669134
rect -5814 633218 -5578 633454
rect -5494 633218 -5258 633454
rect -5814 632898 -5578 633134
rect -5494 632898 -5258 633134
rect -5814 597218 -5578 597454
rect -5494 597218 -5258 597454
rect -5814 596898 -5578 597134
rect -5494 596898 -5258 597134
rect -5814 561218 -5578 561454
rect -5494 561218 -5258 561454
rect -5814 560898 -5578 561134
rect -5494 560898 -5258 561134
rect -5814 525218 -5578 525454
rect -5494 525218 -5258 525454
rect -5814 524898 -5578 525134
rect -5494 524898 -5258 525134
rect -5814 489218 -5578 489454
rect -5494 489218 -5258 489454
rect -5814 488898 -5578 489134
rect -5494 488898 -5258 489134
rect -5814 453218 -5578 453454
rect -5494 453218 -5258 453454
rect -5814 452898 -5578 453134
rect -5494 452898 -5258 453134
rect -5814 417218 -5578 417454
rect -5494 417218 -5258 417454
rect -5814 416898 -5578 417134
rect -5494 416898 -5258 417134
rect -5814 381218 -5578 381454
rect -5494 381218 -5258 381454
rect -5814 380898 -5578 381134
rect -5494 380898 -5258 381134
rect -5814 345218 -5578 345454
rect -5494 345218 -5258 345454
rect -5814 344898 -5578 345134
rect -5494 344898 -5258 345134
rect -5814 309218 -5578 309454
rect -5494 309218 -5258 309454
rect -5814 308898 -5578 309134
rect -5494 308898 -5258 309134
rect -5814 273218 -5578 273454
rect -5494 273218 -5258 273454
rect -5814 272898 -5578 273134
rect -5494 272898 -5258 273134
rect -5814 237218 -5578 237454
rect -5494 237218 -5258 237454
rect -5814 236898 -5578 237134
rect -5494 236898 -5258 237134
rect -5814 201218 -5578 201454
rect -5494 201218 -5258 201454
rect -5814 200898 -5578 201134
rect -5494 200898 -5258 201134
rect -5814 165218 -5578 165454
rect -5494 165218 -5258 165454
rect -5814 164898 -5578 165134
rect -5494 164898 -5258 165134
rect -5814 129218 -5578 129454
rect -5494 129218 -5258 129454
rect -5814 128898 -5578 129134
rect -5494 128898 -5258 129134
rect -5814 93218 -5578 93454
rect -5494 93218 -5258 93454
rect -5814 92898 -5578 93134
rect -5494 92898 -5258 93134
rect -5814 57218 -5578 57454
rect -5494 57218 -5258 57454
rect -5814 56898 -5578 57134
rect -5494 56898 -5258 57134
rect -5814 21218 -5578 21454
rect -5494 21218 -5258 21454
rect -5814 20898 -5578 21134
rect -5494 20898 -5258 21134
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 700718 -4618 700954
rect -4534 700718 -4298 700954
rect -4854 700398 -4618 700634
rect -4534 700398 -4298 700634
rect -4854 664718 -4618 664954
rect -4534 664718 -4298 664954
rect -4854 664398 -4618 664634
rect -4534 664398 -4298 664634
rect -4854 628718 -4618 628954
rect -4534 628718 -4298 628954
rect -4854 628398 -4618 628634
rect -4534 628398 -4298 628634
rect -4854 592718 -4618 592954
rect -4534 592718 -4298 592954
rect -4854 592398 -4618 592634
rect -4534 592398 -4298 592634
rect -4854 556718 -4618 556954
rect -4534 556718 -4298 556954
rect -4854 556398 -4618 556634
rect -4534 556398 -4298 556634
rect -4854 520718 -4618 520954
rect -4534 520718 -4298 520954
rect -4854 520398 -4618 520634
rect -4534 520398 -4298 520634
rect -4854 484718 -4618 484954
rect -4534 484718 -4298 484954
rect -4854 484398 -4618 484634
rect -4534 484398 -4298 484634
rect -4854 448718 -4618 448954
rect -4534 448718 -4298 448954
rect -4854 448398 -4618 448634
rect -4534 448398 -4298 448634
rect -4854 412718 -4618 412954
rect -4534 412718 -4298 412954
rect -4854 412398 -4618 412634
rect -4534 412398 -4298 412634
rect -4854 376718 -4618 376954
rect -4534 376718 -4298 376954
rect -4854 376398 -4618 376634
rect -4534 376398 -4298 376634
rect -4854 340718 -4618 340954
rect -4534 340718 -4298 340954
rect -4854 340398 -4618 340634
rect -4534 340398 -4298 340634
rect -4854 304718 -4618 304954
rect -4534 304718 -4298 304954
rect -4854 304398 -4618 304634
rect -4534 304398 -4298 304634
rect -4854 268718 -4618 268954
rect -4534 268718 -4298 268954
rect -4854 268398 -4618 268634
rect -4534 268398 -4298 268634
rect -4854 232718 -4618 232954
rect -4534 232718 -4298 232954
rect -4854 232398 -4618 232634
rect -4534 232398 -4298 232634
rect -4854 196718 -4618 196954
rect -4534 196718 -4298 196954
rect -4854 196398 -4618 196634
rect -4534 196398 -4298 196634
rect -4854 160718 -4618 160954
rect -4534 160718 -4298 160954
rect -4854 160398 -4618 160634
rect -4534 160398 -4298 160634
rect -4854 124718 -4618 124954
rect -4534 124718 -4298 124954
rect -4854 124398 -4618 124634
rect -4534 124398 -4298 124634
rect -4854 88718 -4618 88954
rect -4534 88718 -4298 88954
rect -4854 88398 -4618 88634
rect -4534 88398 -4298 88634
rect -4854 52718 -4618 52954
rect -4534 52718 -4298 52954
rect -4854 52398 -4618 52634
rect -4534 52398 -4298 52634
rect -4854 16718 -4618 16954
rect -4534 16718 -4298 16954
rect -4854 16398 -4618 16634
rect -4534 16398 -4298 16634
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 696218 -3658 696454
rect -3574 696218 -3338 696454
rect -3894 695898 -3658 696134
rect -3574 695898 -3338 696134
rect -3894 660218 -3658 660454
rect -3574 660218 -3338 660454
rect -3894 659898 -3658 660134
rect -3574 659898 -3338 660134
rect -3894 624218 -3658 624454
rect -3574 624218 -3338 624454
rect -3894 623898 -3658 624134
rect -3574 623898 -3338 624134
rect -3894 588218 -3658 588454
rect -3574 588218 -3338 588454
rect -3894 587898 -3658 588134
rect -3574 587898 -3338 588134
rect -3894 552218 -3658 552454
rect -3574 552218 -3338 552454
rect -3894 551898 -3658 552134
rect -3574 551898 -3338 552134
rect -3894 516218 -3658 516454
rect -3574 516218 -3338 516454
rect -3894 515898 -3658 516134
rect -3574 515898 -3338 516134
rect -3894 480218 -3658 480454
rect -3574 480218 -3338 480454
rect -3894 479898 -3658 480134
rect -3574 479898 -3338 480134
rect -3894 444218 -3658 444454
rect -3574 444218 -3338 444454
rect -3894 443898 -3658 444134
rect -3574 443898 -3338 444134
rect -3894 408218 -3658 408454
rect -3574 408218 -3338 408454
rect -3894 407898 -3658 408134
rect -3574 407898 -3338 408134
rect -3894 372218 -3658 372454
rect -3574 372218 -3338 372454
rect -3894 371898 -3658 372134
rect -3574 371898 -3338 372134
rect -3894 336218 -3658 336454
rect -3574 336218 -3338 336454
rect -3894 335898 -3658 336134
rect -3574 335898 -3338 336134
rect -3894 300218 -3658 300454
rect -3574 300218 -3338 300454
rect -3894 299898 -3658 300134
rect -3574 299898 -3338 300134
rect -3894 264218 -3658 264454
rect -3574 264218 -3338 264454
rect -3894 263898 -3658 264134
rect -3574 263898 -3338 264134
rect -3894 228218 -3658 228454
rect -3574 228218 -3338 228454
rect -3894 227898 -3658 228134
rect -3574 227898 -3338 228134
rect -3894 192218 -3658 192454
rect -3574 192218 -3338 192454
rect -3894 191898 -3658 192134
rect -3574 191898 -3338 192134
rect -3894 156218 -3658 156454
rect -3574 156218 -3338 156454
rect -3894 155898 -3658 156134
rect -3574 155898 -3338 156134
rect -3894 120218 -3658 120454
rect -3574 120218 -3338 120454
rect -3894 119898 -3658 120134
rect -3574 119898 -3338 120134
rect -3894 84218 -3658 84454
rect -3574 84218 -3338 84454
rect -3894 83898 -3658 84134
rect -3574 83898 -3338 84134
rect -3894 48218 -3658 48454
rect -3574 48218 -3338 48454
rect -3894 47898 -3658 48134
rect -3574 47898 -3338 48134
rect -3894 12218 -3658 12454
rect -3574 12218 -3338 12454
rect -3894 11898 -3658 12134
rect -3574 11898 -3338 12134
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 691718 -2698 691954
rect -2614 691718 -2378 691954
rect -2934 691398 -2698 691634
rect -2614 691398 -2378 691634
rect -2934 655718 -2698 655954
rect -2614 655718 -2378 655954
rect -2934 655398 -2698 655634
rect -2614 655398 -2378 655634
rect -2934 619718 -2698 619954
rect -2614 619718 -2378 619954
rect -2934 619398 -2698 619634
rect -2614 619398 -2378 619634
rect -2934 583718 -2698 583954
rect -2614 583718 -2378 583954
rect -2934 583398 -2698 583634
rect -2614 583398 -2378 583634
rect -2934 547718 -2698 547954
rect -2614 547718 -2378 547954
rect -2934 547398 -2698 547634
rect -2614 547398 -2378 547634
rect -2934 511718 -2698 511954
rect -2614 511718 -2378 511954
rect -2934 511398 -2698 511634
rect -2614 511398 -2378 511634
rect -2934 475718 -2698 475954
rect -2614 475718 -2378 475954
rect -2934 475398 -2698 475634
rect -2614 475398 -2378 475634
rect -2934 439718 -2698 439954
rect -2614 439718 -2378 439954
rect -2934 439398 -2698 439634
rect -2614 439398 -2378 439634
rect -2934 403718 -2698 403954
rect -2614 403718 -2378 403954
rect -2934 403398 -2698 403634
rect -2614 403398 -2378 403634
rect -2934 367718 -2698 367954
rect -2614 367718 -2378 367954
rect -2934 367398 -2698 367634
rect -2614 367398 -2378 367634
rect -2934 331718 -2698 331954
rect -2614 331718 -2378 331954
rect -2934 331398 -2698 331634
rect -2614 331398 -2378 331634
rect -2934 295718 -2698 295954
rect -2614 295718 -2378 295954
rect -2934 295398 -2698 295634
rect -2614 295398 -2378 295634
rect -2934 259718 -2698 259954
rect -2614 259718 -2378 259954
rect -2934 259398 -2698 259634
rect -2614 259398 -2378 259634
rect -2934 223718 -2698 223954
rect -2614 223718 -2378 223954
rect -2934 223398 -2698 223634
rect -2614 223398 -2378 223634
rect -2934 187718 -2698 187954
rect -2614 187718 -2378 187954
rect -2934 187398 -2698 187634
rect -2614 187398 -2378 187634
rect -2934 151718 -2698 151954
rect -2614 151718 -2378 151954
rect -2934 151398 -2698 151634
rect -2614 151398 -2378 151634
rect -2934 115718 -2698 115954
rect -2614 115718 -2378 115954
rect -2934 115398 -2698 115634
rect -2614 115398 -2378 115634
rect -2934 79718 -2698 79954
rect -2614 79718 -2378 79954
rect -2934 79398 -2698 79634
rect -2614 79398 -2378 79634
rect -2934 43718 -2698 43954
rect -2614 43718 -2378 43954
rect -2934 43398 -2698 43634
rect -2614 43398 -2378 43634
rect -2934 7718 -2698 7954
rect -2614 7718 -2378 7954
rect -2934 7398 -2698 7634
rect -2614 7398 -2378 7634
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 6326 705562 6562 705798
rect 6646 705562 6882 705798
rect 6326 705242 6562 705478
rect 6646 705242 6882 705478
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1542 6562 -1306
rect 6646 -1542 6882 -1306
rect 6326 -1862 6562 -1626
rect 6646 -1862 6882 -1626
rect 10826 706522 11062 706758
rect 11146 706522 11382 706758
rect 10826 706202 11062 706438
rect 11146 706202 11382 706438
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2502 11062 -2266
rect 11146 -2502 11382 -2266
rect 10826 -2822 11062 -2586
rect 11146 -2822 11382 -2586
rect 15326 707482 15562 707718
rect 15646 707482 15882 707718
rect 15326 707162 15562 707398
rect 15646 707162 15882 707398
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3462 15562 -3226
rect 15646 -3462 15882 -3226
rect 15326 -3782 15562 -3546
rect 15646 -3782 15882 -3546
rect 19826 708442 20062 708678
rect 20146 708442 20382 708678
rect 19826 708122 20062 708358
rect 20146 708122 20382 708358
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4422 20062 -4186
rect 20146 -4422 20382 -4186
rect 19826 -4742 20062 -4506
rect 20146 -4742 20382 -4506
rect 24326 709402 24562 709638
rect 24646 709402 24882 709638
rect 24326 709082 24562 709318
rect 24646 709082 24882 709318
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 24326 133718 24562 133954
rect 24646 133718 24882 133954
rect 24326 133398 24562 133634
rect 24646 133398 24882 133634
rect 24326 97718 24562 97954
rect 24646 97718 24882 97954
rect 24326 97398 24562 97634
rect 24646 97398 24882 97634
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5382 24562 -5146
rect 24646 -5382 24882 -5146
rect 24326 -5702 24562 -5466
rect 24646 -5702 24882 -5466
rect 28826 710362 29062 710598
rect 29146 710362 29382 710598
rect 28826 710042 29062 710278
rect 29146 710042 29382 710278
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 28826 138218 29062 138454
rect 29146 138218 29382 138454
rect 28826 137898 29062 138134
rect 29146 137898 29382 138134
rect 28826 102218 29062 102454
rect 29146 102218 29382 102454
rect 28826 101898 29062 102134
rect 29146 101898 29382 102134
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6342 29062 -6106
rect 29146 -6342 29382 -6106
rect 28826 -6662 29062 -6426
rect 29146 -6662 29382 -6426
rect 33326 711322 33562 711558
rect 33646 711322 33882 711558
rect 33326 711002 33562 711238
rect 33646 711002 33882 711238
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 33326 646718 33562 646954
rect 33646 646718 33882 646954
rect 33326 646398 33562 646634
rect 33646 646398 33882 646634
rect 33326 610718 33562 610954
rect 33646 610718 33882 610954
rect 33326 610398 33562 610634
rect 33646 610398 33882 610634
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 33326 142718 33562 142954
rect 33646 142718 33882 142954
rect 33326 142398 33562 142634
rect 33646 142398 33882 142634
rect 33326 106718 33562 106954
rect 33646 106718 33882 106954
rect 33326 106398 33562 106634
rect 33646 106398 33882 106634
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7302 33562 -7066
rect 33646 -7302 33882 -7066
rect 33326 -7622 33562 -7386
rect 33646 -7622 33882 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 42326 705562 42562 705798
rect 42646 705562 42882 705798
rect 42326 705242 42562 705478
rect 42646 705242 42882 705478
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 42326 655718 42562 655954
rect 42646 655718 42882 655954
rect 42326 655398 42562 655634
rect 42646 655398 42882 655634
rect 42326 619718 42562 619954
rect 42646 619718 42882 619954
rect 42326 619398 42562 619634
rect 42646 619398 42882 619634
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 46826 706522 47062 706758
rect 47146 706522 47382 706758
rect 46826 706202 47062 706438
rect 47146 706202 47382 706438
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 46826 660218 47062 660454
rect 47146 660218 47382 660454
rect 46826 659898 47062 660134
rect 47146 659898 47382 660134
rect 46826 624218 47062 624454
rect 47146 624218 47382 624454
rect 46826 623898 47062 624134
rect 47146 623898 47382 624134
rect 46826 588218 47062 588454
rect 47146 588218 47382 588454
rect 46826 587898 47062 588134
rect 47146 587898 47382 588134
rect 46826 552218 47062 552454
rect 47146 552218 47382 552454
rect 46826 551898 47062 552134
rect 47146 551898 47382 552134
rect 46826 516218 47062 516454
rect 47146 516218 47382 516454
rect 46826 515898 47062 516134
rect 47146 515898 47382 516134
rect 46826 480218 47062 480454
rect 47146 480218 47382 480454
rect 46826 479898 47062 480134
rect 47146 479898 47382 480134
rect 46826 444218 47062 444454
rect 47146 444218 47382 444454
rect 46826 443898 47062 444134
rect 47146 443898 47382 444134
rect 46826 408218 47062 408454
rect 47146 408218 47382 408454
rect 46826 407898 47062 408134
rect 47146 407898 47382 408134
rect 46826 372218 47062 372454
rect 47146 372218 47382 372454
rect 46826 371898 47062 372134
rect 47146 371898 47382 372134
rect 46826 336218 47062 336454
rect 47146 336218 47382 336454
rect 46826 335898 47062 336134
rect 47146 335898 47382 336134
rect 46826 300218 47062 300454
rect 47146 300218 47382 300454
rect 46826 299898 47062 300134
rect 47146 299898 47382 300134
rect 46826 264218 47062 264454
rect 47146 264218 47382 264454
rect 46826 263898 47062 264134
rect 47146 263898 47382 264134
rect 51326 707482 51562 707718
rect 51646 707482 51882 707718
rect 51326 707162 51562 707398
rect 51646 707162 51882 707398
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 51326 664718 51562 664954
rect 51646 664718 51882 664954
rect 51326 664398 51562 664634
rect 51646 664398 51882 664634
rect 51326 628718 51562 628954
rect 51646 628718 51882 628954
rect 51326 628398 51562 628634
rect 51646 628398 51882 628634
rect 51326 592718 51562 592954
rect 51646 592718 51882 592954
rect 51326 592398 51562 592634
rect 51646 592398 51882 592634
rect 51326 556718 51562 556954
rect 51646 556718 51882 556954
rect 51326 556398 51562 556634
rect 51646 556398 51882 556634
rect 51326 520718 51562 520954
rect 51646 520718 51882 520954
rect 51326 520398 51562 520634
rect 51646 520398 51882 520634
rect 51326 484718 51562 484954
rect 51646 484718 51882 484954
rect 51326 484398 51562 484634
rect 51646 484398 51882 484634
rect 51326 448718 51562 448954
rect 51646 448718 51882 448954
rect 51326 448398 51562 448634
rect 51646 448398 51882 448634
rect 51326 412718 51562 412954
rect 51646 412718 51882 412954
rect 51326 412398 51562 412634
rect 51646 412398 51882 412634
rect 51326 376718 51562 376954
rect 51646 376718 51882 376954
rect 51326 376398 51562 376634
rect 51646 376398 51882 376634
rect 51326 340718 51562 340954
rect 51646 340718 51882 340954
rect 51326 340398 51562 340634
rect 51646 340398 51882 340634
rect 51326 304718 51562 304954
rect 51646 304718 51882 304954
rect 51326 304398 51562 304634
rect 51646 304398 51882 304634
rect 51326 268718 51562 268954
rect 51646 268718 51882 268954
rect 51326 268398 51562 268634
rect 51646 268398 51882 268634
rect 55826 708442 56062 708678
rect 56146 708442 56382 708678
rect 55826 708122 56062 708358
rect 56146 708122 56382 708358
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 60326 709402 60562 709638
rect 60646 709402 60882 709638
rect 60326 709082 60562 709318
rect 60646 709082 60882 709318
rect 60326 673718 60562 673954
rect 60646 673718 60882 673954
rect 60326 673398 60562 673634
rect 60646 673398 60882 673634
rect 60326 637718 60562 637954
rect 60646 637718 60882 637954
rect 60326 637398 60562 637634
rect 60646 637398 60882 637634
rect 60326 601718 60562 601954
rect 60646 601718 60882 601954
rect 60326 601398 60562 601634
rect 60646 601398 60882 601634
rect 60326 565718 60562 565954
rect 60646 565718 60882 565954
rect 60326 565398 60562 565634
rect 60646 565398 60882 565634
rect 60326 529718 60562 529954
rect 60646 529718 60882 529954
rect 60326 529398 60562 529634
rect 60646 529398 60882 529634
rect 60326 493718 60562 493954
rect 60646 493718 60882 493954
rect 60326 493398 60562 493634
rect 60646 493398 60882 493634
rect 60326 457718 60562 457954
rect 60646 457718 60882 457954
rect 60326 457398 60562 457634
rect 60646 457398 60882 457634
rect 60326 421718 60562 421954
rect 60646 421718 60882 421954
rect 60326 421398 60562 421634
rect 60646 421398 60882 421634
rect 60326 385718 60562 385954
rect 60646 385718 60882 385954
rect 60326 385398 60562 385634
rect 60646 385398 60882 385634
rect 60326 349718 60562 349954
rect 60646 349718 60882 349954
rect 60326 349398 60562 349634
rect 60646 349398 60882 349634
rect 60326 313718 60562 313954
rect 60646 313718 60882 313954
rect 60326 313398 60562 313634
rect 60646 313398 60882 313634
rect 60326 277718 60562 277954
rect 60646 277718 60882 277954
rect 60326 277398 60562 277634
rect 60646 277398 60882 277634
rect 64826 710362 65062 710598
rect 65146 710362 65382 710598
rect 64826 710042 65062 710278
rect 65146 710042 65382 710278
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 64826 642218 65062 642454
rect 65146 642218 65382 642454
rect 64826 641898 65062 642134
rect 65146 641898 65382 642134
rect 64826 606218 65062 606454
rect 65146 606218 65382 606454
rect 64826 605898 65062 606134
rect 65146 605898 65382 606134
rect 64826 570218 65062 570454
rect 65146 570218 65382 570454
rect 64826 569898 65062 570134
rect 65146 569898 65382 570134
rect 64826 534218 65062 534454
rect 65146 534218 65382 534454
rect 64826 533898 65062 534134
rect 65146 533898 65382 534134
rect 64826 498218 65062 498454
rect 65146 498218 65382 498454
rect 64826 497898 65062 498134
rect 65146 497898 65382 498134
rect 64826 462218 65062 462454
rect 65146 462218 65382 462454
rect 64826 461898 65062 462134
rect 65146 461898 65382 462134
rect 64826 426218 65062 426454
rect 65146 426218 65382 426454
rect 64826 425898 65062 426134
rect 65146 425898 65382 426134
rect 64826 390218 65062 390454
rect 65146 390218 65382 390454
rect 64826 389898 65062 390134
rect 65146 389898 65382 390134
rect 64826 354218 65062 354454
rect 65146 354218 65382 354454
rect 64826 353898 65062 354134
rect 65146 353898 65382 354134
rect 64826 318218 65062 318454
rect 65146 318218 65382 318454
rect 64826 317898 65062 318134
rect 65146 317898 65382 318134
rect 64826 282218 65062 282454
rect 65146 282218 65382 282454
rect 64826 281898 65062 282134
rect 65146 281898 65382 282134
rect 69326 711322 69562 711558
rect 69646 711322 69882 711558
rect 69326 711002 69562 711238
rect 69646 711002 69882 711238
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 69326 646718 69562 646954
rect 69646 646718 69882 646954
rect 69326 646398 69562 646634
rect 69646 646398 69882 646634
rect 69326 610718 69562 610954
rect 69646 610718 69882 610954
rect 69326 610398 69562 610634
rect 69646 610398 69882 610634
rect 69326 574718 69562 574954
rect 69646 574718 69882 574954
rect 69326 574398 69562 574634
rect 69646 574398 69882 574634
rect 69326 538718 69562 538954
rect 69646 538718 69882 538954
rect 69326 538398 69562 538634
rect 69646 538398 69882 538634
rect 69326 502718 69562 502954
rect 69646 502718 69882 502954
rect 69326 502398 69562 502634
rect 69646 502398 69882 502634
rect 69326 466718 69562 466954
rect 69646 466718 69882 466954
rect 69326 466398 69562 466634
rect 69646 466398 69882 466634
rect 69326 430718 69562 430954
rect 69646 430718 69882 430954
rect 69326 430398 69562 430634
rect 69646 430398 69882 430634
rect 69326 394718 69562 394954
rect 69646 394718 69882 394954
rect 69326 394398 69562 394634
rect 69646 394398 69882 394634
rect 69326 358718 69562 358954
rect 69646 358718 69882 358954
rect 69326 358398 69562 358634
rect 69646 358398 69882 358634
rect 69326 322718 69562 322954
rect 69646 322718 69882 322954
rect 69326 322398 69562 322634
rect 69646 322398 69882 322634
rect 69326 286718 69562 286954
rect 69646 286718 69882 286954
rect 69326 286398 69562 286634
rect 69646 286398 69882 286634
rect 69326 250718 69562 250954
rect 69646 250718 69882 250954
rect 69326 250398 69562 250634
rect 69646 250398 69882 250634
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 78326 705562 78562 705798
rect 78646 705562 78882 705798
rect 78326 705242 78562 705478
rect 78646 705242 78882 705478
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 78326 655718 78562 655954
rect 78646 655718 78882 655954
rect 78326 655398 78562 655634
rect 78646 655398 78882 655634
rect 78326 619718 78562 619954
rect 78646 619718 78882 619954
rect 78326 619398 78562 619634
rect 78646 619398 78882 619634
rect 78326 583718 78562 583954
rect 78646 583718 78882 583954
rect 78326 583398 78562 583634
rect 78646 583398 78882 583634
rect 78326 547718 78562 547954
rect 78646 547718 78882 547954
rect 78326 547398 78562 547634
rect 78646 547398 78882 547634
rect 78326 511718 78562 511954
rect 78646 511718 78882 511954
rect 78326 511398 78562 511634
rect 78646 511398 78882 511634
rect 78326 475718 78562 475954
rect 78646 475718 78882 475954
rect 78326 475398 78562 475634
rect 78646 475398 78882 475634
rect 78326 439718 78562 439954
rect 78646 439718 78882 439954
rect 78326 439398 78562 439634
rect 78646 439398 78882 439634
rect 78326 403718 78562 403954
rect 78646 403718 78882 403954
rect 78326 403398 78562 403634
rect 78646 403398 78882 403634
rect 78326 367718 78562 367954
rect 78646 367718 78882 367954
rect 78326 367398 78562 367634
rect 78646 367398 78882 367634
rect 78326 331718 78562 331954
rect 78646 331718 78882 331954
rect 78326 331398 78562 331634
rect 78646 331398 78882 331634
rect 78326 295718 78562 295954
rect 78646 295718 78882 295954
rect 78326 295398 78562 295634
rect 78646 295398 78882 295634
rect 78326 259718 78562 259954
rect 78646 259718 78882 259954
rect 78326 259398 78562 259634
rect 78646 259398 78882 259634
rect 82826 706522 83062 706758
rect 83146 706522 83382 706758
rect 82826 706202 83062 706438
rect 83146 706202 83382 706438
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 82826 660218 83062 660454
rect 83146 660218 83382 660454
rect 82826 659898 83062 660134
rect 83146 659898 83382 660134
rect 82826 624218 83062 624454
rect 83146 624218 83382 624454
rect 82826 623898 83062 624134
rect 83146 623898 83382 624134
rect 82826 588218 83062 588454
rect 83146 588218 83382 588454
rect 82826 587898 83062 588134
rect 83146 587898 83382 588134
rect 82826 552218 83062 552454
rect 83146 552218 83382 552454
rect 82826 551898 83062 552134
rect 83146 551898 83382 552134
rect 82826 516218 83062 516454
rect 83146 516218 83382 516454
rect 82826 515898 83062 516134
rect 83146 515898 83382 516134
rect 82826 480218 83062 480454
rect 83146 480218 83382 480454
rect 82826 479898 83062 480134
rect 83146 479898 83382 480134
rect 82826 444218 83062 444454
rect 83146 444218 83382 444454
rect 82826 443898 83062 444134
rect 83146 443898 83382 444134
rect 82826 408218 83062 408454
rect 83146 408218 83382 408454
rect 82826 407898 83062 408134
rect 83146 407898 83382 408134
rect 82826 372218 83062 372454
rect 83146 372218 83382 372454
rect 82826 371898 83062 372134
rect 83146 371898 83382 372134
rect 82826 336218 83062 336454
rect 83146 336218 83382 336454
rect 82826 335898 83062 336134
rect 83146 335898 83382 336134
rect 82826 300218 83062 300454
rect 83146 300218 83382 300454
rect 82826 299898 83062 300134
rect 83146 299898 83382 300134
rect 82826 264218 83062 264454
rect 83146 264218 83382 264454
rect 82826 263898 83062 264134
rect 83146 263898 83382 264134
rect 87326 707482 87562 707718
rect 87646 707482 87882 707718
rect 87326 707162 87562 707398
rect 87646 707162 87882 707398
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 87326 664718 87562 664954
rect 87646 664718 87882 664954
rect 87326 664398 87562 664634
rect 87646 664398 87882 664634
rect 87326 628718 87562 628954
rect 87646 628718 87882 628954
rect 87326 628398 87562 628634
rect 87646 628398 87882 628634
rect 87326 592718 87562 592954
rect 87646 592718 87882 592954
rect 87326 592398 87562 592634
rect 87646 592398 87882 592634
rect 87326 556718 87562 556954
rect 87646 556718 87882 556954
rect 87326 556398 87562 556634
rect 87646 556398 87882 556634
rect 87326 520718 87562 520954
rect 87646 520718 87882 520954
rect 87326 520398 87562 520634
rect 87646 520398 87882 520634
rect 87326 484718 87562 484954
rect 87646 484718 87882 484954
rect 87326 484398 87562 484634
rect 87646 484398 87882 484634
rect 87326 448718 87562 448954
rect 87646 448718 87882 448954
rect 87326 448398 87562 448634
rect 87646 448398 87882 448634
rect 87326 412718 87562 412954
rect 87646 412718 87882 412954
rect 87326 412398 87562 412634
rect 87646 412398 87882 412634
rect 87326 376718 87562 376954
rect 87646 376718 87882 376954
rect 87326 376398 87562 376634
rect 87646 376398 87882 376634
rect 87326 340718 87562 340954
rect 87646 340718 87882 340954
rect 87326 340398 87562 340634
rect 87646 340398 87882 340634
rect 87326 304718 87562 304954
rect 87646 304718 87882 304954
rect 87326 304398 87562 304634
rect 87646 304398 87882 304634
rect 87326 268718 87562 268954
rect 87646 268718 87882 268954
rect 87326 268398 87562 268634
rect 87646 268398 87882 268634
rect 91826 708442 92062 708678
rect 92146 708442 92382 708678
rect 91826 708122 92062 708358
rect 92146 708122 92382 708358
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 96326 709402 96562 709638
rect 96646 709402 96882 709638
rect 96326 709082 96562 709318
rect 96646 709082 96882 709318
rect 96326 673718 96562 673954
rect 96646 673718 96882 673954
rect 96326 673398 96562 673634
rect 96646 673398 96882 673634
rect 96326 637718 96562 637954
rect 96646 637718 96882 637954
rect 96326 637398 96562 637634
rect 96646 637398 96882 637634
rect 96326 601718 96562 601954
rect 96646 601718 96882 601954
rect 96326 601398 96562 601634
rect 96646 601398 96882 601634
rect 96326 565718 96562 565954
rect 96646 565718 96882 565954
rect 96326 565398 96562 565634
rect 96646 565398 96882 565634
rect 96326 529718 96562 529954
rect 96646 529718 96882 529954
rect 96326 529398 96562 529634
rect 96646 529398 96882 529634
rect 96326 493718 96562 493954
rect 96646 493718 96882 493954
rect 96326 493398 96562 493634
rect 96646 493398 96882 493634
rect 96326 457718 96562 457954
rect 96646 457718 96882 457954
rect 96326 457398 96562 457634
rect 96646 457398 96882 457634
rect 96326 421718 96562 421954
rect 96646 421718 96882 421954
rect 96326 421398 96562 421634
rect 96646 421398 96882 421634
rect 96326 385718 96562 385954
rect 96646 385718 96882 385954
rect 96326 385398 96562 385634
rect 96646 385398 96882 385634
rect 96326 349718 96562 349954
rect 96646 349718 96882 349954
rect 96326 349398 96562 349634
rect 96646 349398 96882 349634
rect 96326 313718 96562 313954
rect 96646 313718 96882 313954
rect 96326 313398 96562 313634
rect 96646 313398 96882 313634
rect 96326 277718 96562 277954
rect 96646 277718 96882 277954
rect 96326 277398 96562 277634
rect 96646 277398 96882 277634
rect 100826 710362 101062 710598
rect 101146 710362 101382 710598
rect 100826 710042 101062 710278
rect 101146 710042 101382 710278
rect 100826 678218 101062 678454
rect 101146 678218 101382 678454
rect 100826 677898 101062 678134
rect 101146 677898 101382 678134
rect 100826 642218 101062 642454
rect 101146 642218 101382 642454
rect 100826 641898 101062 642134
rect 101146 641898 101382 642134
rect 100826 606218 101062 606454
rect 101146 606218 101382 606454
rect 100826 605898 101062 606134
rect 101146 605898 101382 606134
rect 100826 570218 101062 570454
rect 101146 570218 101382 570454
rect 100826 569898 101062 570134
rect 101146 569898 101382 570134
rect 100826 534218 101062 534454
rect 101146 534218 101382 534454
rect 100826 533898 101062 534134
rect 101146 533898 101382 534134
rect 100826 498218 101062 498454
rect 101146 498218 101382 498454
rect 100826 497898 101062 498134
rect 101146 497898 101382 498134
rect 100826 462218 101062 462454
rect 101146 462218 101382 462454
rect 100826 461898 101062 462134
rect 101146 461898 101382 462134
rect 100826 426218 101062 426454
rect 101146 426218 101382 426454
rect 100826 425898 101062 426134
rect 101146 425898 101382 426134
rect 100826 390218 101062 390454
rect 101146 390218 101382 390454
rect 100826 389898 101062 390134
rect 101146 389898 101382 390134
rect 100826 354218 101062 354454
rect 101146 354218 101382 354454
rect 100826 353898 101062 354134
rect 101146 353898 101382 354134
rect 100826 318218 101062 318454
rect 101146 318218 101382 318454
rect 100826 317898 101062 318134
rect 101146 317898 101382 318134
rect 100826 282218 101062 282454
rect 101146 282218 101382 282454
rect 100826 281898 101062 282134
rect 101146 281898 101382 282134
rect 105326 711322 105562 711558
rect 105646 711322 105882 711558
rect 105326 711002 105562 711238
rect 105646 711002 105882 711238
rect 105326 682718 105562 682954
rect 105646 682718 105882 682954
rect 105326 682398 105562 682634
rect 105646 682398 105882 682634
rect 105326 646718 105562 646954
rect 105646 646718 105882 646954
rect 105326 646398 105562 646634
rect 105646 646398 105882 646634
rect 105326 610718 105562 610954
rect 105646 610718 105882 610954
rect 105326 610398 105562 610634
rect 105646 610398 105882 610634
rect 105326 574718 105562 574954
rect 105646 574718 105882 574954
rect 105326 574398 105562 574634
rect 105646 574398 105882 574634
rect 105326 538718 105562 538954
rect 105646 538718 105882 538954
rect 105326 538398 105562 538634
rect 105646 538398 105882 538634
rect 105326 502718 105562 502954
rect 105646 502718 105882 502954
rect 105326 502398 105562 502634
rect 105646 502398 105882 502634
rect 105326 466718 105562 466954
rect 105646 466718 105882 466954
rect 105326 466398 105562 466634
rect 105646 466398 105882 466634
rect 105326 430718 105562 430954
rect 105646 430718 105882 430954
rect 105326 430398 105562 430634
rect 105646 430398 105882 430634
rect 105326 394718 105562 394954
rect 105646 394718 105882 394954
rect 105326 394398 105562 394634
rect 105646 394398 105882 394634
rect 105326 358718 105562 358954
rect 105646 358718 105882 358954
rect 105326 358398 105562 358634
rect 105646 358398 105882 358634
rect 105326 322718 105562 322954
rect 105646 322718 105882 322954
rect 105326 322398 105562 322634
rect 105646 322398 105882 322634
rect 105326 286718 105562 286954
rect 105646 286718 105882 286954
rect 105326 286398 105562 286634
rect 105646 286398 105882 286634
rect 105326 250718 105562 250954
rect 105646 250718 105882 250954
rect 105326 250398 105562 250634
rect 105646 250398 105882 250634
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 114326 705562 114562 705798
rect 114646 705562 114882 705798
rect 114326 705242 114562 705478
rect 114646 705242 114882 705478
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 114326 655718 114562 655954
rect 114646 655718 114882 655954
rect 114326 655398 114562 655634
rect 114646 655398 114882 655634
rect 114326 619718 114562 619954
rect 114646 619718 114882 619954
rect 114326 619398 114562 619634
rect 114646 619398 114882 619634
rect 114326 583718 114562 583954
rect 114646 583718 114882 583954
rect 114326 583398 114562 583634
rect 114646 583398 114882 583634
rect 114326 547718 114562 547954
rect 114646 547718 114882 547954
rect 114326 547398 114562 547634
rect 114646 547398 114882 547634
rect 114326 511718 114562 511954
rect 114646 511718 114882 511954
rect 114326 511398 114562 511634
rect 114646 511398 114882 511634
rect 114326 475718 114562 475954
rect 114646 475718 114882 475954
rect 114326 475398 114562 475634
rect 114646 475398 114882 475634
rect 114326 439718 114562 439954
rect 114646 439718 114882 439954
rect 114326 439398 114562 439634
rect 114646 439398 114882 439634
rect 114326 403718 114562 403954
rect 114646 403718 114882 403954
rect 114326 403398 114562 403634
rect 114646 403398 114882 403634
rect 114326 367718 114562 367954
rect 114646 367718 114882 367954
rect 114326 367398 114562 367634
rect 114646 367398 114882 367634
rect 114326 331718 114562 331954
rect 114646 331718 114882 331954
rect 114326 331398 114562 331634
rect 114646 331398 114882 331634
rect 114326 295718 114562 295954
rect 114646 295718 114882 295954
rect 114326 295398 114562 295634
rect 114646 295398 114882 295634
rect 114326 259718 114562 259954
rect 114646 259718 114882 259954
rect 114326 259398 114562 259634
rect 114646 259398 114882 259634
rect 118826 706522 119062 706758
rect 119146 706522 119382 706758
rect 118826 706202 119062 706438
rect 119146 706202 119382 706438
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 118826 660218 119062 660454
rect 119146 660218 119382 660454
rect 118826 659898 119062 660134
rect 119146 659898 119382 660134
rect 118826 624218 119062 624454
rect 119146 624218 119382 624454
rect 118826 623898 119062 624134
rect 119146 623898 119382 624134
rect 118826 588218 119062 588454
rect 119146 588218 119382 588454
rect 118826 587898 119062 588134
rect 119146 587898 119382 588134
rect 118826 552218 119062 552454
rect 119146 552218 119382 552454
rect 118826 551898 119062 552134
rect 119146 551898 119382 552134
rect 118826 516218 119062 516454
rect 119146 516218 119382 516454
rect 118826 515898 119062 516134
rect 119146 515898 119382 516134
rect 118826 480218 119062 480454
rect 119146 480218 119382 480454
rect 118826 479898 119062 480134
rect 119146 479898 119382 480134
rect 118826 444218 119062 444454
rect 119146 444218 119382 444454
rect 118826 443898 119062 444134
rect 119146 443898 119382 444134
rect 118826 408218 119062 408454
rect 119146 408218 119382 408454
rect 118826 407898 119062 408134
rect 119146 407898 119382 408134
rect 118826 372218 119062 372454
rect 119146 372218 119382 372454
rect 118826 371898 119062 372134
rect 119146 371898 119382 372134
rect 118826 336218 119062 336454
rect 119146 336218 119382 336454
rect 118826 335898 119062 336134
rect 119146 335898 119382 336134
rect 118826 300218 119062 300454
rect 119146 300218 119382 300454
rect 118826 299898 119062 300134
rect 119146 299898 119382 300134
rect 118826 264218 119062 264454
rect 119146 264218 119382 264454
rect 118826 263898 119062 264134
rect 119146 263898 119382 264134
rect 123326 707482 123562 707718
rect 123646 707482 123882 707718
rect 123326 707162 123562 707398
rect 123646 707162 123882 707398
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 123326 664718 123562 664954
rect 123646 664718 123882 664954
rect 123326 664398 123562 664634
rect 123646 664398 123882 664634
rect 123326 628718 123562 628954
rect 123646 628718 123882 628954
rect 123326 628398 123562 628634
rect 123646 628398 123882 628634
rect 123326 592718 123562 592954
rect 123646 592718 123882 592954
rect 123326 592398 123562 592634
rect 123646 592398 123882 592634
rect 123326 556718 123562 556954
rect 123646 556718 123882 556954
rect 123326 556398 123562 556634
rect 123646 556398 123882 556634
rect 123326 520718 123562 520954
rect 123646 520718 123882 520954
rect 123326 520398 123562 520634
rect 123646 520398 123882 520634
rect 123326 484718 123562 484954
rect 123646 484718 123882 484954
rect 123326 484398 123562 484634
rect 123646 484398 123882 484634
rect 123326 448718 123562 448954
rect 123646 448718 123882 448954
rect 123326 448398 123562 448634
rect 123646 448398 123882 448634
rect 123326 412718 123562 412954
rect 123646 412718 123882 412954
rect 123326 412398 123562 412634
rect 123646 412398 123882 412634
rect 123326 376718 123562 376954
rect 123646 376718 123882 376954
rect 123326 376398 123562 376634
rect 123646 376398 123882 376634
rect 123326 340718 123562 340954
rect 123646 340718 123882 340954
rect 123326 340398 123562 340634
rect 123646 340398 123882 340634
rect 123326 304718 123562 304954
rect 123646 304718 123882 304954
rect 123326 304398 123562 304634
rect 123646 304398 123882 304634
rect 123326 268718 123562 268954
rect 123646 268718 123882 268954
rect 123326 268398 123562 268634
rect 123646 268398 123882 268634
rect 127826 708442 128062 708678
rect 128146 708442 128382 708678
rect 127826 708122 128062 708358
rect 128146 708122 128382 708358
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 132326 709402 132562 709638
rect 132646 709402 132882 709638
rect 132326 709082 132562 709318
rect 132646 709082 132882 709318
rect 132326 673718 132562 673954
rect 132646 673718 132882 673954
rect 132326 673398 132562 673634
rect 132646 673398 132882 673634
rect 132326 637718 132562 637954
rect 132646 637718 132882 637954
rect 132326 637398 132562 637634
rect 132646 637398 132882 637634
rect 132326 601718 132562 601954
rect 132646 601718 132882 601954
rect 132326 601398 132562 601634
rect 132646 601398 132882 601634
rect 132326 565718 132562 565954
rect 132646 565718 132882 565954
rect 132326 565398 132562 565634
rect 132646 565398 132882 565634
rect 132326 529718 132562 529954
rect 132646 529718 132882 529954
rect 132326 529398 132562 529634
rect 132646 529398 132882 529634
rect 132326 493718 132562 493954
rect 132646 493718 132882 493954
rect 132326 493398 132562 493634
rect 132646 493398 132882 493634
rect 132326 457718 132562 457954
rect 132646 457718 132882 457954
rect 132326 457398 132562 457634
rect 132646 457398 132882 457634
rect 132326 421718 132562 421954
rect 132646 421718 132882 421954
rect 132326 421398 132562 421634
rect 132646 421398 132882 421634
rect 132326 385718 132562 385954
rect 132646 385718 132882 385954
rect 132326 385398 132562 385634
rect 132646 385398 132882 385634
rect 132326 349718 132562 349954
rect 132646 349718 132882 349954
rect 132326 349398 132562 349634
rect 132646 349398 132882 349634
rect 132326 313718 132562 313954
rect 132646 313718 132882 313954
rect 132326 313398 132562 313634
rect 132646 313398 132882 313634
rect 132326 277718 132562 277954
rect 132646 277718 132882 277954
rect 132326 277398 132562 277634
rect 132646 277398 132882 277634
rect 136826 710362 137062 710598
rect 137146 710362 137382 710598
rect 136826 710042 137062 710278
rect 137146 710042 137382 710278
rect 136826 678218 137062 678454
rect 137146 678218 137382 678454
rect 136826 677898 137062 678134
rect 137146 677898 137382 678134
rect 136826 642218 137062 642454
rect 137146 642218 137382 642454
rect 136826 641898 137062 642134
rect 137146 641898 137382 642134
rect 136826 606218 137062 606454
rect 137146 606218 137382 606454
rect 136826 605898 137062 606134
rect 137146 605898 137382 606134
rect 136826 570218 137062 570454
rect 137146 570218 137382 570454
rect 136826 569898 137062 570134
rect 137146 569898 137382 570134
rect 136826 534218 137062 534454
rect 137146 534218 137382 534454
rect 136826 533898 137062 534134
rect 137146 533898 137382 534134
rect 136826 498218 137062 498454
rect 137146 498218 137382 498454
rect 136826 497898 137062 498134
rect 137146 497898 137382 498134
rect 136826 462218 137062 462454
rect 137146 462218 137382 462454
rect 136826 461898 137062 462134
rect 137146 461898 137382 462134
rect 136826 426218 137062 426454
rect 137146 426218 137382 426454
rect 136826 425898 137062 426134
rect 137146 425898 137382 426134
rect 136826 390218 137062 390454
rect 137146 390218 137382 390454
rect 136826 389898 137062 390134
rect 137146 389898 137382 390134
rect 136826 354218 137062 354454
rect 137146 354218 137382 354454
rect 136826 353898 137062 354134
rect 137146 353898 137382 354134
rect 136826 318218 137062 318454
rect 137146 318218 137382 318454
rect 136826 317898 137062 318134
rect 137146 317898 137382 318134
rect 136826 282218 137062 282454
rect 137146 282218 137382 282454
rect 136826 281898 137062 282134
rect 137146 281898 137382 282134
rect 141326 711322 141562 711558
rect 141646 711322 141882 711558
rect 141326 711002 141562 711238
rect 141646 711002 141882 711238
rect 141326 682718 141562 682954
rect 141646 682718 141882 682954
rect 141326 682398 141562 682634
rect 141646 682398 141882 682634
rect 141326 646718 141562 646954
rect 141646 646718 141882 646954
rect 141326 646398 141562 646634
rect 141646 646398 141882 646634
rect 141326 610718 141562 610954
rect 141646 610718 141882 610954
rect 141326 610398 141562 610634
rect 141646 610398 141882 610634
rect 141326 574718 141562 574954
rect 141646 574718 141882 574954
rect 141326 574398 141562 574634
rect 141646 574398 141882 574634
rect 141326 538718 141562 538954
rect 141646 538718 141882 538954
rect 141326 538398 141562 538634
rect 141646 538398 141882 538634
rect 141326 502718 141562 502954
rect 141646 502718 141882 502954
rect 141326 502398 141562 502634
rect 141646 502398 141882 502634
rect 141326 466718 141562 466954
rect 141646 466718 141882 466954
rect 141326 466398 141562 466634
rect 141646 466398 141882 466634
rect 141326 430718 141562 430954
rect 141646 430718 141882 430954
rect 141326 430398 141562 430634
rect 141646 430398 141882 430634
rect 141326 394718 141562 394954
rect 141646 394718 141882 394954
rect 141326 394398 141562 394634
rect 141646 394398 141882 394634
rect 141326 358718 141562 358954
rect 141646 358718 141882 358954
rect 141326 358398 141562 358634
rect 141646 358398 141882 358634
rect 141326 322718 141562 322954
rect 141646 322718 141882 322954
rect 141326 322398 141562 322634
rect 141646 322398 141882 322634
rect 141326 286718 141562 286954
rect 141646 286718 141882 286954
rect 141326 286398 141562 286634
rect 141646 286398 141882 286634
rect 141326 250718 141562 250954
rect 141646 250718 141882 250954
rect 141326 250398 141562 250634
rect 141646 250398 141882 250634
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 150326 705562 150562 705798
rect 150646 705562 150882 705798
rect 150326 705242 150562 705478
rect 150646 705242 150882 705478
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 150326 655718 150562 655954
rect 150646 655718 150882 655954
rect 150326 655398 150562 655634
rect 150646 655398 150882 655634
rect 150326 619718 150562 619954
rect 150646 619718 150882 619954
rect 150326 619398 150562 619634
rect 150646 619398 150882 619634
rect 150326 583718 150562 583954
rect 150646 583718 150882 583954
rect 150326 583398 150562 583634
rect 150646 583398 150882 583634
rect 150326 547718 150562 547954
rect 150646 547718 150882 547954
rect 150326 547398 150562 547634
rect 150646 547398 150882 547634
rect 150326 511718 150562 511954
rect 150646 511718 150882 511954
rect 150326 511398 150562 511634
rect 150646 511398 150882 511634
rect 150326 475718 150562 475954
rect 150646 475718 150882 475954
rect 150326 475398 150562 475634
rect 150646 475398 150882 475634
rect 150326 439718 150562 439954
rect 150646 439718 150882 439954
rect 150326 439398 150562 439634
rect 150646 439398 150882 439634
rect 150326 403718 150562 403954
rect 150646 403718 150882 403954
rect 150326 403398 150562 403634
rect 150646 403398 150882 403634
rect 150326 367718 150562 367954
rect 150646 367718 150882 367954
rect 150326 367398 150562 367634
rect 150646 367398 150882 367634
rect 150326 331718 150562 331954
rect 150646 331718 150882 331954
rect 150326 331398 150562 331634
rect 150646 331398 150882 331634
rect 150326 295718 150562 295954
rect 150646 295718 150882 295954
rect 150326 295398 150562 295634
rect 150646 295398 150882 295634
rect 150326 259718 150562 259954
rect 150646 259718 150882 259954
rect 150326 259398 150562 259634
rect 150646 259398 150882 259634
rect 154826 706522 155062 706758
rect 155146 706522 155382 706758
rect 154826 706202 155062 706438
rect 155146 706202 155382 706438
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 154826 660218 155062 660454
rect 155146 660218 155382 660454
rect 154826 659898 155062 660134
rect 155146 659898 155382 660134
rect 154826 624218 155062 624454
rect 155146 624218 155382 624454
rect 154826 623898 155062 624134
rect 155146 623898 155382 624134
rect 154826 588218 155062 588454
rect 155146 588218 155382 588454
rect 154826 587898 155062 588134
rect 155146 587898 155382 588134
rect 154826 552218 155062 552454
rect 155146 552218 155382 552454
rect 154826 551898 155062 552134
rect 155146 551898 155382 552134
rect 154826 516218 155062 516454
rect 155146 516218 155382 516454
rect 154826 515898 155062 516134
rect 155146 515898 155382 516134
rect 154826 480218 155062 480454
rect 155146 480218 155382 480454
rect 154826 479898 155062 480134
rect 155146 479898 155382 480134
rect 154826 444218 155062 444454
rect 155146 444218 155382 444454
rect 154826 443898 155062 444134
rect 155146 443898 155382 444134
rect 154826 408218 155062 408454
rect 155146 408218 155382 408454
rect 154826 407898 155062 408134
rect 155146 407898 155382 408134
rect 154826 372218 155062 372454
rect 155146 372218 155382 372454
rect 154826 371898 155062 372134
rect 155146 371898 155382 372134
rect 154826 336218 155062 336454
rect 155146 336218 155382 336454
rect 154826 335898 155062 336134
rect 155146 335898 155382 336134
rect 154826 300218 155062 300454
rect 155146 300218 155382 300454
rect 154826 299898 155062 300134
rect 155146 299898 155382 300134
rect 154826 264218 155062 264454
rect 155146 264218 155382 264454
rect 154826 263898 155062 264134
rect 155146 263898 155382 264134
rect 159326 707482 159562 707718
rect 159646 707482 159882 707718
rect 159326 707162 159562 707398
rect 159646 707162 159882 707398
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 159326 664718 159562 664954
rect 159646 664718 159882 664954
rect 159326 664398 159562 664634
rect 159646 664398 159882 664634
rect 159326 628718 159562 628954
rect 159646 628718 159882 628954
rect 159326 628398 159562 628634
rect 159646 628398 159882 628634
rect 159326 592718 159562 592954
rect 159646 592718 159882 592954
rect 159326 592398 159562 592634
rect 159646 592398 159882 592634
rect 159326 556718 159562 556954
rect 159646 556718 159882 556954
rect 159326 556398 159562 556634
rect 159646 556398 159882 556634
rect 159326 520718 159562 520954
rect 159646 520718 159882 520954
rect 159326 520398 159562 520634
rect 159646 520398 159882 520634
rect 159326 484718 159562 484954
rect 159646 484718 159882 484954
rect 159326 484398 159562 484634
rect 159646 484398 159882 484634
rect 159326 448718 159562 448954
rect 159646 448718 159882 448954
rect 159326 448398 159562 448634
rect 159646 448398 159882 448634
rect 159326 412718 159562 412954
rect 159646 412718 159882 412954
rect 159326 412398 159562 412634
rect 159646 412398 159882 412634
rect 159326 376718 159562 376954
rect 159646 376718 159882 376954
rect 159326 376398 159562 376634
rect 159646 376398 159882 376634
rect 159326 340718 159562 340954
rect 159646 340718 159882 340954
rect 159326 340398 159562 340634
rect 159646 340398 159882 340634
rect 159326 304718 159562 304954
rect 159646 304718 159882 304954
rect 159326 304398 159562 304634
rect 159646 304398 159882 304634
rect 159326 268718 159562 268954
rect 159646 268718 159882 268954
rect 159326 268398 159562 268634
rect 159646 268398 159882 268634
rect 163826 708442 164062 708678
rect 164146 708442 164382 708678
rect 163826 708122 164062 708358
rect 164146 708122 164382 708358
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 168326 709402 168562 709638
rect 168646 709402 168882 709638
rect 168326 709082 168562 709318
rect 168646 709082 168882 709318
rect 168326 673718 168562 673954
rect 168646 673718 168882 673954
rect 168326 673398 168562 673634
rect 168646 673398 168882 673634
rect 168326 637718 168562 637954
rect 168646 637718 168882 637954
rect 168326 637398 168562 637634
rect 168646 637398 168882 637634
rect 168326 601718 168562 601954
rect 168646 601718 168882 601954
rect 168326 601398 168562 601634
rect 168646 601398 168882 601634
rect 168326 565718 168562 565954
rect 168646 565718 168882 565954
rect 168326 565398 168562 565634
rect 168646 565398 168882 565634
rect 168326 529718 168562 529954
rect 168646 529718 168882 529954
rect 168326 529398 168562 529634
rect 168646 529398 168882 529634
rect 168326 493718 168562 493954
rect 168646 493718 168882 493954
rect 168326 493398 168562 493634
rect 168646 493398 168882 493634
rect 168326 457718 168562 457954
rect 168646 457718 168882 457954
rect 168326 457398 168562 457634
rect 168646 457398 168882 457634
rect 168326 421718 168562 421954
rect 168646 421718 168882 421954
rect 168326 421398 168562 421634
rect 168646 421398 168882 421634
rect 168326 385718 168562 385954
rect 168646 385718 168882 385954
rect 168326 385398 168562 385634
rect 168646 385398 168882 385634
rect 168326 349718 168562 349954
rect 168646 349718 168882 349954
rect 168326 349398 168562 349634
rect 168646 349398 168882 349634
rect 168326 313718 168562 313954
rect 168646 313718 168882 313954
rect 168326 313398 168562 313634
rect 168646 313398 168882 313634
rect 168326 277718 168562 277954
rect 168646 277718 168882 277954
rect 168326 277398 168562 277634
rect 168646 277398 168882 277634
rect 172826 710362 173062 710598
rect 173146 710362 173382 710598
rect 172826 710042 173062 710278
rect 173146 710042 173382 710278
rect 172826 678218 173062 678454
rect 173146 678218 173382 678454
rect 172826 677898 173062 678134
rect 173146 677898 173382 678134
rect 172826 642218 173062 642454
rect 173146 642218 173382 642454
rect 172826 641898 173062 642134
rect 173146 641898 173382 642134
rect 172826 606218 173062 606454
rect 173146 606218 173382 606454
rect 172826 605898 173062 606134
rect 173146 605898 173382 606134
rect 172826 570218 173062 570454
rect 173146 570218 173382 570454
rect 172826 569898 173062 570134
rect 173146 569898 173382 570134
rect 172826 534218 173062 534454
rect 173146 534218 173382 534454
rect 172826 533898 173062 534134
rect 173146 533898 173382 534134
rect 172826 498218 173062 498454
rect 173146 498218 173382 498454
rect 172826 497898 173062 498134
rect 173146 497898 173382 498134
rect 172826 462218 173062 462454
rect 173146 462218 173382 462454
rect 172826 461898 173062 462134
rect 173146 461898 173382 462134
rect 172826 426218 173062 426454
rect 173146 426218 173382 426454
rect 172826 425898 173062 426134
rect 173146 425898 173382 426134
rect 172826 390218 173062 390454
rect 173146 390218 173382 390454
rect 172826 389898 173062 390134
rect 173146 389898 173382 390134
rect 172826 354218 173062 354454
rect 173146 354218 173382 354454
rect 172826 353898 173062 354134
rect 173146 353898 173382 354134
rect 172826 318218 173062 318454
rect 173146 318218 173382 318454
rect 172826 317898 173062 318134
rect 173146 317898 173382 318134
rect 172826 282218 173062 282454
rect 173146 282218 173382 282454
rect 172826 281898 173062 282134
rect 173146 281898 173382 282134
rect 177326 711322 177562 711558
rect 177646 711322 177882 711558
rect 177326 711002 177562 711238
rect 177646 711002 177882 711238
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 177326 646718 177562 646954
rect 177646 646718 177882 646954
rect 177326 646398 177562 646634
rect 177646 646398 177882 646634
rect 177326 610718 177562 610954
rect 177646 610718 177882 610954
rect 177326 610398 177562 610634
rect 177646 610398 177882 610634
rect 177326 574718 177562 574954
rect 177646 574718 177882 574954
rect 177326 574398 177562 574634
rect 177646 574398 177882 574634
rect 177326 538718 177562 538954
rect 177646 538718 177882 538954
rect 177326 538398 177562 538634
rect 177646 538398 177882 538634
rect 177326 502718 177562 502954
rect 177646 502718 177882 502954
rect 177326 502398 177562 502634
rect 177646 502398 177882 502634
rect 177326 466718 177562 466954
rect 177646 466718 177882 466954
rect 177326 466398 177562 466634
rect 177646 466398 177882 466634
rect 177326 430718 177562 430954
rect 177646 430718 177882 430954
rect 177326 430398 177562 430634
rect 177646 430398 177882 430634
rect 177326 394718 177562 394954
rect 177646 394718 177882 394954
rect 177326 394398 177562 394634
rect 177646 394398 177882 394634
rect 177326 358718 177562 358954
rect 177646 358718 177882 358954
rect 177326 358398 177562 358634
rect 177646 358398 177882 358634
rect 177326 322718 177562 322954
rect 177646 322718 177882 322954
rect 177326 322398 177562 322634
rect 177646 322398 177882 322634
rect 177326 286718 177562 286954
rect 177646 286718 177882 286954
rect 177326 286398 177562 286634
rect 177646 286398 177882 286634
rect 177326 250718 177562 250954
rect 177646 250718 177882 250954
rect 177326 250398 177562 250634
rect 177646 250398 177882 250634
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 186326 705562 186562 705798
rect 186646 705562 186882 705798
rect 186326 705242 186562 705478
rect 186646 705242 186882 705478
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 186326 655718 186562 655954
rect 186646 655718 186882 655954
rect 186326 655398 186562 655634
rect 186646 655398 186882 655634
rect 186326 619718 186562 619954
rect 186646 619718 186882 619954
rect 186326 619398 186562 619634
rect 186646 619398 186882 619634
rect 186326 583718 186562 583954
rect 186646 583718 186882 583954
rect 186326 583398 186562 583634
rect 186646 583398 186882 583634
rect 186326 547718 186562 547954
rect 186646 547718 186882 547954
rect 186326 547398 186562 547634
rect 186646 547398 186882 547634
rect 186326 511718 186562 511954
rect 186646 511718 186882 511954
rect 186326 511398 186562 511634
rect 186646 511398 186882 511634
rect 186326 475718 186562 475954
rect 186646 475718 186882 475954
rect 186326 475398 186562 475634
rect 186646 475398 186882 475634
rect 186326 439718 186562 439954
rect 186646 439718 186882 439954
rect 186326 439398 186562 439634
rect 186646 439398 186882 439634
rect 186326 403718 186562 403954
rect 186646 403718 186882 403954
rect 186326 403398 186562 403634
rect 186646 403398 186882 403634
rect 186326 367718 186562 367954
rect 186646 367718 186882 367954
rect 186326 367398 186562 367634
rect 186646 367398 186882 367634
rect 186326 331718 186562 331954
rect 186646 331718 186882 331954
rect 186326 331398 186562 331634
rect 186646 331398 186882 331634
rect 186326 295718 186562 295954
rect 186646 295718 186882 295954
rect 186326 295398 186562 295634
rect 186646 295398 186882 295634
rect 186326 259718 186562 259954
rect 186646 259718 186882 259954
rect 186326 259398 186562 259634
rect 186646 259398 186882 259634
rect 190826 706522 191062 706758
rect 191146 706522 191382 706758
rect 190826 706202 191062 706438
rect 191146 706202 191382 706438
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 190826 660218 191062 660454
rect 191146 660218 191382 660454
rect 190826 659898 191062 660134
rect 191146 659898 191382 660134
rect 190826 624218 191062 624454
rect 191146 624218 191382 624454
rect 190826 623898 191062 624134
rect 191146 623898 191382 624134
rect 190826 588218 191062 588454
rect 191146 588218 191382 588454
rect 190826 587898 191062 588134
rect 191146 587898 191382 588134
rect 190826 552218 191062 552454
rect 191146 552218 191382 552454
rect 190826 551898 191062 552134
rect 191146 551898 191382 552134
rect 190826 516218 191062 516454
rect 191146 516218 191382 516454
rect 190826 515898 191062 516134
rect 191146 515898 191382 516134
rect 190826 480218 191062 480454
rect 191146 480218 191382 480454
rect 190826 479898 191062 480134
rect 191146 479898 191382 480134
rect 190826 444218 191062 444454
rect 191146 444218 191382 444454
rect 190826 443898 191062 444134
rect 191146 443898 191382 444134
rect 190826 408218 191062 408454
rect 191146 408218 191382 408454
rect 190826 407898 191062 408134
rect 191146 407898 191382 408134
rect 190826 372218 191062 372454
rect 191146 372218 191382 372454
rect 190826 371898 191062 372134
rect 191146 371898 191382 372134
rect 190826 336218 191062 336454
rect 191146 336218 191382 336454
rect 190826 335898 191062 336134
rect 191146 335898 191382 336134
rect 190826 300218 191062 300454
rect 191146 300218 191382 300454
rect 190826 299898 191062 300134
rect 191146 299898 191382 300134
rect 190826 264218 191062 264454
rect 191146 264218 191382 264454
rect 190826 263898 191062 264134
rect 191146 263898 191382 264134
rect 195326 707482 195562 707718
rect 195646 707482 195882 707718
rect 195326 707162 195562 707398
rect 195646 707162 195882 707398
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 195326 664718 195562 664954
rect 195646 664718 195882 664954
rect 195326 664398 195562 664634
rect 195646 664398 195882 664634
rect 195326 628718 195562 628954
rect 195646 628718 195882 628954
rect 195326 628398 195562 628634
rect 195646 628398 195882 628634
rect 195326 592718 195562 592954
rect 195646 592718 195882 592954
rect 195326 592398 195562 592634
rect 195646 592398 195882 592634
rect 195326 556718 195562 556954
rect 195646 556718 195882 556954
rect 195326 556398 195562 556634
rect 195646 556398 195882 556634
rect 195326 520718 195562 520954
rect 195646 520718 195882 520954
rect 195326 520398 195562 520634
rect 195646 520398 195882 520634
rect 195326 484718 195562 484954
rect 195646 484718 195882 484954
rect 195326 484398 195562 484634
rect 195646 484398 195882 484634
rect 195326 448718 195562 448954
rect 195646 448718 195882 448954
rect 195326 448398 195562 448634
rect 195646 448398 195882 448634
rect 195326 412718 195562 412954
rect 195646 412718 195882 412954
rect 195326 412398 195562 412634
rect 195646 412398 195882 412634
rect 195326 376718 195562 376954
rect 195646 376718 195882 376954
rect 195326 376398 195562 376634
rect 195646 376398 195882 376634
rect 195326 340718 195562 340954
rect 195646 340718 195882 340954
rect 195326 340398 195562 340634
rect 195646 340398 195882 340634
rect 195326 304718 195562 304954
rect 195646 304718 195882 304954
rect 195326 304398 195562 304634
rect 195646 304398 195882 304634
rect 195326 268718 195562 268954
rect 195646 268718 195882 268954
rect 195326 268398 195562 268634
rect 195646 268398 195882 268634
rect 199826 708442 200062 708678
rect 200146 708442 200382 708678
rect 199826 708122 200062 708358
rect 200146 708122 200382 708358
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 204326 709402 204562 709638
rect 204646 709402 204882 709638
rect 204326 709082 204562 709318
rect 204646 709082 204882 709318
rect 204326 673718 204562 673954
rect 204646 673718 204882 673954
rect 204326 673398 204562 673634
rect 204646 673398 204882 673634
rect 204326 637718 204562 637954
rect 204646 637718 204882 637954
rect 204326 637398 204562 637634
rect 204646 637398 204882 637634
rect 204326 601718 204562 601954
rect 204646 601718 204882 601954
rect 204326 601398 204562 601634
rect 204646 601398 204882 601634
rect 204326 565718 204562 565954
rect 204646 565718 204882 565954
rect 204326 565398 204562 565634
rect 204646 565398 204882 565634
rect 204326 529718 204562 529954
rect 204646 529718 204882 529954
rect 204326 529398 204562 529634
rect 204646 529398 204882 529634
rect 204326 493718 204562 493954
rect 204646 493718 204882 493954
rect 204326 493398 204562 493634
rect 204646 493398 204882 493634
rect 204326 457718 204562 457954
rect 204646 457718 204882 457954
rect 204326 457398 204562 457634
rect 204646 457398 204882 457634
rect 204326 421718 204562 421954
rect 204646 421718 204882 421954
rect 204326 421398 204562 421634
rect 204646 421398 204882 421634
rect 204326 385718 204562 385954
rect 204646 385718 204882 385954
rect 204326 385398 204562 385634
rect 204646 385398 204882 385634
rect 204326 349718 204562 349954
rect 204646 349718 204882 349954
rect 204326 349398 204562 349634
rect 204646 349398 204882 349634
rect 204326 313718 204562 313954
rect 204646 313718 204882 313954
rect 204326 313398 204562 313634
rect 204646 313398 204882 313634
rect 204326 277718 204562 277954
rect 204646 277718 204882 277954
rect 204326 277398 204562 277634
rect 204646 277398 204882 277634
rect 208826 710362 209062 710598
rect 209146 710362 209382 710598
rect 208826 710042 209062 710278
rect 209146 710042 209382 710278
rect 208826 678218 209062 678454
rect 209146 678218 209382 678454
rect 208826 677898 209062 678134
rect 209146 677898 209382 678134
rect 208826 642218 209062 642454
rect 209146 642218 209382 642454
rect 208826 641898 209062 642134
rect 209146 641898 209382 642134
rect 208826 606218 209062 606454
rect 209146 606218 209382 606454
rect 208826 605898 209062 606134
rect 209146 605898 209382 606134
rect 208826 570218 209062 570454
rect 209146 570218 209382 570454
rect 208826 569898 209062 570134
rect 209146 569898 209382 570134
rect 208826 534218 209062 534454
rect 209146 534218 209382 534454
rect 208826 533898 209062 534134
rect 209146 533898 209382 534134
rect 208826 498218 209062 498454
rect 209146 498218 209382 498454
rect 208826 497898 209062 498134
rect 209146 497898 209382 498134
rect 208826 462218 209062 462454
rect 209146 462218 209382 462454
rect 208826 461898 209062 462134
rect 209146 461898 209382 462134
rect 208826 426218 209062 426454
rect 209146 426218 209382 426454
rect 208826 425898 209062 426134
rect 209146 425898 209382 426134
rect 208826 390218 209062 390454
rect 209146 390218 209382 390454
rect 208826 389898 209062 390134
rect 209146 389898 209382 390134
rect 208826 354218 209062 354454
rect 209146 354218 209382 354454
rect 208826 353898 209062 354134
rect 209146 353898 209382 354134
rect 208826 318218 209062 318454
rect 209146 318218 209382 318454
rect 208826 317898 209062 318134
rect 209146 317898 209382 318134
rect 208826 282218 209062 282454
rect 209146 282218 209382 282454
rect 208826 281898 209062 282134
rect 209146 281898 209382 282134
rect 213326 711322 213562 711558
rect 213646 711322 213882 711558
rect 213326 711002 213562 711238
rect 213646 711002 213882 711238
rect 213326 682718 213562 682954
rect 213646 682718 213882 682954
rect 213326 682398 213562 682634
rect 213646 682398 213882 682634
rect 213326 646718 213562 646954
rect 213646 646718 213882 646954
rect 213326 646398 213562 646634
rect 213646 646398 213882 646634
rect 213326 610718 213562 610954
rect 213646 610718 213882 610954
rect 213326 610398 213562 610634
rect 213646 610398 213882 610634
rect 213326 574718 213562 574954
rect 213646 574718 213882 574954
rect 213326 574398 213562 574634
rect 213646 574398 213882 574634
rect 213326 538718 213562 538954
rect 213646 538718 213882 538954
rect 213326 538398 213562 538634
rect 213646 538398 213882 538634
rect 213326 502718 213562 502954
rect 213646 502718 213882 502954
rect 213326 502398 213562 502634
rect 213646 502398 213882 502634
rect 213326 466718 213562 466954
rect 213646 466718 213882 466954
rect 213326 466398 213562 466634
rect 213646 466398 213882 466634
rect 213326 430718 213562 430954
rect 213646 430718 213882 430954
rect 213326 430398 213562 430634
rect 213646 430398 213882 430634
rect 213326 394718 213562 394954
rect 213646 394718 213882 394954
rect 213326 394398 213562 394634
rect 213646 394398 213882 394634
rect 213326 358718 213562 358954
rect 213646 358718 213882 358954
rect 213326 358398 213562 358634
rect 213646 358398 213882 358634
rect 213326 322718 213562 322954
rect 213646 322718 213882 322954
rect 213326 322398 213562 322634
rect 213646 322398 213882 322634
rect 213326 286718 213562 286954
rect 213646 286718 213882 286954
rect 213326 286398 213562 286634
rect 213646 286398 213882 286634
rect 213326 250718 213562 250954
rect 213646 250718 213882 250954
rect 213326 250398 213562 250634
rect 213646 250398 213882 250634
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 222326 705562 222562 705798
rect 222646 705562 222882 705798
rect 222326 705242 222562 705478
rect 222646 705242 222882 705478
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 222326 655718 222562 655954
rect 222646 655718 222882 655954
rect 222326 655398 222562 655634
rect 222646 655398 222882 655634
rect 222326 619718 222562 619954
rect 222646 619718 222882 619954
rect 222326 619398 222562 619634
rect 222646 619398 222882 619634
rect 222326 583718 222562 583954
rect 222646 583718 222882 583954
rect 222326 583398 222562 583634
rect 222646 583398 222882 583634
rect 222326 547718 222562 547954
rect 222646 547718 222882 547954
rect 222326 547398 222562 547634
rect 222646 547398 222882 547634
rect 222326 511718 222562 511954
rect 222646 511718 222882 511954
rect 222326 511398 222562 511634
rect 222646 511398 222882 511634
rect 222326 475718 222562 475954
rect 222646 475718 222882 475954
rect 222326 475398 222562 475634
rect 222646 475398 222882 475634
rect 222326 439718 222562 439954
rect 222646 439718 222882 439954
rect 222326 439398 222562 439634
rect 222646 439398 222882 439634
rect 222326 403718 222562 403954
rect 222646 403718 222882 403954
rect 222326 403398 222562 403634
rect 222646 403398 222882 403634
rect 222326 367718 222562 367954
rect 222646 367718 222882 367954
rect 222326 367398 222562 367634
rect 222646 367398 222882 367634
rect 222326 331718 222562 331954
rect 222646 331718 222882 331954
rect 222326 331398 222562 331634
rect 222646 331398 222882 331634
rect 222326 295718 222562 295954
rect 222646 295718 222882 295954
rect 222326 295398 222562 295634
rect 222646 295398 222882 295634
rect 222326 259718 222562 259954
rect 222646 259718 222882 259954
rect 222326 259398 222562 259634
rect 222646 259398 222882 259634
rect 226826 706522 227062 706758
rect 227146 706522 227382 706758
rect 226826 706202 227062 706438
rect 227146 706202 227382 706438
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 226826 660218 227062 660454
rect 227146 660218 227382 660454
rect 226826 659898 227062 660134
rect 227146 659898 227382 660134
rect 226826 624218 227062 624454
rect 227146 624218 227382 624454
rect 226826 623898 227062 624134
rect 227146 623898 227382 624134
rect 226826 588218 227062 588454
rect 227146 588218 227382 588454
rect 226826 587898 227062 588134
rect 227146 587898 227382 588134
rect 226826 552218 227062 552454
rect 227146 552218 227382 552454
rect 226826 551898 227062 552134
rect 227146 551898 227382 552134
rect 226826 516218 227062 516454
rect 227146 516218 227382 516454
rect 226826 515898 227062 516134
rect 227146 515898 227382 516134
rect 226826 480218 227062 480454
rect 227146 480218 227382 480454
rect 226826 479898 227062 480134
rect 227146 479898 227382 480134
rect 226826 444218 227062 444454
rect 227146 444218 227382 444454
rect 226826 443898 227062 444134
rect 227146 443898 227382 444134
rect 226826 408218 227062 408454
rect 227146 408218 227382 408454
rect 226826 407898 227062 408134
rect 227146 407898 227382 408134
rect 226826 372218 227062 372454
rect 227146 372218 227382 372454
rect 226826 371898 227062 372134
rect 227146 371898 227382 372134
rect 226826 336218 227062 336454
rect 227146 336218 227382 336454
rect 226826 335898 227062 336134
rect 227146 335898 227382 336134
rect 226826 300218 227062 300454
rect 227146 300218 227382 300454
rect 226826 299898 227062 300134
rect 227146 299898 227382 300134
rect 226826 264218 227062 264454
rect 227146 264218 227382 264454
rect 226826 263898 227062 264134
rect 227146 263898 227382 264134
rect 231326 707482 231562 707718
rect 231646 707482 231882 707718
rect 231326 707162 231562 707398
rect 231646 707162 231882 707398
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 231326 664718 231562 664954
rect 231646 664718 231882 664954
rect 231326 664398 231562 664634
rect 231646 664398 231882 664634
rect 231326 628718 231562 628954
rect 231646 628718 231882 628954
rect 231326 628398 231562 628634
rect 231646 628398 231882 628634
rect 231326 592718 231562 592954
rect 231646 592718 231882 592954
rect 231326 592398 231562 592634
rect 231646 592398 231882 592634
rect 231326 556718 231562 556954
rect 231646 556718 231882 556954
rect 231326 556398 231562 556634
rect 231646 556398 231882 556634
rect 231326 520718 231562 520954
rect 231646 520718 231882 520954
rect 231326 520398 231562 520634
rect 231646 520398 231882 520634
rect 231326 484718 231562 484954
rect 231646 484718 231882 484954
rect 231326 484398 231562 484634
rect 231646 484398 231882 484634
rect 231326 448718 231562 448954
rect 231646 448718 231882 448954
rect 231326 448398 231562 448634
rect 231646 448398 231882 448634
rect 231326 412718 231562 412954
rect 231646 412718 231882 412954
rect 231326 412398 231562 412634
rect 231646 412398 231882 412634
rect 231326 376718 231562 376954
rect 231646 376718 231882 376954
rect 231326 376398 231562 376634
rect 231646 376398 231882 376634
rect 231326 340718 231562 340954
rect 231646 340718 231882 340954
rect 231326 340398 231562 340634
rect 231646 340398 231882 340634
rect 231326 304718 231562 304954
rect 231646 304718 231882 304954
rect 231326 304398 231562 304634
rect 231646 304398 231882 304634
rect 231326 268718 231562 268954
rect 231646 268718 231882 268954
rect 231326 268398 231562 268634
rect 231646 268398 231882 268634
rect 235826 708442 236062 708678
rect 236146 708442 236382 708678
rect 235826 708122 236062 708358
rect 236146 708122 236382 708358
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 240326 709402 240562 709638
rect 240646 709402 240882 709638
rect 240326 709082 240562 709318
rect 240646 709082 240882 709318
rect 240326 673718 240562 673954
rect 240646 673718 240882 673954
rect 240326 673398 240562 673634
rect 240646 673398 240882 673634
rect 240326 637718 240562 637954
rect 240646 637718 240882 637954
rect 240326 637398 240562 637634
rect 240646 637398 240882 637634
rect 240326 601718 240562 601954
rect 240646 601718 240882 601954
rect 240326 601398 240562 601634
rect 240646 601398 240882 601634
rect 240326 565718 240562 565954
rect 240646 565718 240882 565954
rect 240326 565398 240562 565634
rect 240646 565398 240882 565634
rect 240326 529718 240562 529954
rect 240646 529718 240882 529954
rect 240326 529398 240562 529634
rect 240646 529398 240882 529634
rect 240326 493718 240562 493954
rect 240646 493718 240882 493954
rect 240326 493398 240562 493634
rect 240646 493398 240882 493634
rect 240326 457718 240562 457954
rect 240646 457718 240882 457954
rect 240326 457398 240562 457634
rect 240646 457398 240882 457634
rect 240326 421718 240562 421954
rect 240646 421718 240882 421954
rect 240326 421398 240562 421634
rect 240646 421398 240882 421634
rect 240326 385718 240562 385954
rect 240646 385718 240882 385954
rect 240326 385398 240562 385634
rect 240646 385398 240882 385634
rect 240326 349718 240562 349954
rect 240646 349718 240882 349954
rect 240326 349398 240562 349634
rect 240646 349398 240882 349634
rect 240326 313718 240562 313954
rect 240646 313718 240882 313954
rect 240326 313398 240562 313634
rect 240646 313398 240882 313634
rect 240326 277718 240562 277954
rect 240646 277718 240882 277954
rect 240326 277398 240562 277634
rect 240646 277398 240882 277634
rect 244826 710362 245062 710598
rect 245146 710362 245382 710598
rect 244826 710042 245062 710278
rect 245146 710042 245382 710278
rect 244826 678218 245062 678454
rect 245146 678218 245382 678454
rect 244826 677898 245062 678134
rect 245146 677898 245382 678134
rect 244826 642218 245062 642454
rect 245146 642218 245382 642454
rect 244826 641898 245062 642134
rect 245146 641898 245382 642134
rect 244826 606218 245062 606454
rect 245146 606218 245382 606454
rect 244826 605898 245062 606134
rect 245146 605898 245382 606134
rect 244826 570218 245062 570454
rect 245146 570218 245382 570454
rect 244826 569898 245062 570134
rect 245146 569898 245382 570134
rect 244826 534218 245062 534454
rect 245146 534218 245382 534454
rect 244826 533898 245062 534134
rect 245146 533898 245382 534134
rect 244826 498218 245062 498454
rect 245146 498218 245382 498454
rect 244826 497898 245062 498134
rect 245146 497898 245382 498134
rect 244826 462218 245062 462454
rect 245146 462218 245382 462454
rect 244826 461898 245062 462134
rect 245146 461898 245382 462134
rect 244826 426218 245062 426454
rect 245146 426218 245382 426454
rect 244826 425898 245062 426134
rect 245146 425898 245382 426134
rect 244826 390218 245062 390454
rect 245146 390218 245382 390454
rect 244826 389898 245062 390134
rect 245146 389898 245382 390134
rect 244826 354218 245062 354454
rect 245146 354218 245382 354454
rect 244826 353898 245062 354134
rect 245146 353898 245382 354134
rect 244826 318218 245062 318454
rect 245146 318218 245382 318454
rect 244826 317898 245062 318134
rect 245146 317898 245382 318134
rect 244826 282218 245062 282454
rect 245146 282218 245382 282454
rect 244826 281898 245062 282134
rect 245146 281898 245382 282134
rect 249326 711322 249562 711558
rect 249646 711322 249882 711558
rect 249326 711002 249562 711238
rect 249646 711002 249882 711238
rect 249326 682718 249562 682954
rect 249646 682718 249882 682954
rect 249326 682398 249562 682634
rect 249646 682398 249882 682634
rect 249326 646718 249562 646954
rect 249646 646718 249882 646954
rect 249326 646398 249562 646634
rect 249646 646398 249882 646634
rect 249326 610718 249562 610954
rect 249646 610718 249882 610954
rect 249326 610398 249562 610634
rect 249646 610398 249882 610634
rect 249326 574718 249562 574954
rect 249646 574718 249882 574954
rect 249326 574398 249562 574634
rect 249646 574398 249882 574634
rect 249326 538718 249562 538954
rect 249646 538718 249882 538954
rect 249326 538398 249562 538634
rect 249646 538398 249882 538634
rect 249326 502718 249562 502954
rect 249646 502718 249882 502954
rect 249326 502398 249562 502634
rect 249646 502398 249882 502634
rect 249326 466718 249562 466954
rect 249646 466718 249882 466954
rect 249326 466398 249562 466634
rect 249646 466398 249882 466634
rect 249326 430718 249562 430954
rect 249646 430718 249882 430954
rect 249326 430398 249562 430634
rect 249646 430398 249882 430634
rect 249326 394718 249562 394954
rect 249646 394718 249882 394954
rect 249326 394398 249562 394634
rect 249646 394398 249882 394634
rect 249326 358718 249562 358954
rect 249646 358718 249882 358954
rect 249326 358398 249562 358634
rect 249646 358398 249882 358634
rect 249326 322718 249562 322954
rect 249646 322718 249882 322954
rect 249326 322398 249562 322634
rect 249646 322398 249882 322634
rect 249326 286718 249562 286954
rect 249646 286718 249882 286954
rect 249326 286398 249562 286634
rect 249646 286398 249882 286634
rect 249326 250718 249562 250954
rect 249646 250718 249882 250954
rect 249326 250398 249562 250634
rect 249646 250398 249882 250634
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 258326 705562 258562 705798
rect 258646 705562 258882 705798
rect 258326 705242 258562 705478
rect 258646 705242 258882 705478
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 258326 655718 258562 655954
rect 258646 655718 258882 655954
rect 258326 655398 258562 655634
rect 258646 655398 258882 655634
rect 258326 619718 258562 619954
rect 258646 619718 258882 619954
rect 258326 619398 258562 619634
rect 258646 619398 258882 619634
rect 258326 583718 258562 583954
rect 258646 583718 258882 583954
rect 258326 583398 258562 583634
rect 258646 583398 258882 583634
rect 258326 547718 258562 547954
rect 258646 547718 258882 547954
rect 258326 547398 258562 547634
rect 258646 547398 258882 547634
rect 258326 511718 258562 511954
rect 258646 511718 258882 511954
rect 258326 511398 258562 511634
rect 258646 511398 258882 511634
rect 258326 475718 258562 475954
rect 258646 475718 258882 475954
rect 258326 475398 258562 475634
rect 258646 475398 258882 475634
rect 258326 439718 258562 439954
rect 258646 439718 258882 439954
rect 258326 439398 258562 439634
rect 258646 439398 258882 439634
rect 258326 403718 258562 403954
rect 258646 403718 258882 403954
rect 258326 403398 258562 403634
rect 258646 403398 258882 403634
rect 258326 367718 258562 367954
rect 258646 367718 258882 367954
rect 258326 367398 258562 367634
rect 258646 367398 258882 367634
rect 258326 331718 258562 331954
rect 258646 331718 258882 331954
rect 258326 331398 258562 331634
rect 258646 331398 258882 331634
rect 258326 295718 258562 295954
rect 258646 295718 258882 295954
rect 258326 295398 258562 295634
rect 258646 295398 258882 295634
rect 258326 259718 258562 259954
rect 258646 259718 258882 259954
rect 258326 259398 258562 259634
rect 258646 259398 258882 259634
rect 262826 706522 263062 706758
rect 263146 706522 263382 706758
rect 262826 706202 263062 706438
rect 263146 706202 263382 706438
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 262826 660218 263062 660454
rect 263146 660218 263382 660454
rect 262826 659898 263062 660134
rect 263146 659898 263382 660134
rect 262826 624218 263062 624454
rect 263146 624218 263382 624454
rect 262826 623898 263062 624134
rect 263146 623898 263382 624134
rect 262826 588218 263062 588454
rect 263146 588218 263382 588454
rect 262826 587898 263062 588134
rect 263146 587898 263382 588134
rect 262826 552218 263062 552454
rect 263146 552218 263382 552454
rect 262826 551898 263062 552134
rect 263146 551898 263382 552134
rect 262826 516218 263062 516454
rect 263146 516218 263382 516454
rect 262826 515898 263062 516134
rect 263146 515898 263382 516134
rect 262826 480218 263062 480454
rect 263146 480218 263382 480454
rect 262826 479898 263062 480134
rect 263146 479898 263382 480134
rect 262826 444218 263062 444454
rect 263146 444218 263382 444454
rect 262826 443898 263062 444134
rect 263146 443898 263382 444134
rect 262826 408218 263062 408454
rect 263146 408218 263382 408454
rect 262826 407898 263062 408134
rect 263146 407898 263382 408134
rect 262826 372218 263062 372454
rect 263146 372218 263382 372454
rect 262826 371898 263062 372134
rect 263146 371898 263382 372134
rect 262826 336218 263062 336454
rect 263146 336218 263382 336454
rect 262826 335898 263062 336134
rect 263146 335898 263382 336134
rect 262826 300218 263062 300454
rect 263146 300218 263382 300454
rect 262826 299898 263062 300134
rect 263146 299898 263382 300134
rect 262826 264218 263062 264454
rect 263146 264218 263382 264454
rect 262826 263898 263062 264134
rect 263146 263898 263382 264134
rect 267326 707482 267562 707718
rect 267646 707482 267882 707718
rect 267326 707162 267562 707398
rect 267646 707162 267882 707398
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 267326 664718 267562 664954
rect 267646 664718 267882 664954
rect 267326 664398 267562 664634
rect 267646 664398 267882 664634
rect 267326 628718 267562 628954
rect 267646 628718 267882 628954
rect 267326 628398 267562 628634
rect 267646 628398 267882 628634
rect 267326 592718 267562 592954
rect 267646 592718 267882 592954
rect 267326 592398 267562 592634
rect 267646 592398 267882 592634
rect 267326 556718 267562 556954
rect 267646 556718 267882 556954
rect 267326 556398 267562 556634
rect 267646 556398 267882 556634
rect 267326 520718 267562 520954
rect 267646 520718 267882 520954
rect 267326 520398 267562 520634
rect 267646 520398 267882 520634
rect 267326 484718 267562 484954
rect 267646 484718 267882 484954
rect 267326 484398 267562 484634
rect 267646 484398 267882 484634
rect 267326 448718 267562 448954
rect 267646 448718 267882 448954
rect 267326 448398 267562 448634
rect 267646 448398 267882 448634
rect 267326 412718 267562 412954
rect 267646 412718 267882 412954
rect 267326 412398 267562 412634
rect 267646 412398 267882 412634
rect 267326 376718 267562 376954
rect 267646 376718 267882 376954
rect 267326 376398 267562 376634
rect 267646 376398 267882 376634
rect 267326 340718 267562 340954
rect 267646 340718 267882 340954
rect 267326 340398 267562 340634
rect 267646 340398 267882 340634
rect 267326 304718 267562 304954
rect 267646 304718 267882 304954
rect 267326 304398 267562 304634
rect 267646 304398 267882 304634
rect 267326 268718 267562 268954
rect 267646 268718 267882 268954
rect 267326 268398 267562 268634
rect 267646 268398 267882 268634
rect 271826 708442 272062 708678
rect 272146 708442 272382 708678
rect 271826 708122 272062 708358
rect 272146 708122 272382 708358
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 276326 709402 276562 709638
rect 276646 709402 276882 709638
rect 276326 709082 276562 709318
rect 276646 709082 276882 709318
rect 276326 673718 276562 673954
rect 276646 673718 276882 673954
rect 276326 673398 276562 673634
rect 276646 673398 276882 673634
rect 276326 637718 276562 637954
rect 276646 637718 276882 637954
rect 276326 637398 276562 637634
rect 276646 637398 276882 637634
rect 276326 601718 276562 601954
rect 276646 601718 276882 601954
rect 276326 601398 276562 601634
rect 276646 601398 276882 601634
rect 276326 565718 276562 565954
rect 276646 565718 276882 565954
rect 276326 565398 276562 565634
rect 276646 565398 276882 565634
rect 276326 529718 276562 529954
rect 276646 529718 276882 529954
rect 276326 529398 276562 529634
rect 276646 529398 276882 529634
rect 276326 493718 276562 493954
rect 276646 493718 276882 493954
rect 276326 493398 276562 493634
rect 276646 493398 276882 493634
rect 276326 457718 276562 457954
rect 276646 457718 276882 457954
rect 276326 457398 276562 457634
rect 276646 457398 276882 457634
rect 276326 421718 276562 421954
rect 276646 421718 276882 421954
rect 276326 421398 276562 421634
rect 276646 421398 276882 421634
rect 276326 385718 276562 385954
rect 276646 385718 276882 385954
rect 276326 385398 276562 385634
rect 276646 385398 276882 385634
rect 276326 349718 276562 349954
rect 276646 349718 276882 349954
rect 276326 349398 276562 349634
rect 276646 349398 276882 349634
rect 276326 313718 276562 313954
rect 276646 313718 276882 313954
rect 276326 313398 276562 313634
rect 276646 313398 276882 313634
rect 276326 277718 276562 277954
rect 276646 277718 276882 277954
rect 276326 277398 276562 277634
rect 276646 277398 276882 277634
rect 280826 710362 281062 710598
rect 281146 710362 281382 710598
rect 280826 710042 281062 710278
rect 281146 710042 281382 710278
rect 280826 678218 281062 678454
rect 281146 678218 281382 678454
rect 280826 677898 281062 678134
rect 281146 677898 281382 678134
rect 280826 642218 281062 642454
rect 281146 642218 281382 642454
rect 280826 641898 281062 642134
rect 281146 641898 281382 642134
rect 280826 606218 281062 606454
rect 281146 606218 281382 606454
rect 280826 605898 281062 606134
rect 281146 605898 281382 606134
rect 280826 570218 281062 570454
rect 281146 570218 281382 570454
rect 280826 569898 281062 570134
rect 281146 569898 281382 570134
rect 280826 534218 281062 534454
rect 281146 534218 281382 534454
rect 280826 533898 281062 534134
rect 281146 533898 281382 534134
rect 280826 498218 281062 498454
rect 281146 498218 281382 498454
rect 280826 497898 281062 498134
rect 281146 497898 281382 498134
rect 280826 462218 281062 462454
rect 281146 462218 281382 462454
rect 280826 461898 281062 462134
rect 281146 461898 281382 462134
rect 280826 426218 281062 426454
rect 281146 426218 281382 426454
rect 280826 425898 281062 426134
rect 281146 425898 281382 426134
rect 280826 390218 281062 390454
rect 281146 390218 281382 390454
rect 280826 389898 281062 390134
rect 281146 389898 281382 390134
rect 280826 354218 281062 354454
rect 281146 354218 281382 354454
rect 280826 353898 281062 354134
rect 281146 353898 281382 354134
rect 280826 318218 281062 318454
rect 281146 318218 281382 318454
rect 280826 317898 281062 318134
rect 281146 317898 281382 318134
rect 280826 282218 281062 282454
rect 281146 282218 281382 282454
rect 280826 281898 281062 282134
rect 281146 281898 281382 282134
rect 285326 711322 285562 711558
rect 285646 711322 285882 711558
rect 285326 711002 285562 711238
rect 285646 711002 285882 711238
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 285326 610718 285562 610954
rect 285646 610718 285882 610954
rect 285326 610398 285562 610634
rect 285646 610398 285882 610634
rect 285326 574718 285562 574954
rect 285646 574718 285882 574954
rect 285326 574398 285562 574634
rect 285646 574398 285882 574634
rect 285326 538718 285562 538954
rect 285646 538718 285882 538954
rect 285326 538398 285562 538634
rect 285646 538398 285882 538634
rect 285326 502718 285562 502954
rect 285646 502718 285882 502954
rect 285326 502398 285562 502634
rect 285646 502398 285882 502634
rect 285326 466718 285562 466954
rect 285646 466718 285882 466954
rect 285326 466398 285562 466634
rect 285646 466398 285882 466634
rect 285326 430718 285562 430954
rect 285646 430718 285882 430954
rect 285326 430398 285562 430634
rect 285646 430398 285882 430634
rect 285326 394718 285562 394954
rect 285646 394718 285882 394954
rect 285326 394398 285562 394634
rect 285646 394398 285882 394634
rect 285326 358718 285562 358954
rect 285646 358718 285882 358954
rect 285326 358398 285562 358634
rect 285646 358398 285882 358634
rect 285326 322718 285562 322954
rect 285646 322718 285882 322954
rect 285326 322398 285562 322634
rect 285646 322398 285882 322634
rect 285326 286718 285562 286954
rect 285646 286718 285882 286954
rect 285326 286398 285562 286634
rect 285646 286398 285882 286634
rect 285326 250718 285562 250954
rect 285646 250718 285882 250954
rect 285326 250398 285562 250634
rect 285646 250398 285882 250634
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 294326 705562 294562 705798
rect 294646 705562 294882 705798
rect 294326 705242 294562 705478
rect 294646 705242 294882 705478
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 294326 619718 294562 619954
rect 294646 619718 294882 619954
rect 294326 619398 294562 619634
rect 294646 619398 294882 619634
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 294326 547718 294562 547954
rect 294646 547718 294882 547954
rect 294326 547398 294562 547634
rect 294646 547398 294882 547634
rect 294326 511718 294562 511954
rect 294646 511718 294882 511954
rect 294326 511398 294562 511634
rect 294646 511398 294882 511634
rect 294326 475718 294562 475954
rect 294646 475718 294882 475954
rect 294326 475398 294562 475634
rect 294646 475398 294882 475634
rect 294326 439718 294562 439954
rect 294646 439718 294882 439954
rect 294326 439398 294562 439634
rect 294646 439398 294882 439634
rect 294326 403718 294562 403954
rect 294646 403718 294882 403954
rect 294326 403398 294562 403634
rect 294646 403398 294882 403634
rect 294326 367718 294562 367954
rect 294646 367718 294882 367954
rect 294326 367398 294562 367634
rect 294646 367398 294882 367634
rect 294326 331718 294562 331954
rect 294646 331718 294882 331954
rect 294326 331398 294562 331634
rect 294646 331398 294882 331634
rect 294326 295718 294562 295954
rect 294646 295718 294882 295954
rect 294326 295398 294562 295634
rect 294646 295398 294882 295634
rect 294326 259718 294562 259954
rect 294646 259718 294882 259954
rect 294326 259398 294562 259634
rect 294646 259398 294882 259634
rect 298826 706522 299062 706758
rect 299146 706522 299382 706758
rect 298826 706202 299062 706438
rect 299146 706202 299382 706438
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 298826 660218 299062 660454
rect 299146 660218 299382 660454
rect 298826 659898 299062 660134
rect 299146 659898 299382 660134
rect 298826 624218 299062 624454
rect 299146 624218 299382 624454
rect 298826 623898 299062 624134
rect 299146 623898 299382 624134
rect 298826 588218 299062 588454
rect 299146 588218 299382 588454
rect 298826 587898 299062 588134
rect 299146 587898 299382 588134
rect 298826 552218 299062 552454
rect 299146 552218 299382 552454
rect 298826 551898 299062 552134
rect 299146 551898 299382 552134
rect 298826 516218 299062 516454
rect 299146 516218 299382 516454
rect 298826 515898 299062 516134
rect 299146 515898 299382 516134
rect 298826 480218 299062 480454
rect 299146 480218 299382 480454
rect 298826 479898 299062 480134
rect 299146 479898 299382 480134
rect 298826 444218 299062 444454
rect 299146 444218 299382 444454
rect 298826 443898 299062 444134
rect 299146 443898 299382 444134
rect 298826 408218 299062 408454
rect 299146 408218 299382 408454
rect 298826 407898 299062 408134
rect 299146 407898 299382 408134
rect 298826 372218 299062 372454
rect 299146 372218 299382 372454
rect 298826 371898 299062 372134
rect 299146 371898 299382 372134
rect 298826 336218 299062 336454
rect 299146 336218 299382 336454
rect 298826 335898 299062 336134
rect 299146 335898 299382 336134
rect 298826 300218 299062 300454
rect 299146 300218 299382 300454
rect 298826 299898 299062 300134
rect 299146 299898 299382 300134
rect 298826 264218 299062 264454
rect 299146 264218 299382 264454
rect 298826 263898 299062 264134
rect 299146 263898 299382 264134
rect 303326 707482 303562 707718
rect 303646 707482 303882 707718
rect 303326 707162 303562 707398
rect 303646 707162 303882 707398
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 303326 664718 303562 664954
rect 303646 664718 303882 664954
rect 303326 664398 303562 664634
rect 303646 664398 303882 664634
rect 303326 628718 303562 628954
rect 303646 628718 303882 628954
rect 303326 628398 303562 628634
rect 303646 628398 303882 628634
rect 303326 592718 303562 592954
rect 303646 592718 303882 592954
rect 303326 592398 303562 592634
rect 303646 592398 303882 592634
rect 303326 556718 303562 556954
rect 303646 556718 303882 556954
rect 303326 556398 303562 556634
rect 303646 556398 303882 556634
rect 303326 520718 303562 520954
rect 303646 520718 303882 520954
rect 303326 520398 303562 520634
rect 303646 520398 303882 520634
rect 303326 484718 303562 484954
rect 303646 484718 303882 484954
rect 303326 484398 303562 484634
rect 303646 484398 303882 484634
rect 303326 448718 303562 448954
rect 303646 448718 303882 448954
rect 303326 448398 303562 448634
rect 303646 448398 303882 448634
rect 303326 412718 303562 412954
rect 303646 412718 303882 412954
rect 303326 412398 303562 412634
rect 303646 412398 303882 412634
rect 303326 376718 303562 376954
rect 303646 376718 303882 376954
rect 303326 376398 303562 376634
rect 303646 376398 303882 376634
rect 303326 340718 303562 340954
rect 303646 340718 303882 340954
rect 303326 340398 303562 340634
rect 303646 340398 303882 340634
rect 303326 304718 303562 304954
rect 303646 304718 303882 304954
rect 303326 304398 303562 304634
rect 303646 304398 303882 304634
rect 303326 268718 303562 268954
rect 303646 268718 303882 268954
rect 303326 268398 303562 268634
rect 303646 268398 303882 268634
rect 307826 708442 308062 708678
rect 308146 708442 308382 708678
rect 307826 708122 308062 708358
rect 308146 708122 308382 708358
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 312326 709402 312562 709638
rect 312646 709402 312882 709638
rect 312326 709082 312562 709318
rect 312646 709082 312882 709318
rect 312326 673718 312562 673954
rect 312646 673718 312882 673954
rect 312326 673398 312562 673634
rect 312646 673398 312882 673634
rect 312326 637718 312562 637954
rect 312646 637718 312882 637954
rect 312326 637398 312562 637634
rect 312646 637398 312882 637634
rect 312326 601718 312562 601954
rect 312646 601718 312882 601954
rect 312326 601398 312562 601634
rect 312646 601398 312882 601634
rect 312326 565718 312562 565954
rect 312646 565718 312882 565954
rect 312326 565398 312562 565634
rect 312646 565398 312882 565634
rect 312326 529718 312562 529954
rect 312646 529718 312882 529954
rect 312326 529398 312562 529634
rect 312646 529398 312882 529634
rect 312326 493718 312562 493954
rect 312646 493718 312882 493954
rect 312326 493398 312562 493634
rect 312646 493398 312882 493634
rect 312326 457718 312562 457954
rect 312646 457718 312882 457954
rect 312326 457398 312562 457634
rect 312646 457398 312882 457634
rect 312326 421718 312562 421954
rect 312646 421718 312882 421954
rect 312326 421398 312562 421634
rect 312646 421398 312882 421634
rect 312326 385718 312562 385954
rect 312646 385718 312882 385954
rect 312326 385398 312562 385634
rect 312646 385398 312882 385634
rect 312326 349718 312562 349954
rect 312646 349718 312882 349954
rect 312326 349398 312562 349634
rect 312646 349398 312882 349634
rect 312326 313718 312562 313954
rect 312646 313718 312882 313954
rect 312326 313398 312562 313634
rect 312646 313398 312882 313634
rect 312326 277718 312562 277954
rect 312646 277718 312882 277954
rect 312326 277398 312562 277634
rect 312646 277398 312882 277634
rect 316826 710362 317062 710598
rect 317146 710362 317382 710598
rect 316826 710042 317062 710278
rect 317146 710042 317382 710278
rect 316826 678218 317062 678454
rect 317146 678218 317382 678454
rect 316826 677898 317062 678134
rect 317146 677898 317382 678134
rect 316826 642218 317062 642454
rect 317146 642218 317382 642454
rect 316826 641898 317062 642134
rect 317146 641898 317382 642134
rect 316826 606218 317062 606454
rect 317146 606218 317382 606454
rect 316826 605898 317062 606134
rect 317146 605898 317382 606134
rect 316826 570218 317062 570454
rect 317146 570218 317382 570454
rect 316826 569898 317062 570134
rect 317146 569898 317382 570134
rect 316826 534218 317062 534454
rect 317146 534218 317382 534454
rect 316826 533898 317062 534134
rect 317146 533898 317382 534134
rect 316826 498218 317062 498454
rect 317146 498218 317382 498454
rect 316826 497898 317062 498134
rect 317146 497898 317382 498134
rect 316826 462218 317062 462454
rect 317146 462218 317382 462454
rect 316826 461898 317062 462134
rect 317146 461898 317382 462134
rect 316826 426218 317062 426454
rect 317146 426218 317382 426454
rect 316826 425898 317062 426134
rect 317146 425898 317382 426134
rect 316826 390218 317062 390454
rect 317146 390218 317382 390454
rect 316826 389898 317062 390134
rect 317146 389898 317382 390134
rect 316826 354218 317062 354454
rect 317146 354218 317382 354454
rect 316826 353898 317062 354134
rect 317146 353898 317382 354134
rect 316826 318218 317062 318454
rect 317146 318218 317382 318454
rect 316826 317898 317062 318134
rect 317146 317898 317382 318134
rect 316826 282218 317062 282454
rect 317146 282218 317382 282454
rect 316826 281898 317062 282134
rect 317146 281898 317382 282134
rect 321326 711322 321562 711558
rect 321646 711322 321882 711558
rect 321326 711002 321562 711238
rect 321646 711002 321882 711238
rect 321326 682718 321562 682954
rect 321646 682718 321882 682954
rect 321326 682398 321562 682634
rect 321646 682398 321882 682634
rect 321326 646718 321562 646954
rect 321646 646718 321882 646954
rect 321326 646398 321562 646634
rect 321646 646398 321882 646634
rect 321326 610718 321562 610954
rect 321646 610718 321882 610954
rect 321326 610398 321562 610634
rect 321646 610398 321882 610634
rect 321326 574718 321562 574954
rect 321646 574718 321882 574954
rect 321326 574398 321562 574634
rect 321646 574398 321882 574634
rect 321326 538718 321562 538954
rect 321646 538718 321882 538954
rect 321326 538398 321562 538634
rect 321646 538398 321882 538634
rect 321326 502718 321562 502954
rect 321646 502718 321882 502954
rect 321326 502398 321562 502634
rect 321646 502398 321882 502634
rect 321326 466718 321562 466954
rect 321646 466718 321882 466954
rect 321326 466398 321562 466634
rect 321646 466398 321882 466634
rect 321326 430718 321562 430954
rect 321646 430718 321882 430954
rect 321326 430398 321562 430634
rect 321646 430398 321882 430634
rect 321326 394718 321562 394954
rect 321646 394718 321882 394954
rect 321326 394398 321562 394634
rect 321646 394398 321882 394634
rect 321326 358718 321562 358954
rect 321646 358718 321882 358954
rect 321326 358398 321562 358634
rect 321646 358398 321882 358634
rect 321326 322718 321562 322954
rect 321646 322718 321882 322954
rect 321326 322398 321562 322634
rect 321646 322398 321882 322634
rect 321326 286718 321562 286954
rect 321646 286718 321882 286954
rect 321326 286398 321562 286634
rect 321646 286398 321882 286634
rect 321326 250718 321562 250954
rect 321646 250718 321882 250954
rect 321326 250398 321562 250634
rect 321646 250398 321882 250634
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 330326 705562 330562 705798
rect 330646 705562 330882 705798
rect 330326 705242 330562 705478
rect 330646 705242 330882 705478
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 330326 655718 330562 655954
rect 330646 655718 330882 655954
rect 330326 655398 330562 655634
rect 330646 655398 330882 655634
rect 330326 619718 330562 619954
rect 330646 619718 330882 619954
rect 330326 619398 330562 619634
rect 330646 619398 330882 619634
rect 330326 583718 330562 583954
rect 330646 583718 330882 583954
rect 330326 583398 330562 583634
rect 330646 583398 330882 583634
rect 330326 547718 330562 547954
rect 330646 547718 330882 547954
rect 330326 547398 330562 547634
rect 330646 547398 330882 547634
rect 330326 511718 330562 511954
rect 330646 511718 330882 511954
rect 330326 511398 330562 511634
rect 330646 511398 330882 511634
rect 330326 475718 330562 475954
rect 330646 475718 330882 475954
rect 330326 475398 330562 475634
rect 330646 475398 330882 475634
rect 330326 439718 330562 439954
rect 330646 439718 330882 439954
rect 330326 439398 330562 439634
rect 330646 439398 330882 439634
rect 330326 403718 330562 403954
rect 330646 403718 330882 403954
rect 330326 403398 330562 403634
rect 330646 403398 330882 403634
rect 330326 367718 330562 367954
rect 330646 367718 330882 367954
rect 330326 367398 330562 367634
rect 330646 367398 330882 367634
rect 330326 331718 330562 331954
rect 330646 331718 330882 331954
rect 330326 331398 330562 331634
rect 330646 331398 330882 331634
rect 330326 295718 330562 295954
rect 330646 295718 330882 295954
rect 330326 295398 330562 295634
rect 330646 295398 330882 295634
rect 330326 259718 330562 259954
rect 330646 259718 330882 259954
rect 330326 259398 330562 259634
rect 330646 259398 330882 259634
rect 334826 706522 335062 706758
rect 335146 706522 335382 706758
rect 334826 706202 335062 706438
rect 335146 706202 335382 706438
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 334826 660218 335062 660454
rect 335146 660218 335382 660454
rect 334826 659898 335062 660134
rect 335146 659898 335382 660134
rect 334826 624218 335062 624454
rect 335146 624218 335382 624454
rect 334826 623898 335062 624134
rect 335146 623898 335382 624134
rect 334826 588218 335062 588454
rect 335146 588218 335382 588454
rect 334826 587898 335062 588134
rect 335146 587898 335382 588134
rect 334826 552218 335062 552454
rect 335146 552218 335382 552454
rect 334826 551898 335062 552134
rect 335146 551898 335382 552134
rect 334826 516218 335062 516454
rect 335146 516218 335382 516454
rect 334826 515898 335062 516134
rect 335146 515898 335382 516134
rect 334826 480218 335062 480454
rect 335146 480218 335382 480454
rect 334826 479898 335062 480134
rect 335146 479898 335382 480134
rect 334826 444218 335062 444454
rect 335146 444218 335382 444454
rect 334826 443898 335062 444134
rect 335146 443898 335382 444134
rect 334826 408218 335062 408454
rect 335146 408218 335382 408454
rect 334826 407898 335062 408134
rect 335146 407898 335382 408134
rect 334826 372218 335062 372454
rect 335146 372218 335382 372454
rect 334826 371898 335062 372134
rect 335146 371898 335382 372134
rect 334826 336218 335062 336454
rect 335146 336218 335382 336454
rect 334826 335898 335062 336134
rect 335146 335898 335382 336134
rect 334826 300218 335062 300454
rect 335146 300218 335382 300454
rect 334826 299898 335062 300134
rect 335146 299898 335382 300134
rect 334826 264218 335062 264454
rect 335146 264218 335382 264454
rect 334826 263898 335062 264134
rect 335146 263898 335382 264134
rect 339326 707482 339562 707718
rect 339646 707482 339882 707718
rect 339326 707162 339562 707398
rect 339646 707162 339882 707398
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 339326 664718 339562 664954
rect 339646 664718 339882 664954
rect 339326 664398 339562 664634
rect 339646 664398 339882 664634
rect 339326 628718 339562 628954
rect 339646 628718 339882 628954
rect 339326 628398 339562 628634
rect 339646 628398 339882 628634
rect 339326 592718 339562 592954
rect 339646 592718 339882 592954
rect 339326 592398 339562 592634
rect 339646 592398 339882 592634
rect 339326 556718 339562 556954
rect 339646 556718 339882 556954
rect 339326 556398 339562 556634
rect 339646 556398 339882 556634
rect 339326 520718 339562 520954
rect 339646 520718 339882 520954
rect 339326 520398 339562 520634
rect 339646 520398 339882 520634
rect 339326 484718 339562 484954
rect 339646 484718 339882 484954
rect 339326 484398 339562 484634
rect 339646 484398 339882 484634
rect 339326 448718 339562 448954
rect 339646 448718 339882 448954
rect 339326 448398 339562 448634
rect 339646 448398 339882 448634
rect 339326 412718 339562 412954
rect 339646 412718 339882 412954
rect 339326 412398 339562 412634
rect 339646 412398 339882 412634
rect 339326 376718 339562 376954
rect 339646 376718 339882 376954
rect 339326 376398 339562 376634
rect 339646 376398 339882 376634
rect 339326 340718 339562 340954
rect 339646 340718 339882 340954
rect 339326 340398 339562 340634
rect 339646 340398 339882 340634
rect 339326 304718 339562 304954
rect 339646 304718 339882 304954
rect 339326 304398 339562 304634
rect 339646 304398 339882 304634
rect 339326 268718 339562 268954
rect 339646 268718 339882 268954
rect 339326 268398 339562 268634
rect 339646 268398 339882 268634
rect 343826 708442 344062 708678
rect 344146 708442 344382 708678
rect 343826 708122 344062 708358
rect 344146 708122 344382 708358
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 348326 709402 348562 709638
rect 348646 709402 348882 709638
rect 348326 709082 348562 709318
rect 348646 709082 348882 709318
rect 348326 673718 348562 673954
rect 348646 673718 348882 673954
rect 348326 673398 348562 673634
rect 348646 673398 348882 673634
rect 348326 637718 348562 637954
rect 348646 637718 348882 637954
rect 348326 637398 348562 637634
rect 348646 637398 348882 637634
rect 348326 601718 348562 601954
rect 348646 601718 348882 601954
rect 348326 601398 348562 601634
rect 348646 601398 348882 601634
rect 348326 565718 348562 565954
rect 348646 565718 348882 565954
rect 348326 565398 348562 565634
rect 348646 565398 348882 565634
rect 348326 529718 348562 529954
rect 348646 529718 348882 529954
rect 348326 529398 348562 529634
rect 348646 529398 348882 529634
rect 348326 493718 348562 493954
rect 348646 493718 348882 493954
rect 348326 493398 348562 493634
rect 348646 493398 348882 493634
rect 348326 457718 348562 457954
rect 348646 457718 348882 457954
rect 348326 457398 348562 457634
rect 348646 457398 348882 457634
rect 348326 421718 348562 421954
rect 348646 421718 348882 421954
rect 348326 421398 348562 421634
rect 348646 421398 348882 421634
rect 348326 385718 348562 385954
rect 348646 385718 348882 385954
rect 348326 385398 348562 385634
rect 348646 385398 348882 385634
rect 348326 349718 348562 349954
rect 348646 349718 348882 349954
rect 348326 349398 348562 349634
rect 348646 349398 348882 349634
rect 348326 313718 348562 313954
rect 348646 313718 348882 313954
rect 348326 313398 348562 313634
rect 348646 313398 348882 313634
rect 348326 277718 348562 277954
rect 348646 277718 348882 277954
rect 348326 277398 348562 277634
rect 348646 277398 348882 277634
rect 352826 710362 353062 710598
rect 353146 710362 353382 710598
rect 352826 710042 353062 710278
rect 353146 710042 353382 710278
rect 352826 678218 353062 678454
rect 353146 678218 353382 678454
rect 352826 677898 353062 678134
rect 353146 677898 353382 678134
rect 352826 642218 353062 642454
rect 353146 642218 353382 642454
rect 352826 641898 353062 642134
rect 353146 641898 353382 642134
rect 352826 606218 353062 606454
rect 353146 606218 353382 606454
rect 352826 605898 353062 606134
rect 353146 605898 353382 606134
rect 352826 570218 353062 570454
rect 353146 570218 353382 570454
rect 352826 569898 353062 570134
rect 353146 569898 353382 570134
rect 352826 534218 353062 534454
rect 353146 534218 353382 534454
rect 352826 533898 353062 534134
rect 353146 533898 353382 534134
rect 352826 498218 353062 498454
rect 353146 498218 353382 498454
rect 352826 497898 353062 498134
rect 353146 497898 353382 498134
rect 352826 462218 353062 462454
rect 353146 462218 353382 462454
rect 352826 461898 353062 462134
rect 353146 461898 353382 462134
rect 352826 426218 353062 426454
rect 353146 426218 353382 426454
rect 352826 425898 353062 426134
rect 353146 425898 353382 426134
rect 352826 390218 353062 390454
rect 353146 390218 353382 390454
rect 352826 389898 353062 390134
rect 353146 389898 353382 390134
rect 352826 354218 353062 354454
rect 353146 354218 353382 354454
rect 352826 353898 353062 354134
rect 353146 353898 353382 354134
rect 352826 318218 353062 318454
rect 353146 318218 353382 318454
rect 352826 317898 353062 318134
rect 353146 317898 353382 318134
rect 352826 282218 353062 282454
rect 353146 282218 353382 282454
rect 352826 281898 353062 282134
rect 353146 281898 353382 282134
rect 357326 711322 357562 711558
rect 357646 711322 357882 711558
rect 357326 711002 357562 711238
rect 357646 711002 357882 711238
rect 357326 682718 357562 682954
rect 357646 682718 357882 682954
rect 357326 682398 357562 682634
rect 357646 682398 357882 682634
rect 357326 646718 357562 646954
rect 357646 646718 357882 646954
rect 357326 646398 357562 646634
rect 357646 646398 357882 646634
rect 357326 610718 357562 610954
rect 357646 610718 357882 610954
rect 357326 610398 357562 610634
rect 357646 610398 357882 610634
rect 357326 574718 357562 574954
rect 357646 574718 357882 574954
rect 357326 574398 357562 574634
rect 357646 574398 357882 574634
rect 357326 538718 357562 538954
rect 357646 538718 357882 538954
rect 357326 538398 357562 538634
rect 357646 538398 357882 538634
rect 357326 502718 357562 502954
rect 357646 502718 357882 502954
rect 357326 502398 357562 502634
rect 357646 502398 357882 502634
rect 357326 466718 357562 466954
rect 357646 466718 357882 466954
rect 357326 466398 357562 466634
rect 357646 466398 357882 466634
rect 357326 430718 357562 430954
rect 357646 430718 357882 430954
rect 357326 430398 357562 430634
rect 357646 430398 357882 430634
rect 357326 394718 357562 394954
rect 357646 394718 357882 394954
rect 357326 394398 357562 394634
rect 357646 394398 357882 394634
rect 357326 358718 357562 358954
rect 357646 358718 357882 358954
rect 357326 358398 357562 358634
rect 357646 358398 357882 358634
rect 357326 322718 357562 322954
rect 357646 322718 357882 322954
rect 357326 322398 357562 322634
rect 357646 322398 357882 322634
rect 357326 286718 357562 286954
rect 357646 286718 357882 286954
rect 357326 286398 357562 286634
rect 357646 286398 357882 286634
rect 357326 250718 357562 250954
rect 357646 250718 357882 250954
rect 357326 250398 357562 250634
rect 357646 250398 357882 250634
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 366326 705562 366562 705798
rect 366646 705562 366882 705798
rect 366326 705242 366562 705478
rect 366646 705242 366882 705478
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 366326 655718 366562 655954
rect 366646 655718 366882 655954
rect 366326 655398 366562 655634
rect 366646 655398 366882 655634
rect 366326 619718 366562 619954
rect 366646 619718 366882 619954
rect 366326 619398 366562 619634
rect 366646 619398 366882 619634
rect 366326 583718 366562 583954
rect 366646 583718 366882 583954
rect 366326 583398 366562 583634
rect 366646 583398 366882 583634
rect 366326 547718 366562 547954
rect 366646 547718 366882 547954
rect 366326 547398 366562 547634
rect 366646 547398 366882 547634
rect 366326 511718 366562 511954
rect 366646 511718 366882 511954
rect 366326 511398 366562 511634
rect 366646 511398 366882 511634
rect 366326 475718 366562 475954
rect 366646 475718 366882 475954
rect 366326 475398 366562 475634
rect 366646 475398 366882 475634
rect 366326 439718 366562 439954
rect 366646 439718 366882 439954
rect 366326 439398 366562 439634
rect 366646 439398 366882 439634
rect 366326 403718 366562 403954
rect 366646 403718 366882 403954
rect 366326 403398 366562 403634
rect 366646 403398 366882 403634
rect 366326 367718 366562 367954
rect 366646 367718 366882 367954
rect 366326 367398 366562 367634
rect 366646 367398 366882 367634
rect 366326 331718 366562 331954
rect 366646 331718 366882 331954
rect 366326 331398 366562 331634
rect 366646 331398 366882 331634
rect 366326 295718 366562 295954
rect 366646 295718 366882 295954
rect 366326 295398 366562 295634
rect 366646 295398 366882 295634
rect 366326 259718 366562 259954
rect 366646 259718 366882 259954
rect 366326 259398 366562 259634
rect 366646 259398 366882 259634
rect 370826 706522 371062 706758
rect 371146 706522 371382 706758
rect 370826 706202 371062 706438
rect 371146 706202 371382 706438
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 370826 660218 371062 660454
rect 371146 660218 371382 660454
rect 370826 659898 371062 660134
rect 371146 659898 371382 660134
rect 370826 624218 371062 624454
rect 371146 624218 371382 624454
rect 370826 623898 371062 624134
rect 371146 623898 371382 624134
rect 370826 588218 371062 588454
rect 371146 588218 371382 588454
rect 370826 587898 371062 588134
rect 371146 587898 371382 588134
rect 370826 552218 371062 552454
rect 371146 552218 371382 552454
rect 370826 551898 371062 552134
rect 371146 551898 371382 552134
rect 370826 516218 371062 516454
rect 371146 516218 371382 516454
rect 370826 515898 371062 516134
rect 371146 515898 371382 516134
rect 370826 480218 371062 480454
rect 371146 480218 371382 480454
rect 370826 479898 371062 480134
rect 371146 479898 371382 480134
rect 370826 444218 371062 444454
rect 371146 444218 371382 444454
rect 370826 443898 371062 444134
rect 371146 443898 371382 444134
rect 370826 408218 371062 408454
rect 371146 408218 371382 408454
rect 370826 407898 371062 408134
rect 371146 407898 371382 408134
rect 370826 372218 371062 372454
rect 371146 372218 371382 372454
rect 370826 371898 371062 372134
rect 371146 371898 371382 372134
rect 370826 336218 371062 336454
rect 371146 336218 371382 336454
rect 370826 335898 371062 336134
rect 371146 335898 371382 336134
rect 370826 300218 371062 300454
rect 371146 300218 371382 300454
rect 370826 299898 371062 300134
rect 371146 299898 371382 300134
rect 370826 264218 371062 264454
rect 371146 264218 371382 264454
rect 370826 263898 371062 264134
rect 371146 263898 371382 264134
rect 375326 707482 375562 707718
rect 375646 707482 375882 707718
rect 375326 707162 375562 707398
rect 375646 707162 375882 707398
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 375326 664718 375562 664954
rect 375646 664718 375882 664954
rect 375326 664398 375562 664634
rect 375646 664398 375882 664634
rect 375326 628718 375562 628954
rect 375646 628718 375882 628954
rect 375326 628398 375562 628634
rect 375646 628398 375882 628634
rect 375326 592718 375562 592954
rect 375646 592718 375882 592954
rect 375326 592398 375562 592634
rect 375646 592398 375882 592634
rect 375326 556718 375562 556954
rect 375646 556718 375882 556954
rect 375326 556398 375562 556634
rect 375646 556398 375882 556634
rect 375326 520718 375562 520954
rect 375646 520718 375882 520954
rect 375326 520398 375562 520634
rect 375646 520398 375882 520634
rect 375326 484718 375562 484954
rect 375646 484718 375882 484954
rect 375326 484398 375562 484634
rect 375646 484398 375882 484634
rect 375326 448718 375562 448954
rect 375646 448718 375882 448954
rect 375326 448398 375562 448634
rect 375646 448398 375882 448634
rect 375326 412718 375562 412954
rect 375646 412718 375882 412954
rect 375326 412398 375562 412634
rect 375646 412398 375882 412634
rect 375326 376718 375562 376954
rect 375646 376718 375882 376954
rect 375326 376398 375562 376634
rect 375646 376398 375882 376634
rect 375326 340718 375562 340954
rect 375646 340718 375882 340954
rect 375326 340398 375562 340634
rect 375646 340398 375882 340634
rect 375326 304718 375562 304954
rect 375646 304718 375882 304954
rect 375326 304398 375562 304634
rect 375646 304398 375882 304634
rect 375326 268718 375562 268954
rect 375646 268718 375882 268954
rect 375326 268398 375562 268634
rect 375646 268398 375882 268634
rect 379826 708442 380062 708678
rect 380146 708442 380382 708678
rect 379826 708122 380062 708358
rect 380146 708122 380382 708358
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 384326 709402 384562 709638
rect 384646 709402 384882 709638
rect 384326 709082 384562 709318
rect 384646 709082 384882 709318
rect 384326 673718 384562 673954
rect 384646 673718 384882 673954
rect 384326 673398 384562 673634
rect 384646 673398 384882 673634
rect 384326 637718 384562 637954
rect 384646 637718 384882 637954
rect 384326 637398 384562 637634
rect 384646 637398 384882 637634
rect 384326 601718 384562 601954
rect 384646 601718 384882 601954
rect 384326 601398 384562 601634
rect 384646 601398 384882 601634
rect 384326 565718 384562 565954
rect 384646 565718 384882 565954
rect 384326 565398 384562 565634
rect 384646 565398 384882 565634
rect 384326 529718 384562 529954
rect 384646 529718 384882 529954
rect 384326 529398 384562 529634
rect 384646 529398 384882 529634
rect 384326 493718 384562 493954
rect 384646 493718 384882 493954
rect 384326 493398 384562 493634
rect 384646 493398 384882 493634
rect 384326 457718 384562 457954
rect 384646 457718 384882 457954
rect 384326 457398 384562 457634
rect 384646 457398 384882 457634
rect 384326 421718 384562 421954
rect 384646 421718 384882 421954
rect 384326 421398 384562 421634
rect 384646 421398 384882 421634
rect 384326 385718 384562 385954
rect 384646 385718 384882 385954
rect 384326 385398 384562 385634
rect 384646 385398 384882 385634
rect 384326 349718 384562 349954
rect 384646 349718 384882 349954
rect 384326 349398 384562 349634
rect 384646 349398 384882 349634
rect 384326 313718 384562 313954
rect 384646 313718 384882 313954
rect 384326 313398 384562 313634
rect 384646 313398 384882 313634
rect 384326 277718 384562 277954
rect 384646 277718 384882 277954
rect 384326 277398 384562 277634
rect 384646 277398 384882 277634
rect 388826 710362 389062 710598
rect 389146 710362 389382 710598
rect 388826 710042 389062 710278
rect 389146 710042 389382 710278
rect 388826 678218 389062 678454
rect 389146 678218 389382 678454
rect 388826 677898 389062 678134
rect 389146 677898 389382 678134
rect 388826 642218 389062 642454
rect 389146 642218 389382 642454
rect 388826 641898 389062 642134
rect 389146 641898 389382 642134
rect 388826 606218 389062 606454
rect 389146 606218 389382 606454
rect 388826 605898 389062 606134
rect 389146 605898 389382 606134
rect 388826 570218 389062 570454
rect 389146 570218 389382 570454
rect 388826 569898 389062 570134
rect 389146 569898 389382 570134
rect 388826 534218 389062 534454
rect 389146 534218 389382 534454
rect 388826 533898 389062 534134
rect 389146 533898 389382 534134
rect 388826 498218 389062 498454
rect 389146 498218 389382 498454
rect 388826 497898 389062 498134
rect 389146 497898 389382 498134
rect 388826 462218 389062 462454
rect 389146 462218 389382 462454
rect 388826 461898 389062 462134
rect 389146 461898 389382 462134
rect 388826 426218 389062 426454
rect 389146 426218 389382 426454
rect 388826 425898 389062 426134
rect 389146 425898 389382 426134
rect 388826 390218 389062 390454
rect 389146 390218 389382 390454
rect 388826 389898 389062 390134
rect 389146 389898 389382 390134
rect 388826 354218 389062 354454
rect 389146 354218 389382 354454
rect 388826 353898 389062 354134
rect 389146 353898 389382 354134
rect 388826 318218 389062 318454
rect 389146 318218 389382 318454
rect 388826 317898 389062 318134
rect 389146 317898 389382 318134
rect 388826 282218 389062 282454
rect 389146 282218 389382 282454
rect 388826 281898 389062 282134
rect 389146 281898 389382 282134
rect 393326 711322 393562 711558
rect 393646 711322 393882 711558
rect 393326 711002 393562 711238
rect 393646 711002 393882 711238
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 393326 610718 393562 610954
rect 393646 610718 393882 610954
rect 393326 610398 393562 610634
rect 393646 610398 393882 610634
rect 393326 574718 393562 574954
rect 393646 574718 393882 574954
rect 393326 574398 393562 574634
rect 393646 574398 393882 574634
rect 393326 538718 393562 538954
rect 393646 538718 393882 538954
rect 393326 538398 393562 538634
rect 393646 538398 393882 538634
rect 393326 502718 393562 502954
rect 393646 502718 393882 502954
rect 393326 502398 393562 502634
rect 393646 502398 393882 502634
rect 393326 466718 393562 466954
rect 393646 466718 393882 466954
rect 393326 466398 393562 466634
rect 393646 466398 393882 466634
rect 393326 430718 393562 430954
rect 393646 430718 393882 430954
rect 393326 430398 393562 430634
rect 393646 430398 393882 430634
rect 393326 394718 393562 394954
rect 393646 394718 393882 394954
rect 393326 394398 393562 394634
rect 393646 394398 393882 394634
rect 393326 358718 393562 358954
rect 393646 358718 393882 358954
rect 393326 358398 393562 358634
rect 393646 358398 393882 358634
rect 393326 322718 393562 322954
rect 393646 322718 393882 322954
rect 393326 322398 393562 322634
rect 393646 322398 393882 322634
rect 393326 286718 393562 286954
rect 393646 286718 393882 286954
rect 393326 286398 393562 286634
rect 393646 286398 393882 286634
rect 393326 250718 393562 250954
rect 393646 250718 393882 250954
rect 393326 250398 393562 250634
rect 393646 250398 393882 250634
rect 65342 246067 65578 246303
rect 65662 246067 65898 246303
rect 65982 246067 66218 246303
rect 66302 246067 66538 246303
rect 66622 246067 66858 246303
rect 66942 246067 67178 246303
rect 67262 246067 67498 246303
rect 67582 246067 67818 246303
rect 67902 246067 68138 246303
rect 68222 246067 68458 246303
rect 68542 246067 68778 246303
rect 68862 246067 69098 246303
rect 69182 246067 69418 246303
rect 69502 246067 69738 246303
rect 69822 246067 70058 246303
rect 65462 241717 65698 241953
rect 65782 241717 66018 241953
rect 66102 241717 66338 241953
rect 66422 241717 66658 241953
rect 66742 241717 66978 241953
rect 67062 241717 67298 241953
rect 67382 241717 67618 241953
rect 67702 241717 67938 241953
rect 68022 241717 68258 241953
rect 68342 241717 68578 241953
rect 68662 241717 68898 241953
rect 68982 241717 69218 241953
rect 69302 241717 69538 241953
rect 69622 241717 69858 241953
rect 69942 241717 70178 241953
rect 70262 241717 70498 241953
rect 70582 241717 70818 241953
rect 70902 241717 71138 241953
rect 65462 241397 65698 241633
rect 65782 241397 66018 241633
rect 66102 241397 66338 241633
rect 66422 241397 66658 241633
rect 66742 241397 66978 241633
rect 67062 241397 67298 241633
rect 67382 241397 67618 241633
rect 67702 241397 67938 241633
rect 68022 241397 68258 241633
rect 68342 241397 68578 241633
rect 68662 241397 68898 241633
rect 68982 241397 69218 241633
rect 69302 241397 69538 241633
rect 69622 241397 69858 241633
rect 69942 241397 70178 241633
rect 70262 241397 70498 241633
rect 70582 241397 70818 241633
rect 70902 241397 71138 241633
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 42326 151718 42562 151954
rect 42646 151718 42882 151954
rect 42326 151398 42562 151634
rect 42646 151398 42882 151634
rect 42326 115718 42562 115954
rect 42646 115718 42882 115954
rect 42326 115398 42562 115634
rect 42646 115398 42882 115634
rect 42326 79718 42562 79954
rect 42646 79718 42882 79954
rect 42326 79398 42562 79634
rect 42646 79398 42882 79634
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1542 42562 -1306
rect 42646 -1542 42882 -1306
rect 42326 -1862 42562 -1626
rect 42646 -1862 42882 -1626
rect 46826 228217 47062 228453
rect 47146 228217 47382 228453
rect 46826 227897 47062 228133
rect 47146 227897 47382 228133
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 46826 84218 47062 84454
rect 47146 84218 47382 84454
rect 46826 83898 47062 84134
rect 47146 83898 47382 84134
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2502 47062 -2266
rect 47146 -2502 47382 -2266
rect 46826 -2822 47062 -2586
rect 47146 -2822 47382 -2586
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 51326 124718 51562 124954
rect 51646 124718 51882 124954
rect 51326 124398 51562 124634
rect 51646 124398 51882 124634
rect 51326 88718 51562 88954
rect 51646 88718 51882 88954
rect 51326 88398 51562 88634
rect 51646 88398 51882 88634
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3462 51562 -3226
rect 51646 -3462 51882 -3226
rect 51326 -3782 51562 -3546
rect 51646 -3782 51882 -3546
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4422 56062 -4186
rect 56146 -4422 56382 -4186
rect 55826 -4742 56062 -4506
rect 56146 -4742 56382 -4506
rect 60326 205718 60562 205954
rect 60646 205718 60882 205954
rect 60326 205398 60562 205634
rect 60646 205398 60882 205634
rect 60326 169718 60562 169954
rect 60646 169718 60882 169954
rect 60326 169398 60562 169634
rect 60646 169398 60882 169634
rect 60326 133718 60562 133954
rect 60646 133718 60882 133954
rect 60326 133398 60562 133634
rect 60646 133398 60882 133634
rect 60326 97718 60562 97954
rect 60646 97718 60882 97954
rect 60326 97398 60562 97634
rect 60646 97398 60882 97634
rect 60326 61718 60562 61954
rect 60646 61718 60882 61954
rect 60326 61398 60562 61634
rect 60646 61398 60882 61634
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 60326 -5382 60562 -5146
rect 60646 -5382 60882 -5146
rect 60326 -5702 60562 -5466
rect 60646 -5702 60882 -5466
rect 64826 210218 65062 210454
rect 65146 210218 65382 210454
rect 64826 209898 65062 210134
rect 65146 209898 65382 210134
rect 64826 174218 65062 174454
rect 65146 174218 65382 174454
rect 64826 173898 65062 174134
rect 65146 173898 65382 174134
rect 64826 138218 65062 138454
rect 65146 138218 65382 138454
rect 64826 137898 65062 138134
rect 65146 137898 65382 138134
rect 64826 102218 65062 102454
rect 65146 102218 65382 102454
rect 64826 101898 65062 102134
rect 65146 101898 65382 102134
rect 64826 66218 65062 66454
rect 65146 66218 65382 66454
rect 64826 65898 65062 66134
rect 65146 65898 65382 66134
rect 64826 30218 65062 30454
rect 65146 30218 65382 30454
rect 64826 29898 65062 30134
rect 65146 29898 65382 30134
rect 64826 -6342 65062 -6106
rect 65146 -6342 65382 -6106
rect 64826 -6662 65062 -6426
rect 65146 -6662 65382 -6426
rect 69326 214718 69562 214954
rect 69646 214718 69882 214954
rect 69326 214398 69562 214634
rect 69646 214398 69882 214634
rect 69326 178718 69562 178954
rect 69646 178718 69882 178954
rect 69326 178398 69562 178634
rect 69646 178398 69882 178634
rect 69326 142718 69562 142954
rect 69646 142718 69882 142954
rect 69326 142398 69562 142634
rect 69646 142398 69882 142634
rect 69326 106718 69562 106954
rect 69646 106718 69882 106954
rect 69326 106398 69562 106634
rect 69646 106398 69882 106634
rect 69326 70718 69562 70954
rect 69646 70718 69882 70954
rect 69326 70398 69562 70634
rect 69646 70398 69882 70634
rect 69326 34718 69562 34954
rect 69646 34718 69882 34954
rect 69326 34398 69562 34634
rect 69646 34398 69882 34634
rect 69326 -7302 69562 -7066
rect 69646 -7302 69882 -7066
rect 69326 -7622 69562 -7386
rect 69646 -7622 69882 -7386
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 78326 223718 78562 223954
rect 78646 223718 78882 223954
rect 78326 223398 78562 223634
rect 78646 223398 78882 223634
rect 78326 187718 78562 187954
rect 78646 187718 78882 187954
rect 78326 187398 78562 187634
rect 78646 187398 78882 187634
rect 78326 151718 78562 151954
rect 78646 151718 78882 151954
rect 78326 151398 78562 151634
rect 78646 151398 78882 151634
rect 78326 115718 78562 115954
rect 78646 115718 78882 115954
rect 78326 115398 78562 115634
rect 78646 115398 78882 115634
rect 78326 79718 78562 79954
rect 78646 79718 78882 79954
rect 78326 79398 78562 79634
rect 78646 79398 78882 79634
rect 78326 43718 78562 43954
rect 78646 43718 78882 43954
rect 78326 43398 78562 43634
rect 78646 43398 78882 43634
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1542 78562 -1306
rect 78646 -1542 78882 -1306
rect 78326 -1862 78562 -1626
rect 78646 -1862 78882 -1626
rect 82826 228217 83062 228453
rect 83146 228217 83382 228453
rect 82826 227897 83062 228133
rect 83146 227897 83382 228133
rect 82826 192218 83062 192454
rect 83146 192218 83382 192454
rect 82826 191898 83062 192134
rect 83146 191898 83382 192134
rect 82826 156218 83062 156454
rect 83146 156218 83382 156454
rect 82826 155898 83062 156134
rect 83146 155898 83382 156134
rect 82826 120218 83062 120454
rect 83146 120218 83382 120454
rect 82826 119898 83062 120134
rect 83146 119898 83382 120134
rect 82826 84218 83062 84454
rect 83146 84218 83382 84454
rect 82826 83898 83062 84134
rect 83146 83898 83382 84134
rect 82826 48218 83062 48454
rect 83146 48218 83382 48454
rect 82826 47898 83062 48134
rect 83146 47898 83382 48134
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2502 83062 -2266
rect 83146 -2502 83382 -2266
rect 82826 -2822 83062 -2586
rect 83146 -2822 83382 -2586
rect 87326 196718 87562 196954
rect 87646 196718 87882 196954
rect 87326 196398 87562 196634
rect 87646 196398 87882 196634
rect 87326 160718 87562 160954
rect 87646 160718 87882 160954
rect 87326 160398 87562 160634
rect 87646 160398 87882 160634
rect 87326 124718 87562 124954
rect 87646 124718 87882 124954
rect 87326 124398 87562 124634
rect 87646 124398 87882 124634
rect 87326 88718 87562 88954
rect 87646 88718 87882 88954
rect 87326 88398 87562 88634
rect 87646 88398 87882 88634
rect 87326 52718 87562 52954
rect 87646 52718 87882 52954
rect 87326 52398 87562 52634
rect 87646 52398 87882 52634
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3462 87562 -3226
rect 87646 -3462 87882 -3226
rect 87326 -3782 87562 -3546
rect 87646 -3782 87882 -3546
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4422 92062 -4186
rect 92146 -4422 92382 -4186
rect 91826 -4742 92062 -4506
rect 92146 -4742 92382 -4506
rect 96326 205718 96562 205954
rect 96646 205718 96882 205954
rect 96326 205398 96562 205634
rect 96646 205398 96882 205634
rect 96326 169718 96562 169954
rect 96646 169718 96882 169954
rect 96326 169398 96562 169634
rect 96646 169398 96882 169634
rect 96326 133718 96562 133954
rect 96646 133718 96882 133954
rect 96326 133398 96562 133634
rect 96646 133398 96882 133634
rect 96326 97718 96562 97954
rect 96646 97718 96882 97954
rect 96326 97398 96562 97634
rect 96646 97398 96882 97634
rect 96326 61718 96562 61954
rect 96646 61718 96882 61954
rect 96326 61398 96562 61634
rect 96646 61398 96882 61634
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 96326 -5382 96562 -5146
rect 96646 -5382 96882 -5146
rect 96326 -5702 96562 -5466
rect 96646 -5702 96882 -5466
rect 100826 210218 101062 210454
rect 101146 210218 101382 210454
rect 100826 209898 101062 210134
rect 101146 209898 101382 210134
rect 100826 174218 101062 174454
rect 101146 174218 101382 174454
rect 100826 173898 101062 174134
rect 101146 173898 101382 174134
rect 100826 138218 101062 138454
rect 101146 138218 101382 138454
rect 100826 137898 101062 138134
rect 101146 137898 101382 138134
rect 100826 102218 101062 102454
rect 101146 102218 101382 102454
rect 100826 101898 101062 102134
rect 101146 101898 101382 102134
rect 100826 66218 101062 66454
rect 101146 66218 101382 66454
rect 100826 65898 101062 66134
rect 101146 65898 101382 66134
rect 100826 30218 101062 30454
rect 101146 30218 101382 30454
rect 100826 29898 101062 30134
rect 101146 29898 101382 30134
rect 100826 -6342 101062 -6106
rect 101146 -6342 101382 -6106
rect 100826 -6662 101062 -6426
rect 101146 -6662 101382 -6426
rect 105326 214718 105562 214954
rect 105646 214718 105882 214954
rect 105326 214398 105562 214634
rect 105646 214398 105882 214634
rect 105326 178718 105562 178954
rect 105646 178718 105882 178954
rect 105326 178398 105562 178634
rect 105646 178398 105882 178634
rect 105326 142718 105562 142954
rect 105646 142718 105882 142954
rect 105326 142398 105562 142634
rect 105646 142398 105882 142634
rect 105326 106718 105562 106954
rect 105646 106718 105882 106954
rect 105326 106398 105562 106634
rect 105646 106398 105882 106634
rect 105326 70718 105562 70954
rect 105646 70718 105882 70954
rect 105326 70398 105562 70634
rect 105646 70398 105882 70634
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 105326 -7302 105562 -7066
rect 105646 -7302 105882 -7066
rect 105326 -7622 105562 -7386
rect 105646 -7622 105882 -7386
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 114326 223718 114562 223954
rect 114646 223718 114882 223954
rect 114326 223398 114562 223634
rect 114646 223398 114882 223634
rect 114326 187718 114562 187954
rect 114646 187718 114882 187954
rect 114326 187398 114562 187634
rect 114646 187398 114882 187634
rect 114326 151718 114562 151954
rect 114646 151718 114882 151954
rect 114326 151398 114562 151634
rect 114646 151398 114882 151634
rect 118826 228217 119062 228453
rect 119146 228217 119382 228453
rect 118826 227897 119062 228133
rect 119146 227897 119382 228133
rect 118826 192218 119062 192454
rect 119146 192218 119382 192454
rect 118826 191898 119062 192134
rect 119146 191898 119382 192134
rect 118826 156218 119062 156454
rect 119146 156218 119382 156454
rect 118826 155898 119062 156134
rect 119146 155898 119382 156134
rect 123326 196718 123562 196954
rect 123646 196718 123882 196954
rect 123326 196398 123562 196634
rect 123646 196398 123882 196634
rect 123326 160718 123562 160954
rect 123646 160718 123882 160954
rect 123326 160398 123562 160634
rect 123646 160398 123882 160634
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 172826 210218 173062 210454
rect 173146 210218 173382 210454
rect 172826 209898 173062 210134
rect 173146 209898 173382 210134
rect 132326 205718 132562 205954
rect 132646 205718 132882 205954
rect 132326 205398 132562 205634
rect 132646 205398 132882 205634
rect 136036 205625 136272 205861
rect 136356 205625 136592 205861
rect 136676 205625 136912 205861
rect 136996 205625 137232 205861
rect 137316 205625 137552 205861
rect 137636 205625 137872 205861
rect 137956 205625 138192 205861
rect 138276 205625 138512 205861
rect 138596 205625 138832 205861
rect 138916 205625 139152 205861
rect 139236 205625 139472 205861
rect 139556 205625 139792 205861
rect 139876 205625 140112 205861
rect 140196 205625 140432 205861
rect 140516 205625 140752 205861
rect 140836 205625 141072 205861
rect 141156 205625 141392 205861
rect 141476 205625 141712 205861
rect 141796 205625 142032 205861
rect 142116 205625 142352 205861
rect 142436 205625 142672 205861
rect 142756 205625 142992 205861
rect 143076 205625 143312 205861
rect 143396 205625 143632 205861
rect 143716 205625 143952 205861
rect 144036 205625 144272 205861
rect 144356 205625 144592 205861
rect 144676 205625 144912 205861
rect 144996 205625 145232 205861
rect 145316 205625 145552 205861
rect 145636 205625 145872 205861
rect 145956 205625 146192 205861
rect 146276 205625 146512 205861
rect 146596 205625 146832 205861
rect 146916 205625 147152 205861
rect 147236 205625 147472 205861
rect 147556 205625 147792 205861
rect 147876 205625 148112 205861
rect 148196 205625 148432 205861
rect 148516 205625 148752 205861
rect 148836 205625 149072 205861
rect 149156 205625 149392 205861
rect 149476 205625 149712 205861
rect 149796 205625 150032 205861
rect 150116 205625 150352 205861
rect 150436 205625 150672 205861
rect 150756 205625 150992 205861
rect 151076 205625 151312 205861
rect 151396 205625 151632 205861
rect 151716 205625 151952 205861
rect 152036 205625 152272 205861
rect 152356 205625 152592 205861
rect 152676 205625 152912 205861
rect 152996 205625 153232 205861
rect 153316 205625 153552 205861
rect 153636 205625 153872 205861
rect 153956 205625 154192 205861
rect 154276 205625 154512 205861
rect 154596 205625 154832 205861
rect 154916 205625 155152 205861
rect 155236 205625 155472 205861
rect 155556 205625 155792 205861
rect 155876 205625 156112 205861
rect 156196 205625 156432 205861
rect 156516 205625 156752 205861
rect 156836 205625 157072 205861
rect 157156 205625 157392 205861
rect 157476 205625 157712 205861
rect 157796 205625 158032 205861
rect 158116 205625 158352 205861
rect 158436 205625 158672 205861
rect 158756 205625 158992 205861
rect 159076 205625 159312 205861
rect 159396 205625 159632 205861
rect 159716 205625 159952 205861
rect 160036 205625 160272 205861
rect 160356 205625 160592 205861
rect 160676 205625 160912 205861
rect 160996 205625 161232 205861
rect 161316 205625 161552 205861
rect 161636 205625 161872 205861
rect 161956 205625 162192 205861
rect 162276 205625 162512 205861
rect 162596 205625 162832 205861
rect 162916 205625 163152 205861
rect 163236 205625 163472 205861
rect 163556 205625 163792 205861
rect 163876 205625 164112 205861
rect 164196 205625 164432 205861
rect 164516 205625 164752 205861
rect 164836 205625 165072 205861
rect 165156 205625 165392 205861
rect 137376 201175 137612 201411
rect 137696 201175 137932 201411
rect 138016 201175 138252 201411
rect 138336 201175 138572 201411
rect 138656 201175 138892 201411
rect 138976 201175 139212 201411
rect 139296 201175 139532 201411
rect 139616 201175 139852 201411
rect 139936 201175 140172 201411
rect 140256 201175 140492 201411
rect 140576 201175 140812 201411
rect 140896 201175 141132 201411
rect 141216 201175 141452 201411
rect 141536 201175 141772 201411
rect 141856 201175 142092 201411
rect 142176 201175 142412 201411
rect 142496 201175 142732 201411
rect 142816 201175 143052 201411
rect 143136 201175 143372 201411
rect 143456 201175 143692 201411
rect 143776 201175 144012 201411
rect 144096 201175 144332 201411
rect 144416 201175 144652 201411
rect 144736 201175 144972 201411
rect 145056 201175 145292 201411
rect 145376 201175 145612 201411
rect 145696 201175 145932 201411
rect 146016 201175 146252 201411
rect 146336 201175 146572 201411
rect 146656 201175 146892 201411
rect 146976 201175 147212 201411
rect 147296 201175 147532 201411
rect 147616 201175 147852 201411
rect 147936 201175 148172 201411
rect 148256 201175 148492 201411
rect 148576 201175 148812 201411
rect 148896 201175 149132 201411
rect 149216 201175 149452 201411
rect 149536 201175 149772 201411
rect 149856 201175 150092 201411
rect 150176 201175 150412 201411
rect 150496 201175 150732 201411
rect 150816 201175 151052 201411
rect 151136 201175 151372 201411
rect 151456 201175 151692 201411
rect 151776 201175 152012 201411
rect 152096 201175 152332 201411
rect 152416 201175 152652 201411
rect 152736 201175 152972 201411
rect 153056 201175 153292 201411
rect 153376 201175 153612 201411
rect 153696 201175 153932 201411
rect 154016 201175 154252 201411
rect 154336 201175 154572 201411
rect 154656 201175 154892 201411
rect 154976 201175 155212 201411
rect 155296 201175 155532 201411
rect 155616 201175 155852 201411
rect 155936 201175 156172 201411
rect 156256 201175 156492 201411
rect 156576 201175 156812 201411
rect 156896 201175 157132 201411
rect 157216 201175 157452 201411
rect 157536 201175 157772 201411
rect 157856 201175 158092 201411
rect 158176 201175 158412 201411
rect 158496 201175 158732 201411
rect 158816 201175 159052 201411
rect 159136 201175 159372 201411
rect 159456 201175 159692 201411
rect 159776 201175 160012 201411
rect 160096 201175 160332 201411
rect 160416 201175 160652 201411
rect 160736 201175 160972 201411
rect 161056 201175 161292 201411
rect 161376 201175 161612 201411
rect 161696 201175 161932 201411
rect 162016 201175 162252 201411
rect 162336 201175 162572 201411
rect 162656 201175 162892 201411
rect 162976 201175 163212 201411
rect 163296 201175 163532 201411
rect 163616 201175 163852 201411
rect 163936 201175 164172 201411
rect 164256 201175 164492 201411
rect 164576 201175 164812 201411
rect 164896 201175 165132 201411
rect 165216 201175 165452 201411
rect 137066 174218 137302 174454
rect 137386 174218 137622 174454
rect 137706 174218 137942 174454
rect 138026 174218 138262 174454
rect 138346 174218 138582 174454
rect 138666 174218 138902 174454
rect 138986 174218 139222 174454
rect 139306 174218 139542 174454
rect 139626 174218 139862 174454
rect 139946 174218 140182 174454
rect 140266 174218 140502 174454
rect 140586 174218 140822 174454
rect 140906 174218 141142 174454
rect 141226 174218 141462 174454
rect 137066 173898 137302 174134
rect 137386 173898 137622 174134
rect 137706 173898 137942 174134
rect 138026 173898 138262 174134
rect 138346 173898 138582 174134
rect 138666 173898 138902 174134
rect 138986 173898 139222 174134
rect 139306 173898 139542 174134
rect 139626 173898 139862 174134
rect 139946 173898 140182 174134
rect 140266 173898 140502 174134
rect 140586 173898 140822 174134
rect 140906 173898 141142 174134
rect 141226 173898 141462 174134
rect 132326 169718 132562 169954
rect 132646 169718 132882 169954
rect 132326 169398 132562 169634
rect 132646 169398 132882 169634
rect 172826 174218 173062 174454
rect 173146 174218 173382 174454
rect 172826 173898 173062 174134
rect 173146 173898 173382 174134
rect 177326 214718 177562 214954
rect 177646 214718 177882 214954
rect 177326 214398 177562 214634
rect 177646 214398 177882 214634
rect 177326 178718 177562 178954
rect 177646 178718 177882 178954
rect 177326 178398 177562 178634
rect 177646 178398 177882 178634
rect 177326 142718 177562 142954
rect 177646 142718 177882 142954
rect 177326 142398 177562 142634
rect 177646 142398 177882 142634
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 186326 223718 186562 223954
rect 186646 223718 186882 223954
rect 186326 223398 186562 223634
rect 186646 223398 186882 223634
rect 186326 187718 186562 187954
rect 186646 187718 186882 187954
rect 186326 187398 186562 187634
rect 186646 187398 186882 187634
rect 186326 151718 186562 151954
rect 186646 151718 186882 151954
rect 186326 151398 186562 151634
rect 186646 151398 186882 151634
rect 114326 115718 114562 115954
rect 114646 115718 114882 115954
rect 114326 115398 114562 115634
rect 114646 115398 114882 115634
rect 139610 115718 139846 115954
rect 139610 115398 139846 115634
rect 170330 115718 170566 115954
rect 170330 115398 170566 115634
rect 186326 115718 186562 115954
rect 186646 115718 186882 115954
rect 186326 115398 186562 115634
rect 186646 115398 186882 115634
rect 124250 111218 124486 111454
rect 124250 110898 124486 111134
rect 154970 111218 155206 111454
rect 154970 110898 155206 111134
rect 114326 79718 114562 79954
rect 114646 79718 114882 79954
rect 114326 79398 114562 79634
rect 114646 79398 114882 79634
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1542 114562 -1306
rect 114646 -1542 114882 -1306
rect 114326 -1862 114562 -1626
rect 114646 -1862 114882 -1626
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2502 119062 -2266
rect 119146 -2502 119382 -2266
rect 118826 -2822 119062 -2586
rect 119146 -2822 119382 -2586
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 123326 -3462 123562 -3226
rect 123646 -3462 123882 -3226
rect 123326 -3782 123562 -3546
rect 123646 -3782 123882 -3546
rect 132326 61718 132562 61954
rect 132646 61718 132882 61954
rect 132326 61398 132562 61634
rect 132646 61398 132882 61634
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 127826 -4422 128062 -4186
rect 128146 -4422 128382 -4186
rect 127826 -4742 128062 -4506
rect 128146 -4742 128382 -4506
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 132326 -5382 132562 -5146
rect 132646 -5382 132882 -5146
rect 132326 -5702 132562 -5466
rect 132646 -5702 132882 -5466
rect 141326 70718 141562 70954
rect 141646 70718 141882 70954
rect 141326 70398 141562 70634
rect 141646 70398 141882 70634
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 136826 -6342 137062 -6106
rect 137146 -6342 137382 -6106
rect 136826 -6662 137062 -6426
rect 137146 -6662 137382 -6426
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 141326 -7302 141562 -7066
rect 141646 -7302 141882 -7066
rect 141326 -7622 141562 -7386
rect 141646 -7622 141882 -7386
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 150326 -1542 150562 -1306
rect 150646 -1542 150882 -1306
rect 150326 -1862 150562 -1626
rect 150646 -1862 150882 -1626
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 154826 -2502 155062 -2266
rect 155146 -2502 155382 -2266
rect 154826 -2822 155062 -2586
rect 155146 -2822 155382 -2586
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 159326 -3462 159562 -3226
rect 159646 -3462 159882 -3226
rect 159326 -3782 159562 -3546
rect 159646 -3782 159882 -3546
rect 168326 61718 168562 61954
rect 168646 61718 168882 61954
rect 168326 61398 168562 61634
rect 168646 61398 168882 61634
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 163826 -4422 164062 -4186
rect 164146 -4422 164382 -4186
rect 163826 -4742 164062 -4506
rect 164146 -4742 164382 -4506
rect 186326 79718 186562 79954
rect 186646 79718 186882 79954
rect 186326 79398 186562 79634
rect 186646 79398 186882 79634
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 168326 -5382 168562 -5146
rect 168646 -5382 168882 -5146
rect 168326 -5702 168562 -5466
rect 168646 -5702 168882 -5466
rect 172826 -6342 173062 -6106
rect 173146 -6342 173382 -6106
rect 172826 -6662 173062 -6426
rect 173146 -6662 173382 -6426
rect 177326 70718 177562 70954
rect 177646 70718 177882 70954
rect 177326 70398 177562 70634
rect 177646 70398 177882 70634
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 177326 -7302 177562 -7066
rect 177646 -7302 177882 -7066
rect 177326 -7622 177562 -7386
rect 177646 -7622 177882 -7386
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1542 186562 -1306
rect 186646 -1542 186882 -1306
rect 186326 -1862 186562 -1626
rect 186646 -1862 186882 -1626
rect 190826 228217 191062 228453
rect 191146 228217 191382 228453
rect 190826 227897 191062 228133
rect 191146 227897 191382 228133
rect 190826 192218 191062 192454
rect 191146 192218 191382 192454
rect 190826 191898 191062 192134
rect 191146 191898 191382 192134
rect 190826 156218 191062 156454
rect 191146 156218 191382 156454
rect 190826 155898 191062 156134
rect 191146 155898 191382 156134
rect 190826 120218 191062 120454
rect 191146 120218 191382 120454
rect 190826 119898 191062 120134
rect 191146 119898 191382 120134
rect 190826 84218 191062 84454
rect 191146 84218 191382 84454
rect 190826 83898 191062 84134
rect 191146 83898 191382 84134
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2502 191062 -2266
rect 191146 -2502 191382 -2266
rect 190826 -2822 191062 -2586
rect 191146 -2822 191382 -2586
rect 195326 196718 195562 196954
rect 195646 196718 195882 196954
rect 195326 196398 195562 196634
rect 195646 196398 195882 196634
rect 195326 160718 195562 160954
rect 195646 160718 195882 160954
rect 195326 160398 195562 160634
rect 195646 160398 195882 160634
rect 195326 124718 195562 124954
rect 195646 124718 195882 124954
rect 195326 124398 195562 124634
rect 195646 124398 195882 124634
rect 195326 88718 195562 88954
rect 195646 88718 195882 88954
rect 195326 88398 195562 88634
rect 195646 88398 195882 88634
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3462 195562 -3226
rect 195646 -3462 195882 -3226
rect 195326 -3782 195562 -3546
rect 195646 -3782 195882 -3546
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4422 200062 -4186
rect 200146 -4422 200382 -4186
rect 199826 -4742 200062 -4506
rect 200146 -4742 200382 -4506
rect 204326 205718 204562 205954
rect 204646 205718 204882 205954
rect 204326 205398 204562 205634
rect 204646 205398 204882 205634
rect 204326 169718 204562 169954
rect 204646 169718 204882 169954
rect 204326 169398 204562 169634
rect 204646 169398 204882 169634
rect 204326 133718 204562 133954
rect 204646 133718 204882 133954
rect 204326 133398 204562 133634
rect 204646 133398 204882 133634
rect 204326 97718 204562 97954
rect 204646 97718 204882 97954
rect 204326 97398 204562 97634
rect 204646 97398 204882 97634
rect 204326 61718 204562 61954
rect 204646 61718 204882 61954
rect 204326 61398 204562 61634
rect 204646 61398 204882 61634
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 204326 -5382 204562 -5146
rect 204646 -5382 204882 -5146
rect 204326 -5702 204562 -5466
rect 204646 -5702 204882 -5466
rect 208826 210218 209062 210454
rect 209146 210218 209382 210454
rect 208826 209898 209062 210134
rect 209146 209898 209382 210134
rect 208826 174218 209062 174454
rect 209146 174218 209382 174454
rect 208826 173898 209062 174134
rect 209146 173898 209382 174134
rect 208826 138218 209062 138454
rect 209146 138218 209382 138454
rect 208826 137898 209062 138134
rect 209146 137898 209382 138134
rect 208826 102218 209062 102454
rect 209146 102218 209382 102454
rect 208826 101898 209062 102134
rect 209146 101898 209382 102134
rect 208826 66218 209062 66454
rect 209146 66218 209382 66454
rect 208826 65898 209062 66134
rect 209146 65898 209382 66134
rect 208826 30218 209062 30454
rect 209146 30218 209382 30454
rect 208826 29898 209062 30134
rect 209146 29898 209382 30134
rect 208826 -6342 209062 -6106
rect 209146 -6342 209382 -6106
rect 208826 -6662 209062 -6426
rect 209146 -6662 209382 -6426
rect 213326 214718 213562 214954
rect 213646 214718 213882 214954
rect 213326 214398 213562 214634
rect 213646 214398 213882 214634
rect 213326 178718 213562 178954
rect 213646 178718 213882 178954
rect 213326 178398 213562 178634
rect 213646 178398 213882 178634
rect 213326 142718 213562 142954
rect 213646 142718 213882 142954
rect 213326 142398 213562 142634
rect 213646 142398 213882 142634
rect 213326 106718 213562 106954
rect 213646 106718 213882 106954
rect 213326 106398 213562 106634
rect 213646 106398 213882 106634
rect 213326 70718 213562 70954
rect 213646 70718 213882 70954
rect 213326 70398 213562 70634
rect 213646 70398 213882 70634
rect 213326 34718 213562 34954
rect 213646 34718 213882 34954
rect 213326 34398 213562 34634
rect 213646 34398 213882 34634
rect 213326 -7302 213562 -7066
rect 213646 -7302 213882 -7066
rect 213326 -7622 213562 -7386
rect 213646 -7622 213882 -7386
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 222326 223718 222562 223954
rect 222646 223718 222882 223954
rect 222326 223398 222562 223634
rect 222646 223398 222882 223634
rect 222326 187718 222562 187954
rect 222646 187718 222882 187954
rect 222326 187398 222562 187634
rect 222646 187398 222882 187634
rect 222326 151718 222562 151954
rect 222646 151718 222882 151954
rect 222326 151398 222562 151634
rect 222646 151398 222882 151634
rect 222326 115718 222562 115954
rect 222646 115718 222882 115954
rect 222326 115398 222562 115634
rect 222646 115398 222882 115634
rect 222326 79718 222562 79954
rect 222646 79718 222882 79954
rect 222326 79398 222562 79634
rect 222646 79398 222882 79634
rect 222326 43718 222562 43954
rect 222646 43718 222882 43954
rect 222326 43398 222562 43634
rect 222646 43398 222882 43634
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 222326 -1542 222562 -1306
rect 222646 -1542 222882 -1306
rect 222326 -1862 222562 -1626
rect 222646 -1862 222882 -1626
rect 226826 228217 227062 228453
rect 227146 228217 227382 228453
rect 226826 227897 227062 228133
rect 227146 227897 227382 228133
rect 226826 192218 227062 192454
rect 227146 192218 227382 192454
rect 226826 191898 227062 192134
rect 227146 191898 227382 192134
rect 226826 156218 227062 156454
rect 227146 156218 227382 156454
rect 226826 155898 227062 156134
rect 227146 155898 227382 156134
rect 226826 120218 227062 120454
rect 227146 120218 227382 120454
rect 226826 119898 227062 120134
rect 227146 119898 227382 120134
rect 226826 84218 227062 84454
rect 227146 84218 227382 84454
rect 226826 83898 227062 84134
rect 227146 83898 227382 84134
rect 226826 48218 227062 48454
rect 227146 48218 227382 48454
rect 226826 47898 227062 48134
rect 227146 47898 227382 48134
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2502 227062 -2266
rect 227146 -2502 227382 -2266
rect 226826 -2822 227062 -2586
rect 227146 -2822 227382 -2586
rect 231326 196718 231562 196954
rect 231646 196718 231882 196954
rect 231326 196398 231562 196634
rect 231646 196398 231882 196634
rect 231326 160718 231562 160954
rect 231646 160718 231882 160954
rect 231326 160398 231562 160634
rect 231646 160398 231882 160634
rect 231326 124718 231562 124954
rect 231646 124718 231882 124954
rect 231326 124398 231562 124634
rect 231646 124398 231882 124634
rect 231326 88718 231562 88954
rect 231646 88718 231882 88954
rect 231326 88398 231562 88634
rect 231646 88398 231882 88634
rect 231326 52718 231562 52954
rect 231646 52718 231882 52954
rect 231326 52398 231562 52634
rect 231646 52398 231882 52634
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3462 231562 -3226
rect 231646 -3462 231882 -3226
rect 231326 -3782 231562 -3546
rect 231646 -3782 231882 -3546
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4422 236062 -4186
rect 236146 -4422 236382 -4186
rect 235826 -4742 236062 -4506
rect 236146 -4742 236382 -4506
rect 240326 205718 240562 205954
rect 240646 205718 240882 205954
rect 240326 205398 240562 205634
rect 240646 205398 240882 205634
rect 240326 169718 240562 169954
rect 240646 169718 240882 169954
rect 240326 169398 240562 169634
rect 240646 169398 240882 169634
rect 240326 133718 240562 133954
rect 240646 133718 240882 133954
rect 240326 133398 240562 133634
rect 240646 133398 240882 133634
rect 240326 97718 240562 97954
rect 240646 97718 240882 97954
rect 240326 97398 240562 97634
rect 240646 97398 240882 97634
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 240326 -5382 240562 -5146
rect 240646 -5382 240882 -5146
rect 240326 -5702 240562 -5466
rect 240646 -5702 240882 -5466
rect 244826 210218 245062 210454
rect 245146 210218 245382 210454
rect 244826 209898 245062 210134
rect 245146 209898 245382 210134
rect 244826 174218 245062 174454
rect 245146 174218 245382 174454
rect 244826 173898 245062 174134
rect 245146 173898 245382 174134
rect 244826 138218 245062 138454
rect 245146 138218 245382 138454
rect 244826 137898 245062 138134
rect 245146 137898 245382 138134
rect 244826 102218 245062 102454
rect 245146 102218 245382 102454
rect 244826 101898 245062 102134
rect 245146 101898 245382 102134
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 244826 30218 245062 30454
rect 245146 30218 245382 30454
rect 244826 29898 245062 30134
rect 245146 29898 245382 30134
rect 244826 -6342 245062 -6106
rect 245146 -6342 245382 -6106
rect 244826 -6662 245062 -6426
rect 245146 -6662 245382 -6426
rect 249326 214718 249562 214954
rect 249646 214718 249882 214954
rect 249326 214398 249562 214634
rect 249646 214398 249882 214634
rect 249326 178718 249562 178954
rect 249646 178718 249882 178954
rect 249326 178398 249562 178634
rect 249646 178398 249882 178634
rect 249326 142718 249562 142954
rect 249646 142718 249882 142954
rect 249326 142398 249562 142634
rect 249646 142398 249882 142634
rect 249326 106718 249562 106954
rect 249646 106718 249882 106954
rect 249326 106398 249562 106634
rect 249646 106398 249882 106634
rect 249326 70718 249562 70954
rect 249646 70718 249882 70954
rect 249326 70398 249562 70634
rect 249646 70398 249882 70634
rect 249326 34718 249562 34954
rect 249646 34718 249882 34954
rect 249326 34398 249562 34634
rect 249646 34398 249882 34634
rect 249326 -7302 249562 -7066
rect 249646 -7302 249882 -7066
rect 249326 -7622 249562 -7386
rect 249646 -7622 249882 -7386
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 258326 223718 258562 223954
rect 258646 223718 258882 223954
rect 258326 223398 258562 223634
rect 258646 223398 258882 223634
rect 258326 187718 258562 187954
rect 258646 187718 258882 187954
rect 258326 187398 258562 187634
rect 258646 187398 258882 187634
rect 258326 151718 258562 151954
rect 258646 151718 258882 151954
rect 258326 151398 258562 151634
rect 258646 151398 258882 151634
rect 258326 115718 258562 115954
rect 258646 115718 258882 115954
rect 258326 115398 258562 115634
rect 258646 115398 258882 115634
rect 258326 79718 258562 79954
rect 258646 79718 258882 79954
rect 258326 79398 258562 79634
rect 258646 79398 258882 79634
rect 258326 43718 258562 43954
rect 258646 43718 258882 43954
rect 258326 43398 258562 43634
rect 258646 43398 258882 43634
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 258326 -1542 258562 -1306
rect 258646 -1542 258882 -1306
rect 258326 -1862 258562 -1626
rect 258646 -1862 258882 -1626
rect 262826 228217 263062 228453
rect 263146 228217 263382 228453
rect 262826 227897 263062 228133
rect 263146 227897 263382 228133
rect 262826 192218 263062 192454
rect 263146 192218 263382 192454
rect 262826 191898 263062 192134
rect 263146 191898 263382 192134
rect 262826 156218 263062 156454
rect 263146 156218 263382 156454
rect 262826 155898 263062 156134
rect 263146 155898 263382 156134
rect 262826 120218 263062 120454
rect 263146 120218 263382 120454
rect 262826 119898 263062 120134
rect 263146 119898 263382 120134
rect 262826 84218 263062 84454
rect 263146 84218 263382 84454
rect 262826 83898 263062 84134
rect 263146 83898 263382 84134
rect 262826 48218 263062 48454
rect 263146 48218 263382 48454
rect 262826 47898 263062 48134
rect 263146 47898 263382 48134
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 262826 -2502 263062 -2266
rect 263146 -2502 263382 -2266
rect 262826 -2822 263062 -2586
rect 263146 -2822 263382 -2586
rect 267326 196718 267562 196954
rect 267646 196718 267882 196954
rect 267326 196398 267562 196634
rect 267646 196398 267882 196634
rect 267326 160718 267562 160954
rect 267646 160718 267882 160954
rect 267326 160398 267562 160634
rect 267646 160398 267882 160634
rect 267326 124718 267562 124954
rect 267646 124718 267882 124954
rect 267326 124398 267562 124634
rect 267646 124398 267882 124634
rect 267326 88718 267562 88954
rect 267646 88718 267882 88954
rect 267326 88398 267562 88634
rect 267646 88398 267882 88634
rect 267326 52718 267562 52954
rect 267646 52718 267882 52954
rect 267326 52398 267562 52634
rect 267646 52398 267882 52634
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3462 267562 -3226
rect 267646 -3462 267882 -3226
rect 267326 -3782 267562 -3546
rect 267646 -3782 267882 -3546
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4422 272062 -4186
rect 272146 -4422 272382 -4186
rect 271826 -4742 272062 -4506
rect 272146 -4742 272382 -4506
rect 276326 205718 276562 205954
rect 276646 205718 276882 205954
rect 276326 205398 276562 205634
rect 276646 205398 276882 205634
rect 276326 169718 276562 169954
rect 276646 169718 276882 169954
rect 276326 169398 276562 169634
rect 276646 169398 276882 169634
rect 276326 133718 276562 133954
rect 276646 133718 276882 133954
rect 276326 133398 276562 133634
rect 276646 133398 276882 133634
rect 276326 97718 276562 97954
rect 276646 97718 276882 97954
rect 276326 97398 276562 97634
rect 276646 97398 276882 97634
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 276326 -5382 276562 -5146
rect 276646 -5382 276882 -5146
rect 276326 -5702 276562 -5466
rect 276646 -5702 276882 -5466
rect 280826 210218 281062 210454
rect 281146 210218 281382 210454
rect 280826 209898 281062 210134
rect 281146 209898 281382 210134
rect 280826 174218 281062 174454
rect 281146 174218 281382 174454
rect 280826 173898 281062 174134
rect 281146 173898 281382 174134
rect 280826 138218 281062 138454
rect 281146 138218 281382 138454
rect 280826 137898 281062 138134
rect 281146 137898 281382 138134
rect 280826 102218 281062 102454
rect 281146 102218 281382 102454
rect 280826 101898 281062 102134
rect 281146 101898 281382 102134
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 280826 30218 281062 30454
rect 281146 30218 281382 30454
rect 280826 29898 281062 30134
rect 281146 29898 281382 30134
rect 280826 -6342 281062 -6106
rect 281146 -6342 281382 -6106
rect 280826 -6662 281062 -6426
rect 281146 -6662 281382 -6426
rect 285326 214718 285562 214954
rect 285646 214718 285882 214954
rect 285326 214398 285562 214634
rect 285646 214398 285882 214634
rect 285326 178718 285562 178954
rect 285646 178718 285882 178954
rect 285326 178398 285562 178634
rect 285646 178398 285882 178634
rect 285326 142718 285562 142954
rect 285646 142718 285882 142954
rect 285326 142398 285562 142634
rect 285646 142398 285882 142634
rect 285326 106718 285562 106954
rect 285646 106718 285882 106954
rect 285326 106398 285562 106634
rect 285646 106398 285882 106634
rect 285326 70718 285562 70954
rect 285646 70718 285882 70954
rect 285326 70398 285562 70634
rect 285646 70398 285882 70634
rect 285326 34718 285562 34954
rect 285646 34718 285882 34954
rect 285326 34398 285562 34634
rect 285646 34398 285882 34634
rect 285326 -7302 285562 -7066
rect 285646 -7302 285882 -7066
rect 285326 -7622 285562 -7386
rect 285646 -7622 285882 -7386
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 294326 223718 294562 223954
rect 294646 223718 294882 223954
rect 294326 223398 294562 223634
rect 294646 223398 294882 223634
rect 294326 187718 294562 187954
rect 294646 187718 294882 187954
rect 294326 187398 294562 187634
rect 294646 187398 294882 187634
rect 294326 151718 294562 151954
rect 294646 151718 294882 151954
rect 294326 151398 294562 151634
rect 294646 151398 294882 151634
rect 294326 115718 294562 115954
rect 294646 115718 294882 115954
rect 294326 115398 294562 115634
rect 294646 115398 294882 115634
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 294326 43718 294562 43954
rect 294646 43718 294882 43954
rect 294326 43398 294562 43634
rect 294646 43398 294882 43634
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 294326 -1542 294562 -1306
rect 294646 -1542 294882 -1306
rect 294326 -1862 294562 -1626
rect 294646 -1862 294882 -1626
rect 298826 228217 299062 228453
rect 299146 228217 299382 228453
rect 298826 227897 299062 228133
rect 299146 227897 299382 228133
rect 298826 192218 299062 192454
rect 299146 192218 299382 192454
rect 298826 191898 299062 192134
rect 299146 191898 299382 192134
rect 298826 156218 299062 156454
rect 299146 156218 299382 156454
rect 298826 155898 299062 156134
rect 299146 155898 299382 156134
rect 298826 120218 299062 120454
rect 299146 120218 299382 120454
rect 298826 119898 299062 120134
rect 299146 119898 299382 120134
rect 298826 84218 299062 84454
rect 299146 84218 299382 84454
rect 298826 83898 299062 84134
rect 299146 83898 299382 84134
rect 298826 48218 299062 48454
rect 299146 48218 299382 48454
rect 298826 47898 299062 48134
rect 299146 47898 299382 48134
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 298826 -2502 299062 -2266
rect 299146 -2502 299382 -2266
rect 298826 -2822 299062 -2586
rect 299146 -2822 299382 -2586
rect 303326 196718 303562 196954
rect 303646 196718 303882 196954
rect 303326 196398 303562 196634
rect 303646 196398 303882 196634
rect 303326 160718 303562 160954
rect 303646 160718 303882 160954
rect 303326 160398 303562 160634
rect 303646 160398 303882 160634
rect 303326 124718 303562 124954
rect 303646 124718 303882 124954
rect 303326 124398 303562 124634
rect 303646 124398 303882 124634
rect 303326 88718 303562 88954
rect 303646 88718 303882 88954
rect 303326 88398 303562 88634
rect 303646 88398 303882 88634
rect 303326 52718 303562 52954
rect 303646 52718 303882 52954
rect 303326 52398 303562 52634
rect 303646 52398 303882 52634
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 303326 -3462 303562 -3226
rect 303646 -3462 303882 -3226
rect 303326 -3782 303562 -3546
rect 303646 -3782 303882 -3546
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4422 308062 -4186
rect 308146 -4422 308382 -4186
rect 307826 -4742 308062 -4506
rect 308146 -4742 308382 -4506
rect 312326 205718 312562 205954
rect 312646 205718 312882 205954
rect 312326 205398 312562 205634
rect 312646 205398 312882 205634
rect 312326 169718 312562 169954
rect 312646 169718 312882 169954
rect 312326 169398 312562 169634
rect 312646 169398 312882 169634
rect 312326 133718 312562 133954
rect 312646 133718 312882 133954
rect 312326 133398 312562 133634
rect 312646 133398 312882 133634
rect 312326 97718 312562 97954
rect 312646 97718 312882 97954
rect 312326 97398 312562 97634
rect 312646 97398 312882 97634
rect 312326 61718 312562 61954
rect 312646 61718 312882 61954
rect 312326 61398 312562 61634
rect 312646 61398 312882 61634
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 312326 -5382 312562 -5146
rect 312646 -5382 312882 -5146
rect 312326 -5702 312562 -5466
rect 312646 -5702 312882 -5466
rect 316826 210218 317062 210454
rect 317146 210218 317382 210454
rect 316826 209898 317062 210134
rect 317146 209898 317382 210134
rect 316826 174218 317062 174454
rect 317146 174218 317382 174454
rect 316826 173898 317062 174134
rect 317146 173898 317382 174134
rect 316826 138218 317062 138454
rect 317146 138218 317382 138454
rect 316826 137898 317062 138134
rect 317146 137898 317382 138134
rect 316826 102218 317062 102454
rect 317146 102218 317382 102454
rect 316826 101898 317062 102134
rect 317146 101898 317382 102134
rect 316826 66218 317062 66454
rect 317146 66218 317382 66454
rect 316826 65898 317062 66134
rect 317146 65898 317382 66134
rect 316826 30218 317062 30454
rect 317146 30218 317382 30454
rect 316826 29898 317062 30134
rect 317146 29898 317382 30134
rect 316826 -6342 317062 -6106
rect 317146 -6342 317382 -6106
rect 316826 -6662 317062 -6426
rect 317146 -6662 317382 -6426
rect 321326 214718 321562 214954
rect 321646 214718 321882 214954
rect 321326 214398 321562 214634
rect 321646 214398 321882 214634
rect 321326 178718 321562 178954
rect 321646 178718 321882 178954
rect 321326 178398 321562 178634
rect 321646 178398 321882 178634
rect 321326 142718 321562 142954
rect 321646 142718 321882 142954
rect 321326 142398 321562 142634
rect 321646 142398 321882 142634
rect 321326 106718 321562 106954
rect 321646 106718 321882 106954
rect 321326 106398 321562 106634
rect 321646 106398 321882 106634
rect 321326 70718 321562 70954
rect 321646 70718 321882 70954
rect 321326 70398 321562 70634
rect 321646 70398 321882 70634
rect 321326 34718 321562 34954
rect 321646 34718 321882 34954
rect 321326 34398 321562 34634
rect 321646 34398 321882 34634
rect 321326 -7302 321562 -7066
rect 321646 -7302 321882 -7066
rect 321326 -7622 321562 -7386
rect 321646 -7622 321882 -7386
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 330326 223718 330562 223954
rect 330646 223718 330882 223954
rect 330326 223398 330562 223634
rect 330646 223398 330882 223634
rect 330326 187718 330562 187954
rect 330646 187718 330882 187954
rect 330326 187398 330562 187634
rect 330646 187398 330882 187634
rect 330326 151718 330562 151954
rect 330646 151718 330882 151954
rect 330326 151398 330562 151634
rect 330646 151398 330882 151634
rect 330326 115718 330562 115954
rect 330646 115718 330882 115954
rect 330326 115398 330562 115634
rect 330646 115398 330882 115634
rect 330326 79718 330562 79954
rect 330646 79718 330882 79954
rect 330326 79398 330562 79634
rect 330646 79398 330882 79634
rect 330326 43718 330562 43954
rect 330646 43718 330882 43954
rect 330326 43398 330562 43634
rect 330646 43398 330882 43634
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1542 330562 -1306
rect 330646 -1542 330882 -1306
rect 330326 -1862 330562 -1626
rect 330646 -1862 330882 -1626
rect 334826 228217 335062 228453
rect 335146 228217 335382 228453
rect 334826 227897 335062 228133
rect 335146 227897 335382 228133
rect 334826 192218 335062 192454
rect 335146 192218 335382 192454
rect 334826 191898 335062 192134
rect 335146 191898 335382 192134
rect 334826 156218 335062 156454
rect 335146 156218 335382 156454
rect 334826 155898 335062 156134
rect 335146 155898 335382 156134
rect 334826 120218 335062 120454
rect 335146 120218 335382 120454
rect 334826 119898 335062 120134
rect 335146 119898 335382 120134
rect 334826 84218 335062 84454
rect 335146 84218 335382 84454
rect 334826 83898 335062 84134
rect 335146 83898 335382 84134
rect 334826 48218 335062 48454
rect 335146 48218 335382 48454
rect 334826 47898 335062 48134
rect 335146 47898 335382 48134
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2502 335062 -2266
rect 335146 -2502 335382 -2266
rect 334826 -2822 335062 -2586
rect 335146 -2822 335382 -2586
rect 339326 196718 339562 196954
rect 339646 196718 339882 196954
rect 339326 196398 339562 196634
rect 339646 196398 339882 196634
rect 339326 160718 339562 160954
rect 339646 160718 339882 160954
rect 339326 160398 339562 160634
rect 339646 160398 339882 160634
rect 339326 124718 339562 124954
rect 339646 124718 339882 124954
rect 339326 124398 339562 124634
rect 339646 124398 339882 124634
rect 339326 88718 339562 88954
rect 339646 88718 339882 88954
rect 339326 88398 339562 88634
rect 339646 88398 339882 88634
rect 339326 52718 339562 52954
rect 339646 52718 339882 52954
rect 339326 52398 339562 52634
rect 339646 52398 339882 52634
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 339326 -3462 339562 -3226
rect 339646 -3462 339882 -3226
rect 339326 -3782 339562 -3546
rect 339646 -3782 339882 -3546
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -4422 344062 -4186
rect 344146 -4422 344382 -4186
rect 343826 -4742 344062 -4506
rect 344146 -4742 344382 -4506
rect 348326 205718 348562 205954
rect 348646 205718 348882 205954
rect 348326 205398 348562 205634
rect 348646 205398 348882 205634
rect 348326 169718 348562 169954
rect 348646 169718 348882 169954
rect 348326 169398 348562 169634
rect 348646 169398 348882 169634
rect 348326 133718 348562 133954
rect 348646 133718 348882 133954
rect 348326 133398 348562 133634
rect 348646 133398 348882 133634
rect 348326 97718 348562 97954
rect 348646 97718 348882 97954
rect 348326 97398 348562 97634
rect 348646 97398 348882 97634
rect 348326 61718 348562 61954
rect 348646 61718 348882 61954
rect 348326 61398 348562 61634
rect 348646 61398 348882 61634
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 348326 -5382 348562 -5146
rect 348646 -5382 348882 -5146
rect 348326 -5702 348562 -5466
rect 348646 -5702 348882 -5466
rect 352826 210218 353062 210454
rect 353146 210218 353382 210454
rect 352826 209898 353062 210134
rect 353146 209898 353382 210134
rect 352826 174218 353062 174454
rect 353146 174218 353382 174454
rect 352826 173898 353062 174134
rect 353146 173898 353382 174134
rect 352826 138218 353062 138454
rect 353146 138218 353382 138454
rect 352826 137898 353062 138134
rect 353146 137898 353382 138134
rect 352826 102218 353062 102454
rect 353146 102218 353382 102454
rect 352826 101898 353062 102134
rect 353146 101898 353382 102134
rect 352826 66218 353062 66454
rect 353146 66218 353382 66454
rect 352826 65898 353062 66134
rect 353146 65898 353382 66134
rect 352826 30218 353062 30454
rect 353146 30218 353382 30454
rect 352826 29898 353062 30134
rect 353146 29898 353382 30134
rect 352826 -6342 353062 -6106
rect 353146 -6342 353382 -6106
rect 352826 -6662 353062 -6426
rect 353146 -6662 353382 -6426
rect 357326 214718 357562 214954
rect 357646 214718 357882 214954
rect 357326 214398 357562 214634
rect 357646 214398 357882 214634
rect 357326 178718 357562 178954
rect 357646 178718 357882 178954
rect 357326 178398 357562 178634
rect 357646 178398 357882 178634
rect 357326 142718 357562 142954
rect 357646 142718 357882 142954
rect 357326 142398 357562 142634
rect 357646 142398 357882 142634
rect 357326 106718 357562 106954
rect 357646 106718 357882 106954
rect 357326 106398 357562 106634
rect 357646 106398 357882 106634
rect 357326 70718 357562 70954
rect 357646 70718 357882 70954
rect 357326 70398 357562 70634
rect 357646 70398 357882 70634
rect 357326 34718 357562 34954
rect 357646 34718 357882 34954
rect 357326 34398 357562 34634
rect 357646 34398 357882 34634
rect 357326 -7302 357562 -7066
rect 357646 -7302 357882 -7066
rect 357326 -7622 357562 -7386
rect 357646 -7622 357882 -7386
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 366326 223718 366562 223954
rect 366646 223718 366882 223954
rect 366326 223398 366562 223634
rect 366646 223398 366882 223634
rect 366326 187718 366562 187954
rect 366646 187718 366882 187954
rect 366326 187398 366562 187634
rect 366646 187398 366882 187634
rect 366326 151718 366562 151954
rect 366646 151718 366882 151954
rect 366326 151398 366562 151634
rect 366646 151398 366882 151634
rect 366326 115718 366562 115954
rect 366646 115718 366882 115954
rect 366326 115398 366562 115634
rect 366646 115398 366882 115634
rect 366326 79718 366562 79954
rect 366646 79718 366882 79954
rect 366326 79398 366562 79634
rect 366646 79398 366882 79634
rect 366326 43718 366562 43954
rect 366646 43718 366882 43954
rect 366326 43398 366562 43634
rect 366646 43398 366882 43634
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 366326 -1542 366562 -1306
rect 366646 -1542 366882 -1306
rect 366326 -1862 366562 -1626
rect 366646 -1862 366882 -1626
rect 370826 228217 371062 228453
rect 371146 228217 371382 228453
rect 370826 227897 371062 228133
rect 371146 227897 371382 228133
rect 370826 192218 371062 192454
rect 371146 192218 371382 192454
rect 370826 191898 371062 192134
rect 371146 191898 371382 192134
rect 370826 156218 371062 156454
rect 371146 156218 371382 156454
rect 370826 155898 371062 156134
rect 371146 155898 371382 156134
rect 370826 120218 371062 120454
rect 371146 120218 371382 120454
rect 370826 119898 371062 120134
rect 371146 119898 371382 120134
rect 370826 84218 371062 84454
rect 371146 84218 371382 84454
rect 370826 83898 371062 84134
rect 371146 83898 371382 84134
rect 370826 48218 371062 48454
rect 371146 48218 371382 48454
rect 370826 47898 371062 48134
rect 371146 47898 371382 48134
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -2502 371062 -2266
rect 371146 -2502 371382 -2266
rect 370826 -2822 371062 -2586
rect 371146 -2822 371382 -2586
rect 375326 196718 375562 196954
rect 375646 196718 375882 196954
rect 375326 196398 375562 196634
rect 375646 196398 375882 196634
rect 375326 160718 375562 160954
rect 375646 160718 375882 160954
rect 375326 160398 375562 160634
rect 375646 160398 375882 160634
rect 375326 124718 375562 124954
rect 375646 124718 375882 124954
rect 375326 124398 375562 124634
rect 375646 124398 375882 124634
rect 375326 88718 375562 88954
rect 375646 88718 375882 88954
rect 375326 88398 375562 88634
rect 375646 88398 375882 88634
rect 375326 52718 375562 52954
rect 375646 52718 375882 52954
rect 375326 52398 375562 52634
rect 375646 52398 375882 52634
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3462 375562 -3226
rect 375646 -3462 375882 -3226
rect 375326 -3782 375562 -3546
rect 375646 -3782 375882 -3546
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4422 380062 -4186
rect 380146 -4422 380382 -4186
rect 379826 -4742 380062 -4506
rect 380146 -4742 380382 -4506
rect 384326 205718 384562 205954
rect 384646 205718 384882 205954
rect 384326 205398 384562 205634
rect 384646 205398 384882 205634
rect 384326 169718 384562 169954
rect 384646 169718 384882 169954
rect 384326 169398 384562 169634
rect 384646 169398 384882 169634
rect 384326 133718 384562 133954
rect 384646 133718 384882 133954
rect 384326 133398 384562 133634
rect 384646 133398 384882 133634
rect 384326 97718 384562 97954
rect 384646 97718 384882 97954
rect 384326 97398 384562 97634
rect 384646 97398 384882 97634
rect 384326 61718 384562 61954
rect 384646 61718 384882 61954
rect 384326 61398 384562 61634
rect 384646 61398 384882 61634
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 384326 -5382 384562 -5146
rect 384646 -5382 384882 -5146
rect 384326 -5702 384562 -5466
rect 384646 -5702 384882 -5466
rect 388826 210218 389062 210454
rect 389146 210218 389382 210454
rect 388826 209898 389062 210134
rect 389146 209898 389382 210134
rect 388826 174218 389062 174454
rect 389146 174218 389382 174454
rect 388826 173898 389062 174134
rect 389146 173898 389382 174134
rect 388826 138218 389062 138454
rect 389146 138218 389382 138454
rect 388826 137898 389062 138134
rect 389146 137898 389382 138134
rect 388826 102218 389062 102454
rect 389146 102218 389382 102454
rect 388826 101898 389062 102134
rect 389146 101898 389382 102134
rect 388826 66218 389062 66454
rect 389146 66218 389382 66454
rect 388826 65898 389062 66134
rect 389146 65898 389382 66134
rect 388826 30218 389062 30454
rect 389146 30218 389382 30454
rect 388826 29898 389062 30134
rect 389146 29898 389382 30134
rect 388826 -6342 389062 -6106
rect 389146 -6342 389382 -6106
rect 388826 -6662 389062 -6426
rect 389146 -6662 389382 -6426
rect 393326 214718 393562 214954
rect 393646 214718 393882 214954
rect 393326 214398 393562 214634
rect 393646 214398 393882 214634
rect 393326 178718 393562 178954
rect 393646 178718 393882 178954
rect 393326 178398 393562 178634
rect 393646 178398 393882 178634
rect 393326 142718 393562 142954
rect 393646 142718 393882 142954
rect 393326 142398 393562 142634
rect 393646 142398 393882 142634
rect 393326 106718 393562 106954
rect 393646 106718 393882 106954
rect 393326 106398 393562 106634
rect 393646 106398 393882 106634
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 402326 705562 402562 705798
rect 402646 705562 402882 705798
rect 402326 705242 402562 705478
rect 402646 705242 402882 705478
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 402326 619718 402562 619954
rect 402646 619718 402882 619954
rect 402326 619398 402562 619634
rect 402646 619398 402882 619634
rect 402326 583718 402562 583954
rect 402646 583718 402882 583954
rect 402326 583398 402562 583634
rect 402646 583398 402882 583634
rect 402326 547718 402562 547954
rect 402646 547718 402882 547954
rect 402326 547398 402562 547634
rect 402646 547398 402882 547634
rect 402326 511718 402562 511954
rect 402646 511718 402882 511954
rect 402326 511398 402562 511634
rect 402646 511398 402882 511634
rect 402326 475718 402562 475954
rect 402646 475718 402882 475954
rect 402326 475398 402562 475634
rect 402646 475398 402882 475634
rect 402326 439718 402562 439954
rect 402646 439718 402882 439954
rect 402326 439398 402562 439634
rect 402646 439398 402882 439634
rect 402326 403718 402562 403954
rect 402646 403718 402882 403954
rect 402326 403398 402562 403634
rect 402646 403398 402882 403634
rect 402326 367718 402562 367954
rect 402646 367718 402882 367954
rect 402326 367398 402562 367634
rect 402646 367398 402882 367634
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 402326 295718 402562 295954
rect 402646 295718 402882 295954
rect 402326 295398 402562 295634
rect 402646 295398 402882 295634
rect 402326 259718 402562 259954
rect 402646 259718 402882 259954
rect 402326 259398 402562 259634
rect 402646 259398 402882 259634
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 393326 70718 393562 70954
rect 393646 70718 393882 70954
rect 393326 70398 393562 70634
rect 393646 70398 393882 70634
rect 393326 34718 393562 34954
rect 393646 34718 393882 34954
rect 393326 34398 393562 34634
rect 393646 34398 393882 34634
rect 393326 -7302 393562 -7066
rect 393646 -7302 393882 -7066
rect 393326 -7622 393562 -7386
rect 393646 -7622 393882 -7386
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 402326 223718 402562 223954
rect 402646 223718 402882 223954
rect 402326 223398 402562 223634
rect 402646 223398 402882 223634
rect 402326 187718 402562 187954
rect 402646 187718 402882 187954
rect 402326 187398 402562 187634
rect 402646 187398 402882 187634
rect 402326 151718 402562 151954
rect 402646 151718 402882 151954
rect 402326 151398 402562 151634
rect 402646 151398 402882 151634
rect 402326 115718 402562 115954
rect 402646 115718 402882 115954
rect 402326 115398 402562 115634
rect 402646 115398 402882 115634
rect 402326 79718 402562 79954
rect 402646 79718 402882 79954
rect 402326 79398 402562 79634
rect 402646 79398 402882 79634
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1542 402562 -1306
rect 402646 -1542 402882 -1306
rect 402326 -1862 402562 -1626
rect 402646 -1862 402882 -1626
rect 406826 706522 407062 706758
rect 407146 706522 407382 706758
rect 406826 706202 407062 706438
rect 407146 706202 407382 706438
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 406826 624218 407062 624454
rect 407146 624218 407382 624454
rect 406826 623898 407062 624134
rect 407146 623898 407382 624134
rect 406826 588218 407062 588454
rect 407146 588218 407382 588454
rect 406826 587898 407062 588134
rect 407146 587898 407382 588134
rect 406826 552218 407062 552454
rect 407146 552218 407382 552454
rect 406826 551898 407062 552134
rect 407146 551898 407382 552134
rect 406826 516218 407062 516454
rect 407146 516218 407382 516454
rect 406826 515898 407062 516134
rect 407146 515898 407382 516134
rect 406826 480218 407062 480454
rect 407146 480218 407382 480454
rect 406826 479898 407062 480134
rect 407146 479898 407382 480134
rect 406826 444218 407062 444454
rect 407146 444218 407382 444454
rect 406826 443898 407062 444134
rect 407146 443898 407382 444134
rect 406826 408218 407062 408454
rect 407146 408218 407382 408454
rect 406826 407898 407062 408134
rect 407146 407898 407382 408134
rect 406826 372218 407062 372454
rect 407146 372218 407382 372454
rect 406826 371898 407062 372134
rect 407146 371898 407382 372134
rect 406826 336218 407062 336454
rect 407146 336218 407382 336454
rect 406826 335898 407062 336134
rect 407146 335898 407382 336134
rect 406826 300218 407062 300454
rect 407146 300218 407382 300454
rect 406826 299898 407062 300134
rect 407146 299898 407382 300134
rect 406826 264218 407062 264454
rect 407146 264218 407382 264454
rect 406826 263898 407062 264134
rect 407146 263898 407382 264134
rect 406826 228218 407062 228454
rect 407146 228218 407382 228454
rect 406826 227898 407062 228134
rect 407146 227898 407382 228134
rect 406826 192218 407062 192454
rect 407146 192218 407382 192454
rect 406826 191898 407062 192134
rect 407146 191898 407382 192134
rect 406826 156218 407062 156454
rect 407146 156218 407382 156454
rect 406826 155898 407062 156134
rect 407146 155898 407382 156134
rect 406826 120218 407062 120454
rect 407146 120218 407382 120454
rect 406826 119898 407062 120134
rect 407146 119898 407382 120134
rect 406826 84218 407062 84454
rect 407146 84218 407382 84454
rect 406826 83898 407062 84134
rect 407146 83898 407382 84134
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2502 407062 -2266
rect 407146 -2502 407382 -2266
rect 406826 -2822 407062 -2586
rect 407146 -2822 407382 -2586
rect 411326 707482 411562 707718
rect 411646 707482 411882 707718
rect 411326 707162 411562 707398
rect 411646 707162 411882 707398
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 411326 664718 411562 664954
rect 411646 664718 411882 664954
rect 411326 664398 411562 664634
rect 411646 664398 411882 664634
rect 411326 628718 411562 628954
rect 411646 628718 411882 628954
rect 411326 628398 411562 628634
rect 411646 628398 411882 628634
rect 411326 592718 411562 592954
rect 411646 592718 411882 592954
rect 411326 592398 411562 592634
rect 411646 592398 411882 592634
rect 411326 556718 411562 556954
rect 411646 556718 411882 556954
rect 411326 556398 411562 556634
rect 411646 556398 411882 556634
rect 411326 520718 411562 520954
rect 411646 520718 411882 520954
rect 411326 520398 411562 520634
rect 411646 520398 411882 520634
rect 411326 484718 411562 484954
rect 411646 484718 411882 484954
rect 411326 484398 411562 484634
rect 411646 484398 411882 484634
rect 411326 448718 411562 448954
rect 411646 448718 411882 448954
rect 411326 448398 411562 448634
rect 411646 448398 411882 448634
rect 411326 412718 411562 412954
rect 411646 412718 411882 412954
rect 411326 412398 411562 412634
rect 411646 412398 411882 412634
rect 411326 376718 411562 376954
rect 411646 376718 411882 376954
rect 411326 376398 411562 376634
rect 411646 376398 411882 376634
rect 411326 340718 411562 340954
rect 411646 340718 411882 340954
rect 411326 340398 411562 340634
rect 411646 340398 411882 340634
rect 411326 304718 411562 304954
rect 411646 304718 411882 304954
rect 411326 304398 411562 304634
rect 411646 304398 411882 304634
rect 411326 268718 411562 268954
rect 411646 268718 411882 268954
rect 411326 268398 411562 268634
rect 411646 268398 411882 268634
rect 411326 232718 411562 232954
rect 411646 232718 411882 232954
rect 411326 232398 411562 232634
rect 411646 232398 411882 232634
rect 411326 196718 411562 196954
rect 411646 196718 411882 196954
rect 411326 196398 411562 196634
rect 411646 196398 411882 196634
rect 411326 160718 411562 160954
rect 411646 160718 411882 160954
rect 411326 160398 411562 160634
rect 411646 160398 411882 160634
rect 411326 124718 411562 124954
rect 411646 124718 411882 124954
rect 411326 124398 411562 124634
rect 411646 124398 411882 124634
rect 411326 88718 411562 88954
rect 411646 88718 411882 88954
rect 411326 88398 411562 88634
rect 411646 88398 411882 88634
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3462 411562 -3226
rect 411646 -3462 411882 -3226
rect 411326 -3782 411562 -3546
rect 411646 -3782 411882 -3546
rect 415826 708442 416062 708678
rect 416146 708442 416382 708678
rect 415826 708122 416062 708358
rect 416146 708122 416382 708358
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4422 416062 -4186
rect 416146 -4422 416382 -4186
rect 415826 -4742 416062 -4506
rect 416146 -4742 416382 -4506
rect 420326 709402 420562 709638
rect 420646 709402 420882 709638
rect 420326 709082 420562 709318
rect 420646 709082 420882 709318
rect 420326 673718 420562 673954
rect 420646 673718 420882 673954
rect 420326 673398 420562 673634
rect 420646 673398 420882 673634
rect 420326 637718 420562 637954
rect 420646 637718 420882 637954
rect 420326 637398 420562 637634
rect 420646 637398 420882 637634
rect 420326 601718 420562 601954
rect 420646 601718 420882 601954
rect 420326 601398 420562 601634
rect 420646 601398 420882 601634
rect 420326 565718 420562 565954
rect 420646 565718 420882 565954
rect 420326 565398 420562 565634
rect 420646 565398 420882 565634
rect 420326 529718 420562 529954
rect 420646 529718 420882 529954
rect 420326 529398 420562 529634
rect 420646 529398 420882 529634
rect 420326 493718 420562 493954
rect 420646 493718 420882 493954
rect 420326 493398 420562 493634
rect 420646 493398 420882 493634
rect 420326 457718 420562 457954
rect 420646 457718 420882 457954
rect 420326 457398 420562 457634
rect 420646 457398 420882 457634
rect 420326 421718 420562 421954
rect 420646 421718 420882 421954
rect 420326 421398 420562 421634
rect 420646 421398 420882 421634
rect 420326 385718 420562 385954
rect 420646 385718 420882 385954
rect 420326 385398 420562 385634
rect 420646 385398 420882 385634
rect 420326 349718 420562 349954
rect 420646 349718 420882 349954
rect 420326 349398 420562 349634
rect 420646 349398 420882 349634
rect 420326 313718 420562 313954
rect 420646 313718 420882 313954
rect 420326 313398 420562 313634
rect 420646 313398 420882 313634
rect 420326 277718 420562 277954
rect 420646 277718 420882 277954
rect 420326 277398 420562 277634
rect 420646 277398 420882 277634
rect 420326 241718 420562 241954
rect 420646 241718 420882 241954
rect 420326 241398 420562 241634
rect 420646 241398 420882 241634
rect 420326 205718 420562 205954
rect 420646 205718 420882 205954
rect 420326 205398 420562 205634
rect 420646 205398 420882 205634
rect 420326 169718 420562 169954
rect 420646 169718 420882 169954
rect 420326 169398 420562 169634
rect 420646 169398 420882 169634
rect 420326 133718 420562 133954
rect 420646 133718 420882 133954
rect 420326 133398 420562 133634
rect 420646 133398 420882 133634
rect 420326 97718 420562 97954
rect 420646 97718 420882 97954
rect 420326 97398 420562 97634
rect 420646 97398 420882 97634
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5382 420562 -5146
rect 420646 -5382 420882 -5146
rect 420326 -5702 420562 -5466
rect 420646 -5702 420882 -5466
rect 424826 710362 425062 710598
rect 425146 710362 425382 710598
rect 424826 710042 425062 710278
rect 425146 710042 425382 710278
rect 424826 678218 425062 678454
rect 425146 678218 425382 678454
rect 424826 677898 425062 678134
rect 425146 677898 425382 678134
rect 424826 642218 425062 642454
rect 425146 642218 425382 642454
rect 424826 641898 425062 642134
rect 425146 641898 425382 642134
rect 424826 606218 425062 606454
rect 425146 606218 425382 606454
rect 424826 605898 425062 606134
rect 425146 605898 425382 606134
rect 424826 570218 425062 570454
rect 425146 570218 425382 570454
rect 424826 569898 425062 570134
rect 425146 569898 425382 570134
rect 424826 534218 425062 534454
rect 425146 534218 425382 534454
rect 424826 533898 425062 534134
rect 425146 533898 425382 534134
rect 424826 498218 425062 498454
rect 425146 498218 425382 498454
rect 424826 497898 425062 498134
rect 425146 497898 425382 498134
rect 424826 462218 425062 462454
rect 425146 462218 425382 462454
rect 424826 461898 425062 462134
rect 425146 461898 425382 462134
rect 424826 426218 425062 426454
rect 425146 426218 425382 426454
rect 424826 425898 425062 426134
rect 425146 425898 425382 426134
rect 424826 390218 425062 390454
rect 425146 390218 425382 390454
rect 424826 389898 425062 390134
rect 425146 389898 425382 390134
rect 424826 354218 425062 354454
rect 425146 354218 425382 354454
rect 424826 353898 425062 354134
rect 425146 353898 425382 354134
rect 424826 318218 425062 318454
rect 425146 318218 425382 318454
rect 424826 317898 425062 318134
rect 425146 317898 425382 318134
rect 424826 282218 425062 282454
rect 425146 282218 425382 282454
rect 424826 281898 425062 282134
rect 425146 281898 425382 282134
rect 424826 246218 425062 246454
rect 425146 246218 425382 246454
rect 424826 245898 425062 246134
rect 425146 245898 425382 246134
rect 424826 210218 425062 210454
rect 425146 210218 425382 210454
rect 424826 209898 425062 210134
rect 425146 209898 425382 210134
rect 424826 174218 425062 174454
rect 425146 174218 425382 174454
rect 424826 173898 425062 174134
rect 425146 173898 425382 174134
rect 424826 138218 425062 138454
rect 425146 138218 425382 138454
rect 424826 137898 425062 138134
rect 425146 137898 425382 138134
rect 424826 102218 425062 102454
rect 425146 102218 425382 102454
rect 424826 101898 425062 102134
rect 425146 101898 425382 102134
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6342 425062 -6106
rect 425146 -6342 425382 -6106
rect 424826 -6662 425062 -6426
rect 425146 -6662 425382 -6426
rect 429326 711322 429562 711558
rect 429646 711322 429882 711558
rect 429326 711002 429562 711238
rect 429646 711002 429882 711238
rect 429326 682718 429562 682954
rect 429646 682718 429882 682954
rect 429326 682398 429562 682634
rect 429646 682398 429882 682634
rect 429326 646718 429562 646954
rect 429646 646718 429882 646954
rect 429326 646398 429562 646634
rect 429646 646398 429882 646634
rect 429326 610718 429562 610954
rect 429646 610718 429882 610954
rect 429326 610398 429562 610634
rect 429646 610398 429882 610634
rect 429326 574718 429562 574954
rect 429646 574718 429882 574954
rect 429326 574398 429562 574634
rect 429646 574398 429882 574634
rect 429326 538718 429562 538954
rect 429646 538718 429882 538954
rect 429326 538398 429562 538634
rect 429646 538398 429882 538634
rect 429326 502718 429562 502954
rect 429646 502718 429882 502954
rect 429326 502398 429562 502634
rect 429646 502398 429882 502634
rect 429326 466718 429562 466954
rect 429646 466718 429882 466954
rect 429326 466398 429562 466634
rect 429646 466398 429882 466634
rect 429326 430718 429562 430954
rect 429646 430718 429882 430954
rect 429326 430398 429562 430634
rect 429646 430398 429882 430634
rect 429326 394718 429562 394954
rect 429646 394718 429882 394954
rect 429326 394398 429562 394634
rect 429646 394398 429882 394634
rect 429326 358718 429562 358954
rect 429646 358718 429882 358954
rect 429326 358398 429562 358634
rect 429646 358398 429882 358634
rect 429326 322718 429562 322954
rect 429646 322718 429882 322954
rect 429326 322398 429562 322634
rect 429646 322398 429882 322634
rect 429326 286718 429562 286954
rect 429646 286718 429882 286954
rect 429326 286398 429562 286634
rect 429646 286398 429882 286634
rect 429326 250718 429562 250954
rect 429646 250718 429882 250954
rect 429326 250398 429562 250634
rect 429646 250398 429882 250634
rect 429326 214718 429562 214954
rect 429646 214718 429882 214954
rect 429326 214398 429562 214634
rect 429646 214398 429882 214634
rect 429326 178718 429562 178954
rect 429646 178718 429882 178954
rect 429326 178398 429562 178634
rect 429646 178398 429882 178634
rect 429326 142718 429562 142954
rect 429646 142718 429882 142954
rect 429326 142398 429562 142634
rect 429646 142398 429882 142634
rect 429326 106718 429562 106954
rect 429646 106718 429882 106954
rect 429326 106398 429562 106634
rect 429646 106398 429882 106634
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7302 429562 -7066
rect 429646 -7302 429882 -7066
rect 429326 -7622 429562 -7386
rect 429646 -7622 429882 -7386
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 438326 705562 438562 705798
rect 438646 705562 438882 705798
rect 438326 705242 438562 705478
rect 438646 705242 438882 705478
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 438326 655718 438562 655954
rect 438646 655718 438882 655954
rect 438326 655398 438562 655634
rect 438646 655398 438882 655634
rect 438326 619718 438562 619954
rect 438646 619718 438882 619954
rect 438326 619398 438562 619634
rect 438646 619398 438882 619634
rect 438326 583718 438562 583954
rect 438646 583718 438882 583954
rect 438326 583398 438562 583634
rect 438646 583398 438882 583634
rect 438326 547718 438562 547954
rect 438646 547718 438882 547954
rect 438326 547398 438562 547634
rect 438646 547398 438882 547634
rect 438326 511718 438562 511954
rect 438646 511718 438882 511954
rect 438326 511398 438562 511634
rect 438646 511398 438882 511634
rect 438326 475718 438562 475954
rect 438646 475718 438882 475954
rect 438326 475398 438562 475634
rect 438646 475398 438882 475634
rect 438326 439718 438562 439954
rect 438646 439718 438882 439954
rect 438326 439398 438562 439634
rect 438646 439398 438882 439634
rect 438326 403718 438562 403954
rect 438646 403718 438882 403954
rect 438326 403398 438562 403634
rect 438646 403398 438882 403634
rect 438326 367718 438562 367954
rect 438646 367718 438882 367954
rect 438326 367398 438562 367634
rect 438646 367398 438882 367634
rect 438326 331718 438562 331954
rect 438646 331718 438882 331954
rect 438326 331398 438562 331634
rect 438646 331398 438882 331634
rect 438326 295718 438562 295954
rect 438646 295718 438882 295954
rect 438326 295398 438562 295634
rect 438646 295398 438882 295634
rect 438326 259718 438562 259954
rect 438646 259718 438882 259954
rect 438326 259398 438562 259634
rect 438646 259398 438882 259634
rect 438326 223718 438562 223954
rect 438646 223718 438882 223954
rect 438326 223398 438562 223634
rect 438646 223398 438882 223634
rect 438326 187718 438562 187954
rect 438646 187718 438882 187954
rect 438326 187398 438562 187634
rect 438646 187398 438882 187634
rect 438326 151718 438562 151954
rect 438646 151718 438882 151954
rect 438326 151398 438562 151634
rect 438646 151398 438882 151634
rect 438326 115718 438562 115954
rect 438646 115718 438882 115954
rect 438326 115398 438562 115634
rect 438646 115398 438882 115634
rect 438326 79718 438562 79954
rect 438646 79718 438882 79954
rect 438326 79398 438562 79634
rect 438646 79398 438882 79634
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1542 438562 -1306
rect 438646 -1542 438882 -1306
rect 438326 -1862 438562 -1626
rect 438646 -1862 438882 -1626
rect 442826 706522 443062 706758
rect 443146 706522 443382 706758
rect 442826 706202 443062 706438
rect 443146 706202 443382 706438
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 442826 660218 443062 660454
rect 443146 660218 443382 660454
rect 442826 659898 443062 660134
rect 443146 659898 443382 660134
rect 442826 624218 443062 624454
rect 443146 624218 443382 624454
rect 442826 623898 443062 624134
rect 443146 623898 443382 624134
rect 442826 588218 443062 588454
rect 443146 588218 443382 588454
rect 442826 587898 443062 588134
rect 443146 587898 443382 588134
rect 442826 552218 443062 552454
rect 443146 552218 443382 552454
rect 442826 551898 443062 552134
rect 443146 551898 443382 552134
rect 442826 516218 443062 516454
rect 443146 516218 443382 516454
rect 442826 515898 443062 516134
rect 443146 515898 443382 516134
rect 442826 480218 443062 480454
rect 443146 480218 443382 480454
rect 442826 479898 443062 480134
rect 443146 479898 443382 480134
rect 442826 444218 443062 444454
rect 443146 444218 443382 444454
rect 442826 443898 443062 444134
rect 443146 443898 443382 444134
rect 442826 408218 443062 408454
rect 443146 408218 443382 408454
rect 442826 407898 443062 408134
rect 443146 407898 443382 408134
rect 442826 372218 443062 372454
rect 443146 372218 443382 372454
rect 442826 371898 443062 372134
rect 443146 371898 443382 372134
rect 442826 336218 443062 336454
rect 443146 336218 443382 336454
rect 442826 335898 443062 336134
rect 443146 335898 443382 336134
rect 442826 300218 443062 300454
rect 443146 300218 443382 300454
rect 442826 299898 443062 300134
rect 443146 299898 443382 300134
rect 442826 264218 443062 264454
rect 443146 264218 443382 264454
rect 442826 263898 443062 264134
rect 443146 263898 443382 264134
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 442826 192218 443062 192454
rect 443146 192218 443382 192454
rect 442826 191898 443062 192134
rect 443146 191898 443382 192134
rect 442826 156218 443062 156454
rect 443146 156218 443382 156454
rect 442826 155898 443062 156134
rect 443146 155898 443382 156134
rect 442826 120218 443062 120454
rect 443146 120218 443382 120454
rect 442826 119898 443062 120134
rect 443146 119898 443382 120134
rect 442826 84218 443062 84454
rect 443146 84218 443382 84454
rect 442826 83898 443062 84134
rect 443146 83898 443382 84134
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2502 443062 -2266
rect 443146 -2502 443382 -2266
rect 442826 -2822 443062 -2586
rect 443146 -2822 443382 -2586
rect 447326 707482 447562 707718
rect 447646 707482 447882 707718
rect 447326 707162 447562 707398
rect 447646 707162 447882 707398
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 447326 664718 447562 664954
rect 447646 664718 447882 664954
rect 447326 664398 447562 664634
rect 447646 664398 447882 664634
rect 447326 628718 447562 628954
rect 447646 628718 447882 628954
rect 447326 628398 447562 628634
rect 447646 628398 447882 628634
rect 447326 592718 447562 592954
rect 447646 592718 447882 592954
rect 447326 592398 447562 592634
rect 447646 592398 447882 592634
rect 447326 556718 447562 556954
rect 447646 556718 447882 556954
rect 447326 556398 447562 556634
rect 447646 556398 447882 556634
rect 447326 520718 447562 520954
rect 447646 520718 447882 520954
rect 447326 520398 447562 520634
rect 447646 520398 447882 520634
rect 447326 484718 447562 484954
rect 447646 484718 447882 484954
rect 447326 484398 447562 484634
rect 447646 484398 447882 484634
rect 447326 448718 447562 448954
rect 447646 448718 447882 448954
rect 447326 448398 447562 448634
rect 447646 448398 447882 448634
rect 447326 412718 447562 412954
rect 447646 412718 447882 412954
rect 447326 412398 447562 412634
rect 447646 412398 447882 412634
rect 447326 376718 447562 376954
rect 447646 376718 447882 376954
rect 447326 376398 447562 376634
rect 447646 376398 447882 376634
rect 447326 340718 447562 340954
rect 447646 340718 447882 340954
rect 447326 340398 447562 340634
rect 447646 340398 447882 340634
rect 447326 304718 447562 304954
rect 447646 304718 447882 304954
rect 447326 304398 447562 304634
rect 447646 304398 447882 304634
rect 447326 268718 447562 268954
rect 447646 268718 447882 268954
rect 447326 268398 447562 268634
rect 447646 268398 447882 268634
rect 447326 232718 447562 232954
rect 447646 232718 447882 232954
rect 447326 232398 447562 232634
rect 447646 232398 447882 232634
rect 447326 196718 447562 196954
rect 447646 196718 447882 196954
rect 447326 196398 447562 196634
rect 447646 196398 447882 196634
rect 447326 160718 447562 160954
rect 447646 160718 447882 160954
rect 447326 160398 447562 160634
rect 447646 160398 447882 160634
rect 447326 124718 447562 124954
rect 447646 124718 447882 124954
rect 447326 124398 447562 124634
rect 447646 124398 447882 124634
rect 447326 88718 447562 88954
rect 447646 88718 447882 88954
rect 447326 88398 447562 88634
rect 447646 88398 447882 88634
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3462 447562 -3226
rect 447646 -3462 447882 -3226
rect 447326 -3782 447562 -3546
rect 447646 -3782 447882 -3546
rect 451826 708442 452062 708678
rect 452146 708442 452382 708678
rect 451826 708122 452062 708358
rect 452146 708122 452382 708358
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4422 452062 -4186
rect 452146 -4422 452382 -4186
rect 451826 -4742 452062 -4506
rect 452146 -4742 452382 -4506
rect 456326 709402 456562 709638
rect 456646 709402 456882 709638
rect 456326 709082 456562 709318
rect 456646 709082 456882 709318
rect 456326 673718 456562 673954
rect 456646 673718 456882 673954
rect 456326 673398 456562 673634
rect 456646 673398 456882 673634
rect 456326 637718 456562 637954
rect 456646 637718 456882 637954
rect 456326 637398 456562 637634
rect 456646 637398 456882 637634
rect 456326 601718 456562 601954
rect 456646 601718 456882 601954
rect 456326 601398 456562 601634
rect 456646 601398 456882 601634
rect 456326 565718 456562 565954
rect 456646 565718 456882 565954
rect 456326 565398 456562 565634
rect 456646 565398 456882 565634
rect 456326 529718 456562 529954
rect 456646 529718 456882 529954
rect 456326 529398 456562 529634
rect 456646 529398 456882 529634
rect 456326 493718 456562 493954
rect 456646 493718 456882 493954
rect 456326 493398 456562 493634
rect 456646 493398 456882 493634
rect 456326 457718 456562 457954
rect 456646 457718 456882 457954
rect 456326 457398 456562 457634
rect 456646 457398 456882 457634
rect 456326 421718 456562 421954
rect 456646 421718 456882 421954
rect 456326 421398 456562 421634
rect 456646 421398 456882 421634
rect 456326 385718 456562 385954
rect 456646 385718 456882 385954
rect 456326 385398 456562 385634
rect 456646 385398 456882 385634
rect 456326 349718 456562 349954
rect 456646 349718 456882 349954
rect 456326 349398 456562 349634
rect 456646 349398 456882 349634
rect 456326 313718 456562 313954
rect 456646 313718 456882 313954
rect 456326 313398 456562 313634
rect 456646 313398 456882 313634
rect 456326 277718 456562 277954
rect 456646 277718 456882 277954
rect 456326 277398 456562 277634
rect 456646 277398 456882 277634
rect 456326 241718 456562 241954
rect 456646 241718 456882 241954
rect 456326 241398 456562 241634
rect 456646 241398 456882 241634
rect 456326 205718 456562 205954
rect 456646 205718 456882 205954
rect 456326 205398 456562 205634
rect 456646 205398 456882 205634
rect 456326 169718 456562 169954
rect 456646 169718 456882 169954
rect 456326 169398 456562 169634
rect 456646 169398 456882 169634
rect 456326 133718 456562 133954
rect 456646 133718 456882 133954
rect 456326 133398 456562 133634
rect 456646 133398 456882 133634
rect 456326 97718 456562 97954
rect 456646 97718 456882 97954
rect 456326 97398 456562 97634
rect 456646 97398 456882 97634
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5382 456562 -5146
rect 456646 -5382 456882 -5146
rect 456326 -5702 456562 -5466
rect 456646 -5702 456882 -5466
rect 460826 710362 461062 710598
rect 461146 710362 461382 710598
rect 460826 710042 461062 710278
rect 461146 710042 461382 710278
rect 460826 678218 461062 678454
rect 461146 678218 461382 678454
rect 460826 677898 461062 678134
rect 461146 677898 461382 678134
rect 460826 642218 461062 642454
rect 461146 642218 461382 642454
rect 460826 641898 461062 642134
rect 461146 641898 461382 642134
rect 460826 606218 461062 606454
rect 461146 606218 461382 606454
rect 460826 605898 461062 606134
rect 461146 605898 461382 606134
rect 460826 570218 461062 570454
rect 461146 570218 461382 570454
rect 460826 569898 461062 570134
rect 461146 569898 461382 570134
rect 460826 534218 461062 534454
rect 461146 534218 461382 534454
rect 460826 533898 461062 534134
rect 461146 533898 461382 534134
rect 460826 498218 461062 498454
rect 461146 498218 461382 498454
rect 460826 497898 461062 498134
rect 461146 497898 461382 498134
rect 460826 462218 461062 462454
rect 461146 462218 461382 462454
rect 460826 461898 461062 462134
rect 461146 461898 461382 462134
rect 460826 426218 461062 426454
rect 461146 426218 461382 426454
rect 460826 425898 461062 426134
rect 461146 425898 461382 426134
rect 460826 390218 461062 390454
rect 461146 390218 461382 390454
rect 460826 389898 461062 390134
rect 461146 389898 461382 390134
rect 460826 354218 461062 354454
rect 461146 354218 461382 354454
rect 460826 353898 461062 354134
rect 461146 353898 461382 354134
rect 460826 318218 461062 318454
rect 461146 318218 461382 318454
rect 460826 317898 461062 318134
rect 461146 317898 461382 318134
rect 460826 282218 461062 282454
rect 461146 282218 461382 282454
rect 460826 281898 461062 282134
rect 461146 281898 461382 282134
rect 460826 246218 461062 246454
rect 461146 246218 461382 246454
rect 460826 245898 461062 246134
rect 461146 245898 461382 246134
rect 460826 210218 461062 210454
rect 461146 210218 461382 210454
rect 460826 209898 461062 210134
rect 461146 209898 461382 210134
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 460826 138218 461062 138454
rect 461146 138218 461382 138454
rect 460826 137898 461062 138134
rect 461146 137898 461382 138134
rect 460826 102218 461062 102454
rect 461146 102218 461382 102454
rect 460826 101898 461062 102134
rect 461146 101898 461382 102134
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6342 461062 -6106
rect 461146 -6342 461382 -6106
rect 460826 -6662 461062 -6426
rect 461146 -6662 461382 -6426
rect 465326 711322 465562 711558
rect 465646 711322 465882 711558
rect 465326 711002 465562 711238
rect 465646 711002 465882 711238
rect 465326 682718 465562 682954
rect 465646 682718 465882 682954
rect 465326 682398 465562 682634
rect 465646 682398 465882 682634
rect 465326 646718 465562 646954
rect 465646 646718 465882 646954
rect 465326 646398 465562 646634
rect 465646 646398 465882 646634
rect 465326 610718 465562 610954
rect 465646 610718 465882 610954
rect 465326 610398 465562 610634
rect 465646 610398 465882 610634
rect 465326 574718 465562 574954
rect 465646 574718 465882 574954
rect 465326 574398 465562 574634
rect 465646 574398 465882 574634
rect 465326 538718 465562 538954
rect 465646 538718 465882 538954
rect 465326 538398 465562 538634
rect 465646 538398 465882 538634
rect 465326 502718 465562 502954
rect 465646 502718 465882 502954
rect 465326 502398 465562 502634
rect 465646 502398 465882 502634
rect 465326 466718 465562 466954
rect 465646 466718 465882 466954
rect 465326 466398 465562 466634
rect 465646 466398 465882 466634
rect 465326 430718 465562 430954
rect 465646 430718 465882 430954
rect 465326 430398 465562 430634
rect 465646 430398 465882 430634
rect 465326 394718 465562 394954
rect 465646 394718 465882 394954
rect 465326 394398 465562 394634
rect 465646 394398 465882 394634
rect 465326 358718 465562 358954
rect 465646 358718 465882 358954
rect 465326 358398 465562 358634
rect 465646 358398 465882 358634
rect 465326 322718 465562 322954
rect 465646 322718 465882 322954
rect 465326 322398 465562 322634
rect 465646 322398 465882 322634
rect 465326 286718 465562 286954
rect 465646 286718 465882 286954
rect 465326 286398 465562 286634
rect 465646 286398 465882 286634
rect 465326 250718 465562 250954
rect 465646 250718 465882 250954
rect 465326 250398 465562 250634
rect 465646 250398 465882 250634
rect 465326 214718 465562 214954
rect 465646 214718 465882 214954
rect 465326 214398 465562 214634
rect 465646 214398 465882 214634
rect 465326 178718 465562 178954
rect 465646 178718 465882 178954
rect 465326 178398 465562 178634
rect 465646 178398 465882 178634
rect 465326 142718 465562 142954
rect 465646 142718 465882 142954
rect 465326 142398 465562 142634
rect 465646 142398 465882 142634
rect 465326 106718 465562 106954
rect 465646 106718 465882 106954
rect 465326 106398 465562 106634
rect 465646 106398 465882 106634
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7302 465562 -7066
rect 465646 -7302 465882 -7066
rect 465326 -7622 465562 -7386
rect 465646 -7622 465882 -7386
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 474326 705562 474562 705798
rect 474646 705562 474882 705798
rect 474326 705242 474562 705478
rect 474646 705242 474882 705478
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 474326 655718 474562 655954
rect 474646 655718 474882 655954
rect 474326 655398 474562 655634
rect 474646 655398 474882 655634
rect 474326 619718 474562 619954
rect 474646 619718 474882 619954
rect 474326 619398 474562 619634
rect 474646 619398 474882 619634
rect 474326 583718 474562 583954
rect 474646 583718 474882 583954
rect 474326 583398 474562 583634
rect 474646 583398 474882 583634
rect 474326 547718 474562 547954
rect 474646 547718 474882 547954
rect 474326 547398 474562 547634
rect 474646 547398 474882 547634
rect 474326 511718 474562 511954
rect 474646 511718 474882 511954
rect 474326 511398 474562 511634
rect 474646 511398 474882 511634
rect 474326 475718 474562 475954
rect 474646 475718 474882 475954
rect 474326 475398 474562 475634
rect 474646 475398 474882 475634
rect 474326 439718 474562 439954
rect 474646 439718 474882 439954
rect 474326 439398 474562 439634
rect 474646 439398 474882 439634
rect 474326 403718 474562 403954
rect 474646 403718 474882 403954
rect 474326 403398 474562 403634
rect 474646 403398 474882 403634
rect 474326 367718 474562 367954
rect 474646 367718 474882 367954
rect 474326 367398 474562 367634
rect 474646 367398 474882 367634
rect 474326 331718 474562 331954
rect 474646 331718 474882 331954
rect 474326 331398 474562 331634
rect 474646 331398 474882 331634
rect 474326 295718 474562 295954
rect 474646 295718 474882 295954
rect 474326 295398 474562 295634
rect 474646 295398 474882 295634
rect 474326 259718 474562 259954
rect 474646 259718 474882 259954
rect 474326 259398 474562 259634
rect 474646 259398 474882 259634
rect 474326 223718 474562 223954
rect 474646 223718 474882 223954
rect 474326 223398 474562 223634
rect 474646 223398 474882 223634
rect 474326 187718 474562 187954
rect 474646 187718 474882 187954
rect 474326 187398 474562 187634
rect 474646 187398 474882 187634
rect 474326 151718 474562 151954
rect 474646 151718 474882 151954
rect 474326 151398 474562 151634
rect 474646 151398 474882 151634
rect 474326 115718 474562 115954
rect 474646 115718 474882 115954
rect 474326 115398 474562 115634
rect 474646 115398 474882 115634
rect 474326 79718 474562 79954
rect 474646 79718 474882 79954
rect 474326 79398 474562 79634
rect 474646 79398 474882 79634
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1542 474562 -1306
rect 474646 -1542 474882 -1306
rect 474326 -1862 474562 -1626
rect 474646 -1862 474882 -1626
rect 478826 706522 479062 706758
rect 479146 706522 479382 706758
rect 478826 706202 479062 706438
rect 479146 706202 479382 706438
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 478826 660218 479062 660454
rect 479146 660218 479382 660454
rect 478826 659898 479062 660134
rect 479146 659898 479382 660134
rect 478826 624218 479062 624454
rect 479146 624218 479382 624454
rect 478826 623898 479062 624134
rect 479146 623898 479382 624134
rect 478826 588218 479062 588454
rect 479146 588218 479382 588454
rect 478826 587898 479062 588134
rect 479146 587898 479382 588134
rect 478826 552218 479062 552454
rect 479146 552218 479382 552454
rect 478826 551898 479062 552134
rect 479146 551898 479382 552134
rect 478826 516218 479062 516454
rect 479146 516218 479382 516454
rect 478826 515898 479062 516134
rect 479146 515898 479382 516134
rect 478826 480218 479062 480454
rect 479146 480218 479382 480454
rect 478826 479898 479062 480134
rect 479146 479898 479382 480134
rect 478826 444218 479062 444454
rect 479146 444218 479382 444454
rect 478826 443898 479062 444134
rect 479146 443898 479382 444134
rect 478826 408218 479062 408454
rect 479146 408218 479382 408454
rect 478826 407898 479062 408134
rect 479146 407898 479382 408134
rect 478826 372218 479062 372454
rect 479146 372218 479382 372454
rect 478826 371898 479062 372134
rect 479146 371898 479382 372134
rect 478826 336218 479062 336454
rect 479146 336218 479382 336454
rect 478826 335898 479062 336134
rect 479146 335898 479382 336134
rect 478826 300218 479062 300454
rect 479146 300218 479382 300454
rect 478826 299898 479062 300134
rect 479146 299898 479382 300134
rect 478826 264218 479062 264454
rect 479146 264218 479382 264454
rect 478826 263898 479062 264134
rect 479146 263898 479382 264134
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 478826 192218 479062 192454
rect 479146 192218 479382 192454
rect 478826 191898 479062 192134
rect 479146 191898 479382 192134
rect 478826 156218 479062 156454
rect 479146 156218 479382 156454
rect 478826 155898 479062 156134
rect 479146 155898 479382 156134
rect 478826 120218 479062 120454
rect 479146 120218 479382 120454
rect 478826 119898 479062 120134
rect 479146 119898 479382 120134
rect 478826 84218 479062 84454
rect 479146 84218 479382 84454
rect 478826 83898 479062 84134
rect 479146 83898 479382 84134
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2502 479062 -2266
rect 479146 -2502 479382 -2266
rect 478826 -2822 479062 -2586
rect 479146 -2822 479382 -2586
rect 483326 707482 483562 707718
rect 483646 707482 483882 707718
rect 483326 707162 483562 707398
rect 483646 707162 483882 707398
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 483326 664718 483562 664954
rect 483646 664718 483882 664954
rect 483326 664398 483562 664634
rect 483646 664398 483882 664634
rect 483326 628718 483562 628954
rect 483646 628718 483882 628954
rect 483326 628398 483562 628634
rect 483646 628398 483882 628634
rect 483326 592718 483562 592954
rect 483646 592718 483882 592954
rect 483326 592398 483562 592634
rect 483646 592398 483882 592634
rect 483326 556718 483562 556954
rect 483646 556718 483882 556954
rect 483326 556398 483562 556634
rect 483646 556398 483882 556634
rect 483326 520718 483562 520954
rect 483646 520718 483882 520954
rect 483326 520398 483562 520634
rect 483646 520398 483882 520634
rect 483326 484718 483562 484954
rect 483646 484718 483882 484954
rect 483326 484398 483562 484634
rect 483646 484398 483882 484634
rect 483326 448718 483562 448954
rect 483646 448718 483882 448954
rect 483326 448398 483562 448634
rect 483646 448398 483882 448634
rect 483326 412718 483562 412954
rect 483646 412718 483882 412954
rect 483326 412398 483562 412634
rect 483646 412398 483882 412634
rect 483326 376718 483562 376954
rect 483646 376718 483882 376954
rect 483326 376398 483562 376634
rect 483646 376398 483882 376634
rect 483326 340718 483562 340954
rect 483646 340718 483882 340954
rect 483326 340398 483562 340634
rect 483646 340398 483882 340634
rect 483326 304718 483562 304954
rect 483646 304718 483882 304954
rect 483326 304398 483562 304634
rect 483646 304398 483882 304634
rect 483326 268718 483562 268954
rect 483646 268718 483882 268954
rect 483326 268398 483562 268634
rect 483646 268398 483882 268634
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 483326 124718 483562 124954
rect 483646 124718 483882 124954
rect 483326 124398 483562 124634
rect 483646 124398 483882 124634
rect 483326 88718 483562 88954
rect 483646 88718 483882 88954
rect 483326 88398 483562 88634
rect 483646 88398 483882 88634
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3462 483562 -3226
rect 483646 -3462 483882 -3226
rect 483326 -3782 483562 -3546
rect 483646 -3782 483882 -3546
rect 487826 708442 488062 708678
rect 488146 708442 488382 708678
rect 487826 708122 488062 708358
rect 488146 708122 488382 708358
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4422 488062 -4186
rect 488146 -4422 488382 -4186
rect 487826 -4742 488062 -4506
rect 488146 -4742 488382 -4506
rect 492326 709402 492562 709638
rect 492646 709402 492882 709638
rect 492326 709082 492562 709318
rect 492646 709082 492882 709318
rect 492326 673718 492562 673954
rect 492646 673718 492882 673954
rect 492326 673398 492562 673634
rect 492646 673398 492882 673634
rect 492326 637718 492562 637954
rect 492646 637718 492882 637954
rect 492326 637398 492562 637634
rect 492646 637398 492882 637634
rect 492326 601718 492562 601954
rect 492646 601718 492882 601954
rect 492326 601398 492562 601634
rect 492646 601398 492882 601634
rect 492326 565718 492562 565954
rect 492646 565718 492882 565954
rect 492326 565398 492562 565634
rect 492646 565398 492882 565634
rect 492326 529718 492562 529954
rect 492646 529718 492882 529954
rect 492326 529398 492562 529634
rect 492646 529398 492882 529634
rect 492326 493718 492562 493954
rect 492646 493718 492882 493954
rect 492326 493398 492562 493634
rect 492646 493398 492882 493634
rect 492326 457718 492562 457954
rect 492646 457718 492882 457954
rect 492326 457398 492562 457634
rect 492646 457398 492882 457634
rect 492326 421718 492562 421954
rect 492646 421718 492882 421954
rect 492326 421398 492562 421634
rect 492646 421398 492882 421634
rect 492326 385718 492562 385954
rect 492646 385718 492882 385954
rect 492326 385398 492562 385634
rect 492646 385398 492882 385634
rect 492326 349718 492562 349954
rect 492646 349718 492882 349954
rect 492326 349398 492562 349634
rect 492646 349398 492882 349634
rect 492326 313718 492562 313954
rect 492646 313718 492882 313954
rect 492326 313398 492562 313634
rect 492646 313398 492882 313634
rect 492326 277718 492562 277954
rect 492646 277718 492882 277954
rect 492326 277398 492562 277634
rect 492646 277398 492882 277634
rect 492326 241718 492562 241954
rect 492646 241718 492882 241954
rect 492326 241398 492562 241634
rect 492646 241398 492882 241634
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 492326 133718 492562 133954
rect 492646 133718 492882 133954
rect 492326 133398 492562 133634
rect 492646 133398 492882 133634
rect 492326 97718 492562 97954
rect 492646 97718 492882 97954
rect 492326 97398 492562 97634
rect 492646 97398 492882 97634
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5382 492562 -5146
rect 492646 -5382 492882 -5146
rect 492326 -5702 492562 -5466
rect 492646 -5702 492882 -5466
rect 496826 710362 497062 710598
rect 497146 710362 497382 710598
rect 496826 710042 497062 710278
rect 497146 710042 497382 710278
rect 496826 678218 497062 678454
rect 497146 678218 497382 678454
rect 496826 677898 497062 678134
rect 497146 677898 497382 678134
rect 496826 642218 497062 642454
rect 497146 642218 497382 642454
rect 496826 641898 497062 642134
rect 497146 641898 497382 642134
rect 496826 606218 497062 606454
rect 497146 606218 497382 606454
rect 496826 605898 497062 606134
rect 497146 605898 497382 606134
rect 496826 570218 497062 570454
rect 497146 570218 497382 570454
rect 496826 569898 497062 570134
rect 497146 569898 497382 570134
rect 496826 534218 497062 534454
rect 497146 534218 497382 534454
rect 496826 533898 497062 534134
rect 497146 533898 497382 534134
rect 496826 498218 497062 498454
rect 497146 498218 497382 498454
rect 496826 497898 497062 498134
rect 497146 497898 497382 498134
rect 496826 462218 497062 462454
rect 497146 462218 497382 462454
rect 496826 461898 497062 462134
rect 497146 461898 497382 462134
rect 496826 426218 497062 426454
rect 497146 426218 497382 426454
rect 496826 425898 497062 426134
rect 497146 425898 497382 426134
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 496826 354218 497062 354454
rect 497146 354218 497382 354454
rect 496826 353898 497062 354134
rect 497146 353898 497382 354134
rect 496826 318218 497062 318454
rect 497146 318218 497382 318454
rect 496826 317898 497062 318134
rect 497146 317898 497382 318134
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 496826 246218 497062 246454
rect 497146 246218 497382 246454
rect 496826 245898 497062 246134
rect 497146 245898 497382 246134
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 496826 138218 497062 138454
rect 497146 138218 497382 138454
rect 496826 137898 497062 138134
rect 497146 137898 497382 138134
rect 496826 102218 497062 102454
rect 497146 102218 497382 102454
rect 496826 101898 497062 102134
rect 497146 101898 497382 102134
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6342 497062 -6106
rect 497146 -6342 497382 -6106
rect 496826 -6662 497062 -6426
rect 497146 -6662 497382 -6426
rect 501326 711322 501562 711558
rect 501646 711322 501882 711558
rect 501326 711002 501562 711238
rect 501646 711002 501882 711238
rect 501326 682718 501562 682954
rect 501646 682718 501882 682954
rect 501326 682398 501562 682634
rect 501646 682398 501882 682634
rect 501326 646718 501562 646954
rect 501646 646718 501882 646954
rect 501326 646398 501562 646634
rect 501646 646398 501882 646634
rect 501326 610718 501562 610954
rect 501646 610718 501882 610954
rect 501326 610398 501562 610634
rect 501646 610398 501882 610634
rect 501326 574718 501562 574954
rect 501646 574718 501882 574954
rect 501326 574398 501562 574634
rect 501646 574398 501882 574634
rect 501326 538718 501562 538954
rect 501646 538718 501882 538954
rect 501326 538398 501562 538634
rect 501646 538398 501882 538634
rect 501326 502718 501562 502954
rect 501646 502718 501882 502954
rect 501326 502398 501562 502634
rect 501646 502398 501882 502634
rect 501326 466718 501562 466954
rect 501646 466718 501882 466954
rect 501326 466398 501562 466634
rect 501646 466398 501882 466634
rect 501326 430718 501562 430954
rect 501646 430718 501882 430954
rect 501326 430398 501562 430634
rect 501646 430398 501882 430634
rect 501326 394718 501562 394954
rect 501646 394718 501882 394954
rect 501326 394398 501562 394634
rect 501646 394398 501882 394634
rect 501326 358718 501562 358954
rect 501646 358718 501882 358954
rect 501326 358398 501562 358634
rect 501646 358398 501882 358634
rect 501326 322718 501562 322954
rect 501646 322718 501882 322954
rect 501326 322398 501562 322634
rect 501646 322398 501882 322634
rect 501326 286718 501562 286954
rect 501646 286718 501882 286954
rect 501326 286398 501562 286634
rect 501646 286398 501882 286634
rect 501326 250718 501562 250954
rect 501646 250718 501882 250954
rect 501326 250398 501562 250634
rect 501646 250398 501882 250634
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 501326 142718 501562 142954
rect 501646 142718 501882 142954
rect 501326 142398 501562 142634
rect 501646 142398 501882 142634
rect 501326 106718 501562 106954
rect 501646 106718 501882 106954
rect 501326 106398 501562 106634
rect 501646 106398 501882 106634
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7302 501562 -7066
rect 501646 -7302 501882 -7066
rect 501326 -7622 501562 -7386
rect 501646 -7622 501882 -7386
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 510326 705562 510562 705798
rect 510646 705562 510882 705798
rect 510326 705242 510562 705478
rect 510646 705242 510882 705478
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 510326 619718 510562 619954
rect 510646 619718 510882 619954
rect 510326 619398 510562 619634
rect 510646 619398 510882 619634
rect 510326 583718 510562 583954
rect 510646 583718 510882 583954
rect 510326 583398 510562 583634
rect 510646 583398 510882 583634
rect 510326 547718 510562 547954
rect 510646 547718 510882 547954
rect 510326 547398 510562 547634
rect 510646 547398 510882 547634
rect 510326 511718 510562 511954
rect 510646 511718 510882 511954
rect 510326 511398 510562 511634
rect 510646 511398 510882 511634
rect 510326 475718 510562 475954
rect 510646 475718 510882 475954
rect 510326 475398 510562 475634
rect 510646 475398 510882 475634
rect 510326 439718 510562 439954
rect 510646 439718 510882 439954
rect 510326 439398 510562 439634
rect 510646 439398 510882 439634
rect 510326 403718 510562 403954
rect 510646 403718 510882 403954
rect 510326 403398 510562 403634
rect 510646 403398 510882 403634
rect 510326 367718 510562 367954
rect 510646 367718 510882 367954
rect 510326 367398 510562 367634
rect 510646 367398 510882 367634
rect 510326 331718 510562 331954
rect 510646 331718 510882 331954
rect 510326 331398 510562 331634
rect 510646 331398 510882 331634
rect 510326 295718 510562 295954
rect 510646 295718 510882 295954
rect 510326 295398 510562 295634
rect 510646 295398 510882 295634
rect 510326 259718 510562 259954
rect 510646 259718 510882 259954
rect 510326 259398 510562 259634
rect 510646 259398 510882 259634
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 510326 151718 510562 151954
rect 510646 151718 510882 151954
rect 510326 151398 510562 151634
rect 510646 151398 510882 151634
rect 510326 115718 510562 115954
rect 510646 115718 510882 115954
rect 510326 115398 510562 115634
rect 510646 115398 510882 115634
rect 510326 79718 510562 79954
rect 510646 79718 510882 79954
rect 510326 79398 510562 79634
rect 510646 79398 510882 79634
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1542 510562 -1306
rect 510646 -1542 510882 -1306
rect 510326 -1862 510562 -1626
rect 510646 -1862 510882 -1626
rect 514826 706522 515062 706758
rect 515146 706522 515382 706758
rect 514826 706202 515062 706438
rect 515146 706202 515382 706438
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 514826 624218 515062 624454
rect 515146 624218 515382 624454
rect 514826 623898 515062 624134
rect 515146 623898 515382 624134
rect 514826 588218 515062 588454
rect 515146 588218 515382 588454
rect 514826 587898 515062 588134
rect 515146 587898 515382 588134
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 514826 516218 515062 516454
rect 515146 516218 515382 516454
rect 514826 515898 515062 516134
rect 515146 515898 515382 516134
rect 514826 480218 515062 480454
rect 515146 480218 515382 480454
rect 514826 479898 515062 480134
rect 515146 479898 515382 480134
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 514826 408218 515062 408454
rect 515146 408218 515382 408454
rect 514826 407898 515062 408134
rect 515146 407898 515382 408134
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 514826 264218 515062 264454
rect 515146 264218 515382 264454
rect 514826 263898 515062 264134
rect 515146 263898 515382 264134
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2502 515062 -2266
rect 515146 -2502 515382 -2266
rect 514826 -2822 515062 -2586
rect 515146 -2822 515382 -2586
rect 519326 707482 519562 707718
rect 519646 707482 519882 707718
rect 519326 707162 519562 707398
rect 519646 707162 519882 707398
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 519326 628718 519562 628954
rect 519646 628718 519882 628954
rect 519326 628398 519562 628634
rect 519646 628398 519882 628634
rect 519326 592718 519562 592954
rect 519646 592718 519882 592954
rect 519326 592398 519562 592634
rect 519646 592398 519882 592634
rect 519326 556718 519562 556954
rect 519646 556718 519882 556954
rect 519326 556398 519562 556634
rect 519646 556398 519882 556634
rect 519326 520718 519562 520954
rect 519646 520718 519882 520954
rect 519326 520398 519562 520634
rect 519646 520398 519882 520634
rect 519326 484718 519562 484954
rect 519646 484718 519882 484954
rect 519326 484398 519562 484634
rect 519646 484398 519882 484634
rect 519326 448718 519562 448954
rect 519646 448718 519882 448954
rect 519326 448398 519562 448634
rect 519646 448398 519882 448634
rect 519326 412718 519562 412954
rect 519646 412718 519882 412954
rect 519326 412398 519562 412634
rect 519646 412398 519882 412634
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 519326 268718 519562 268954
rect 519646 268718 519882 268954
rect 519326 268398 519562 268634
rect 519646 268398 519882 268634
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 519326 124718 519562 124954
rect 519646 124718 519882 124954
rect 519326 124398 519562 124634
rect 519646 124398 519882 124634
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3462 519562 -3226
rect 519646 -3462 519882 -3226
rect 519326 -3782 519562 -3546
rect 519646 -3782 519882 -3546
rect 523826 708442 524062 708678
rect 524146 708442 524382 708678
rect 523826 708122 524062 708358
rect 524146 708122 524382 708358
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4422 524062 -4186
rect 524146 -4422 524382 -4186
rect 523826 -4742 524062 -4506
rect 524146 -4742 524382 -4506
rect 528326 709402 528562 709638
rect 528646 709402 528882 709638
rect 528326 709082 528562 709318
rect 528646 709082 528882 709318
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 528326 565718 528562 565954
rect 528646 565718 528882 565954
rect 528326 565398 528562 565634
rect 528646 565398 528882 565634
rect 528326 529718 528562 529954
rect 528646 529718 528882 529954
rect 528326 529398 528562 529634
rect 528646 529398 528882 529634
rect 528326 493718 528562 493954
rect 528646 493718 528882 493954
rect 528326 493398 528562 493634
rect 528646 493398 528882 493634
rect 528326 457718 528562 457954
rect 528646 457718 528882 457954
rect 528326 457398 528562 457634
rect 528646 457398 528882 457634
rect 528326 421718 528562 421954
rect 528646 421718 528882 421954
rect 528326 421398 528562 421634
rect 528646 421398 528882 421634
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 528326 277718 528562 277954
rect 528646 277718 528882 277954
rect 528326 277398 528562 277634
rect 528646 277398 528882 277634
rect 528326 241718 528562 241954
rect 528646 241718 528882 241954
rect 528326 241398 528562 241634
rect 528646 241398 528882 241634
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 528326 133718 528562 133954
rect 528646 133718 528882 133954
rect 528326 133398 528562 133634
rect 528646 133398 528882 133634
rect 528326 97718 528562 97954
rect 528646 97718 528882 97954
rect 528326 97398 528562 97634
rect 528646 97398 528882 97634
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5382 528562 -5146
rect 528646 -5382 528882 -5146
rect 528326 -5702 528562 -5466
rect 528646 -5702 528882 -5466
rect 532826 710362 533062 710598
rect 533146 710362 533382 710598
rect 532826 710042 533062 710278
rect 533146 710042 533382 710278
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 532826 570218 533062 570454
rect 533146 570218 533382 570454
rect 532826 569898 533062 570134
rect 533146 569898 533382 570134
rect 532826 534218 533062 534454
rect 533146 534218 533382 534454
rect 532826 533898 533062 534134
rect 533146 533898 533382 534134
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 532826 462218 533062 462454
rect 533146 462218 533382 462454
rect 532826 461898 533062 462134
rect 533146 461898 533382 462134
rect 532826 426218 533062 426454
rect 533146 426218 533382 426454
rect 532826 425898 533062 426134
rect 533146 425898 533382 426134
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 532826 246218 533062 246454
rect 533146 246218 533382 246454
rect 532826 245898 533062 246134
rect 533146 245898 533382 246134
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 532826 138218 533062 138454
rect 533146 138218 533382 138454
rect 532826 137898 533062 138134
rect 533146 137898 533382 138134
rect 532826 102218 533062 102454
rect 533146 102218 533382 102454
rect 532826 101898 533062 102134
rect 533146 101898 533382 102134
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6342 533062 -6106
rect 533146 -6342 533382 -6106
rect 532826 -6662 533062 -6426
rect 533146 -6662 533382 -6426
rect 537326 711322 537562 711558
rect 537646 711322 537882 711558
rect 537326 711002 537562 711238
rect 537646 711002 537882 711238
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 537326 250718 537562 250954
rect 537646 250718 537882 250954
rect 537326 250398 537562 250634
rect 537646 250398 537882 250634
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 537326 142718 537562 142954
rect 537646 142718 537882 142954
rect 537326 142398 537562 142634
rect 537646 142398 537882 142634
rect 537326 106718 537562 106954
rect 537646 106718 537882 106954
rect 537326 106398 537562 106634
rect 537646 106398 537882 106634
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7302 537562 -7066
rect 537646 -7302 537882 -7066
rect 537326 -7622 537562 -7386
rect 537646 -7622 537882 -7386
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 546326 705562 546562 705798
rect 546646 705562 546882 705798
rect 546326 705242 546562 705478
rect 546646 705242 546882 705478
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 546326 259718 546562 259954
rect 546646 259718 546882 259954
rect 546326 259398 546562 259634
rect 546646 259398 546882 259634
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1542 546562 -1306
rect 546646 -1542 546882 -1306
rect 546326 -1862 546562 -1626
rect 546646 -1862 546882 -1626
rect 550826 706522 551062 706758
rect 551146 706522 551382 706758
rect 550826 706202 551062 706438
rect 551146 706202 551382 706438
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 550826 300218 551062 300454
rect 551146 300218 551382 300454
rect 550826 299898 551062 300134
rect 551146 299898 551382 300134
rect 550826 264218 551062 264454
rect 551146 264218 551382 264454
rect 550826 263898 551062 264134
rect 551146 263898 551382 264134
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2502 551062 -2266
rect 551146 -2502 551382 -2266
rect 550826 -2822 551062 -2586
rect 551146 -2822 551382 -2586
rect 555326 707482 555562 707718
rect 555646 707482 555882 707718
rect 555326 707162 555562 707398
rect 555646 707162 555882 707398
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3462 555562 -3226
rect 555646 -3462 555882 -3226
rect 555326 -3782 555562 -3546
rect 555646 -3782 555882 -3546
rect 559826 708442 560062 708678
rect 560146 708442 560382 708678
rect 559826 708122 560062 708358
rect 560146 708122 560382 708358
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4422 560062 -4186
rect 560146 -4422 560382 -4186
rect 559826 -4742 560062 -4506
rect 560146 -4742 560382 -4506
rect 564326 709402 564562 709638
rect 564646 709402 564882 709638
rect 564326 709082 564562 709318
rect 564646 709082 564882 709318
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5382 564562 -5146
rect 564646 -5382 564882 -5146
rect 564326 -5702 564562 -5466
rect 564646 -5702 564882 -5466
rect 568826 710362 569062 710598
rect 569146 710362 569382 710598
rect 568826 710042 569062 710278
rect 569146 710042 569382 710278
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6342 569062 -6106
rect 569146 -6342 569382 -6106
rect 568826 -6662 569062 -6426
rect 569146 -6662 569382 -6426
rect 573326 711322 573562 711558
rect 573646 711322 573882 711558
rect 573326 711002 573562 711238
rect 573646 711002 573882 711238
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7302 573562 -7066
rect 573646 -7302 573882 -7066
rect 573326 -7622 573562 -7386
rect 573646 -7622 573882 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 691718 586538 691954
rect 586622 691718 586858 691954
rect 586302 691398 586538 691634
rect 586622 691398 586858 691634
rect 586302 655718 586538 655954
rect 586622 655718 586858 655954
rect 586302 655398 586538 655634
rect 586622 655398 586858 655634
rect 586302 619718 586538 619954
rect 586622 619718 586858 619954
rect 586302 619398 586538 619634
rect 586622 619398 586858 619634
rect 586302 583718 586538 583954
rect 586622 583718 586858 583954
rect 586302 583398 586538 583634
rect 586622 583398 586858 583634
rect 586302 547718 586538 547954
rect 586622 547718 586858 547954
rect 586302 547398 586538 547634
rect 586622 547398 586858 547634
rect 586302 511718 586538 511954
rect 586622 511718 586858 511954
rect 586302 511398 586538 511634
rect 586622 511398 586858 511634
rect 586302 475718 586538 475954
rect 586622 475718 586858 475954
rect 586302 475398 586538 475634
rect 586622 475398 586858 475634
rect 586302 439718 586538 439954
rect 586622 439718 586858 439954
rect 586302 439398 586538 439634
rect 586622 439398 586858 439634
rect 586302 403718 586538 403954
rect 586622 403718 586858 403954
rect 586302 403398 586538 403634
rect 586622 403398 586858 403634
rect 586302 367718 586538 367954
rect 586622 367718 586858 367954
rect 586302 367398 586538 367634
rect 586622 367398 586858 367634
rect 586302 331718 586538 331954
rect 586622 331718 586858 331954
rect 586302 331398 586538 331634
rect 586622 331398 586858 331634
rect 586302 295718 586538 295954
rect 586622 295718 586858 295954
rect 586302 295398 586538 295634
rect 586622 295398 586858 295634
rect 586302 259718 586538 259954
rect 586622 259718 586858 259954
rect 586302 259398 586538 259634
rect 586622 259398 586858 259634
rect 586302 223718 586538 223954
rect 586622 223718 586858 223954
rect 586302 223398 586538 223634
rect 586622 223398 586858 223634
rect 586302 187718 586538 187954
rect 586622 187718 586858 187954
rect 586302 187398 586538 187634
rect 586622 187398 586858 187634
rect 586302 151718 586538 151954
rect 586622 151718 586858 151954
rect 586302 151398 586538 151634
rect 586622 151398 586858 151634
rect 586302 115718 586538 115954
rect 586622 115718 586858 115954
rect 586302 115398 586538 115634
rect 586622 115398 586858 115634
rect 586302 79718 586538 79954
rect 586622 79718 586858 79954
rect 586302 79398 586538 79634
rect 586622 79398 586858 79634
rect 586302 43718 586538 43954
rect 586622 43718 586858 43954
rect 586302 43398 586538 43634
rect 586622 43398 586858 43634
rect 586302 7718 586538 7954
rect 586622 7718 586858 7954
rect 586302 7398 586538 7634
rect 586622 7398 586858 7634
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 696218 587498 696454
rect 587582 696218 587818 696454
rect 587262 695898 587498 696134
rect 587582 695898 587818 696134
rect 587262 660218 587498 660454
rect 587582 660218 587818 660454
rect 587262 659898 587498 660134
rect 587582 659898 587818 660134
rect 587262 624218 587498 624454
rect 587582 624218 587818 624454
rect 587262 623898 587498 624134
rect 587582 623898 587818 624134
rect 587262 588218 587498 588454
rect 587582 588218 587818 588454
rect 587262 587898 587498 588134
rect 587582 587898 587818 588134
rect 587262 552218 587498 552454
rect 587582 552218 587818 552454
rect 587262 551898 587498 552134
rect 587582 551898 587818 552134
rect 587262 516218 587498 516454
rect 587582 516218 587818 516454
rect 587262 515898 587498 516134
rect 587582 515898 587818 516134
rect 587262 480218 587498 480454
rect 587582 480218 587818 480454
rect 587262 479898 587498 480134
rect 587582 479898 587818 480134
rect 587262 444218 587498 444454
rect 587582 444218 587818 444454
rect 587262 443898 587498 444134
rect 587582 443898 587818 444134
rect 587262 408218 587498 408454
rect 587582 408218 587818 408454
rect 587262 407898 587498 408134
rect 587582 407898 587818 408134
rect 587262 372218 587498 372454
rect 587582 372218 587818 372454
rect 587262 371898 587498 372134
rect 587582 371898 587818 372134
rect 587262 336218 587498 336454
rect 587582 336218 587818 336454
rect 587262 335898 587498 336134
rect 587582 335898 587818 336134
rect 587262 300218 587498 300454
rect 587582 300218 587818 300454
rect 587262 299898 587498 300134
rect 587582 299898 587818 300134
rect 587262 264218 587498 264454
rect 587582 264218 587818 264454
rect 587262 263898 587498 264134
rect 587582 263898 587818 264134
rect 587262 228218 587498 228454
rect 587582 228218 587818 228454
rect 587262 227898 587498 228134
rect 587582 227898 587818 228134
rect 587262 192218 587498 192454
rect 587582 192218 587818 192454
rect 587262 191898 587498 192134
rect 587582 191898 587818 192134
rect 587262 156218 587498 156454
rect 587582 156218 587818 156454
rect 587262 155898 587498 156134
rect 587582 155898 587818 156134
rect 587262 120218 587498 120454
rect 587582 120218 587818 120454
rect 587262 119898 587498 120134
rect 587582 119898 587818 120134
rect 587262 84218 587498 84454
rect 587582 84218 587818 84454
rect 587262 83898 587498 84134
rect 587582 83898 587818 84134
rect 587262 48218 587498 48454
rect 587582 48218 587818 48454
rect 587262 47898 587498 48134
rect 587582 47898 587818 48134
rect 587262 12218 587498 12454
rect 587582 12218 587818 12454
rect 587262 11898 587498 12134
rect 587582 11898 587818 12134
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 700718 588458 700954
rect 588542 700718 588778 700954
rect 588222 700398 588458 700634
rect 588542 700398 588778 700634
rect 588222 664718 588458 664954
rect 588542 664718 588778 664954
rect 588222 664398 588458 664634
rect 588542 664398 588778 664634
rect 588222 628718 588458 628954
rect 588542 628718 588778 628954
rect 588222 628398 588458 628634
rect 588542 628398 588778 628634
rect 588222 592718 588458 592954
rect 588542 592718 588778 592954
rect 588222 592398 588458 592634
rect 588542 592398 588778 592634
rect 588222 556718 588458 556954
rect 588542 556718 588778 556954
rect 588222 556398 588458 556634
rect 588542 556398 588778 556634
rect 588222 520718 588458 520954
rect 588542 520718 588778 520954
rect 588222 520398 588458 520634
rect 588542 520398 588778 520634
rect 588222 484718 588458 484954
rect 588542 484718 588778 484954
rect 588222 484398 588458 484634
rect 588542 484398 588778 484634
rect 588222 448718 588458 448954
rect 588542 448718 588778 448954
rect 588222 448398 588458 448634
rect 588542 448398 588778 448634
rect 588222 412718 588458 412954
rect 588542 412718 588778 412954
rect 588222 412398 588458 412634
rect 588542 412398 588778 412634
rect 588222 376718 588458 376954
rect 588542 376718 588778 376954
rect 588222 376398 588458 376634
rect 588542 376398 588778 376634
rect 588222 340718 588458 340954
rect 588542 340718 588778 340954
rect 588222 340398 588458 340634
rect 588542 340398 588778 340634
rect 588222 304718 588458 304954
rect 588542 304718 588778 304954
rect 588222 304398 588458 304634
rect 588542 304398 588778 304634
rect 588222 268718 588458 268954
rect 588542 268718 588778 268954
rect 588222 268398 588458 268634
rect 588542 268398 588778 268634
rect 588222 232718 588458 232954
rect 588542 232718 588778 232954
rect 588222 232398 588458 232634
rect 588542 232398 588778 232634
rect 588222 196718 588458 196954
rect 588542 196718 588778 196954
rect 588222 196398 588458 196634
rect 588542 196398 588778 196634
rect 588222 160718 588458 160954
rect 588542 160718 588778 160954
rect 588222 160398 588458 160634
rect 588542 160398 588778 160634
rect 588222 124718 588458 124954
rect 588542 124718 588778 124954
rect 588222 124398 588458 124634
rect 588542 124398 588778 124634
rect 588222 88718 588458 88954
rect 588542 88718 588778 88954
rect 588222 88398 588458 88634
rect 588542 88398 588778 88634
rect 588222 52718 588458 52954
rect 588542 52718 588778 52954
rect 588222 52398 588458 52634
rect 588542 52398 588778 52634
rect 588222 16718 588458 16954
rect 588542 16718 588778 16954
rect 588222 16398 588458 16634
rect 588542 16398 588778 16634
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 669218 589418 669454
rect 589502 669218 589738 669454
rect 589182 668898 589418 669134
rect 589502 668898 589738 669134
rect 589182 633218 589418 633454
rect 589502 633218 589738 633454
rect 589182 632898 589418 633134
rect 589502 632898 589738 633134
rect 589182 597218 589418 597454
rect 589502 597218 589738 597454
rect 589182 596898 589418 597134
rect 589502 596898 589738 597134
rect 589182 561218 589418 561454
rect 589502 561218 589738 561454
rect 589182 560898 589418 561134
rect 589502 560898 589738 561134
rect 589182 525218 589418 525454
rect 589502 525218 589738 525454
rect 589182 524898 589418 525134
rect 589502 524898 589738 525134
rect 589182 489218 589418 489454
rect 589502 489218 589738 489454
rect 589182 488898 589418 489134
rect 589502 488898 589738 489134
rect 589182 453218 589418 453454
rect 589502 453218 589738 453454
rect 589182 452898 589418 453134
rect 589502 452898 589738 453134
rect 589182 417218 589418 417454
rect 589502 417218 589738 417454
rect 589182 416898 589418 417134
rect 589502 416898 589738 417134
rect 589182 381218 589418 381454
rect 589502 381218 589738 381454
rect 589182 380898 589418 381134
rect 589502 380898 589738 381134
rect 589182 345218 589418 345454
rect 589502 345218 589738 345454
rect 589182 344898 589418 345134
rect 589502 344898 589738 345134
rect 589182 309218 589418 309454
rect 589502 309218 589738 309454
rect 589182 308898 589418 309134
rect 589502 308898 589738 309134
rect 589182 273218 589418 273454
rect 589502 273218 589738 273454
rect 589182 272898 589418 273134
rect 589502 272898 589738 273134
rect 589182 237218 589418 237454
rect 589502 237218 589738 237454
rect 589182 236898 589418 237134
rect 589502 236898 589738 237134
rect 589182 201218 589418 201454
rect 589502 201218 589738 201454
rect 589182 200898 589418 201134
rect 589502 200898 589738 201134
rect 589182 165218 589418 165454
rect 589502 165218 589738 165454
rect 589182 164898 589418 165134
rect 589502 164898 589738 165134
rect 589182 129218 589418 129454
rect 589502 129218 589738 129454
rect 589182 128898 589418 129134
rect 589502 128898 589738 129134
rect 589182 93218 589418 93454
rect 589502 93218 589738 93454
rect 589182 92898 589418 93134
rect 589502 92898 589738 93134
rect 589182 57218 589418 57454
rect 589502 57218 589738 57454
rect 589182 56898 589418 57134
rect 589502 56898 589738 57134
rect 589182 21218 589418 21454
rect 589502 21218 589738 21454
rect 589182 20898 589418 21134
rect 589502 20898 589738 21134
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 673718 590378 673954
rect 590462 673718 590698 673954
rect 590142 673398 590378 673634
rect 590462 673398 590698 673634
rect 590142 637718 590378 637954
rect 590462 637718 590698 637954
rect 590142 637398 590378 637634
rect 590462 637398 590698 637634
rect 590142 601718 590378 601954
rect 590462 601718 590698 601954
rect 590142 601398 590378 601634
rect 590462 601398 590698 601634
rect 590142 565718 590378 565954
rect 590462 565718 590698 565954
rect 590142 565398 590378 565634
rect 590462 565398 590698 565634
rect 590142 529718 590378 529954
rect 590462 529718 590698 529954
rect 590142 529398 590378 529634
rect 590462 529398 590698 529634
rect 590142 493718 590378 493954
rect 590462 493718 590698 493954
rect 590142 493398 590378 493634
rect 590462 493398 590698 493634
rect 590142 457718 590378 457954
rect 590462 457718 590698 457954
rect 590142 457398 590378 457634
rect 590462 457398 590698 457634
rect 590142 421718 590378 421954
rect 590462 421718 590698 421954
rect 590142 421398 590378 421634
rect 590462 421398 590698 421634
rect 590142 385718 590378 385954
rect 590462 385718 590698 385954
rect 590142 385398 590378 385634
rect 590462 385398 590698 385634
rect 590142 349718 590378 349954
rect 590462 349718 590698 349954
rect 590142 349398 590378 349634
rect 590462 349398 590698 349634
rect 590142 313718 590378 313954
rect 590462 313718 590698 313954
rect 590142 313398 590378 313634
rect 590462 313398 590698 313634
rect 590142 277718 590378 277954
rect 590462 277718 590698 277954
rect 590142 277398 590378 277634
rect 590462 277398 590698 277634
rect 590142 241718 590378 241954
rect 590462 241718 590698 241954
rect 590142 241398 590378 241634
rect 590462 241398 590698 241634
rect 590142 205718 590378 205954
rect 590462 205718 590698 205954
rect 590142 205398 590378 205634
rect 590462 205398 590698 205634
rect 590142 169718 590378 169954
rect 590462 169718 590698 169954
rect 590142 169398 590378 169634
rect 590462 169398 590698 169634
rect 590142 133718 590378 133954
rect 590462 133718 590698 133954
rect 590142 133398 590378 133634
rect 590462 133398 590698 133634
rect 590142 97718 590378 97954
rect 590462 97718 590698 97954
rect 590142 97398 590378 97634
rect 590462 97398 590698 97634
rect 590142 61718 590378 61954
rect 590462 61718 590698 61954
rect 590142 61398 590378 61634
rect 590462 61398 590698 61634
rect 590142 25718 590378 25954
rect 590462 25718 590698 25954
rect 590142 25398 590378 25634
rect 590462 25398 590698 25634
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 678218 591338 678454
rect 591422 678218 591658 678454
rect 591102 677898 591338 678134
rect 591422 677898 591658 678134
rect 591102 642218 591338 642454
rect 591422 642218 591658 642454
rect 591102 641898 591338 642134
rect 591422 641898 591658 642134
rect 591102 606218 591338 606454
rect 591422 606218 591658 606454
rect 591102 605898 591338 606134
rect 591422 605898 591658 606134
rect 591102 570218 591338 570454
rect 591422 570218 591658 570454
rect 591102 569898 591338 570134
rect 591422 569898 591658 570134
rect 591102 534218 591338 534454
rect 591422 534218 591658 534454
rect 591102 533898 591338 534134
rect 591422 533898 591658 534134
rect 591102 498218 591338 498454
rect 591422 498218 591658 498454
rect 591102 497898 591338 498134
rect 591422 497898 591658 498134
rect 591102 462218 591338 462454
rect 591422 462218 591658 462454
rect 591102 461898 591338 462134
rect 591422 461898 591658 462134
rect 591102 426218 591338 426454
rect 591422 426218 591658 426454
rect 591102 425898 591338 426134
rect 591422 425898 591658 426134
rect 591102 390218 591338 390454
rect 591422 390218 591658 390454
rect 591102 389898 591338 390134
rect 591422 389898 591658 390134
rect 591102 354218 591338 354454
rect 591422 354218 591658 354454
rect 591102 353898 591338 354134
rect 591422 353898 591658 354134
rect 591102 318218 591338 318454
rect 591422 318218 591658 318454
rect 591102 317898 591338 318134
rect 591422 317898 591658 318134
rect 591102 282218 591338 282454
rect 591422 282218 591658 282454
rect 591102 281898 591338 282134
rect 591422 281898 591658 282134
rect 591102 246218 591338 246454
rect 591422 246218 591658 246454
rect 591102 245898 591338 246134
rect 591422 245898 591658 246134
rect 591102 210218 591338 210454
rect 591422 210218 591658 210454
rect 591102 209898 591338 210134
rect 591422 209898 591658 210134
rect 591102 174218 591338 174454
rect 591422 174218 591658 174454
rect 591102 173898 591338 174134
rect 591422 173898 591658 174134
rect 591102 138218 591338 138454
rect 591422 138218 591658 138454
rect 591102 137898 591338 138134
rect 591422 137898 591658 138134
rect 591102 102218 591338 102454
rect 591422 102218 591658 102454
rect 591102 101898 591338 102134
rect 591422 101898 591658 102134
rect 591102 66218 591338 66454
rect 591422 66218 591658 66454
rect 591102 65898 591338 66134
rect 591422 65898 591658 66134
rect 591102 30218 591338 30454
rect 591422 30218 591658 30454
rect 591102 29898 591338 30134
rect 591422 29898 591658 30134
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 682718 592298 682954
rect 592382 682718 592618 682954
rect 592062 682398 592298 682634
rect 592382 682398 592618 682634
rect 592062 646718 592298 646954
rect 592382 646718 592618 646954
rect 592062 646398 592298 646634
rect 592382 646398 592618 646634
rect 592062 610718 592298 610954
rect 592382 610718 592618 610954
rect 592062 610398 592298 610634
rect 592382 610398 592618 610634
rect 592062 574718 592298 574954
rect 592382 574718 592618 574954
rect 592062 574398 592298 574634
rect 592382 574398 592618 574634
rect 592062 538718 592298 538954
rect 592382 538718 592618 538954
rect 592062 538398 592298 538634
rect 592382 538398 592618 538634
rect 592062 502718 592298 502954
rect 592382 502718 592618 502954
rect 592062 502398 592298 502634
rect 592382 502398 592618 502634
rect 592062 466718 592298 466954
rect 592382 466718 592618 466954
rect 592062 466398 592298 466634
rect 592382 466398 592618 466634
rect 592062 430718 592298 430954
rect 592382 430718 592618 430954
rect 592062 430398 592298 430634
rect 592382 430398 592618 430634
rect 592062 394718 592298 394954
rect 592382 394718 592618 394954
rect 592062 394398 592298 394634
rect 592382 394398 592618 394634
rect 592062 358718 592298 358954
rect 592382 358718 592618 358954
rect 592062 358398 592298 358634
rect 592382 358398 592618 358634
rect 592062 322718 592298 322954
rect 592382 322718 592618 322954
rect 592062 322398 592298 322634
rect 592382 322398 592618 322634
rect 592062 286718 592298 286954
rect 592382 286718 592618 286954
rect 592062 286398 592298 286634
rect 592382 286398 592618 286634
rect 592062 250718 592298 250954
rect 592382 250718 592618 250954
rect 592062 250398 592298 250634
rect 592382 250398 592618 250634
rect 592062 214718 592298 214954
rect 592382 214718 592618 214954
rect 592062 214398 592298 214634
rect 592382 214398 592618 214634
rect 592062 178718 592298 178954
rect 592382 178718 592618 178954
rect 592062 178398 592298 178634
rect 592382 178398 592618 178634
rect 592062 142718 592298 142954
rect 592382 142718 592618 142954
rect 592062 142398 592298 142634
rect 592382 142398 592618 142634
rect 592062 106718 592298 106954
rect 592382 106718 592618 106954
rect 592062 106398 592298 106634
rect 592382 106398 592618 106634
rect 592062 70718 592298 70954
rect 592382 70718 592618 70954
rect 592062 70398 592298 70634
rect 592382 70398 592618 70634
rect 592062 34718 592298 34954
rect 592382 34718 592618 34954
rect 592062 34398 592298 34634
rect 592382 34398 592618 34634
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700954 592650 700986
rect -8726 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 592650 700954
rect -8726 700634 592650 700718
rect -8726 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 592650 700634
rect -8726 700366 592650 700398
rect -8726 696454 592650 696486
rect -8726 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 691954 592650 691986
rect -8726 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 592650 691954
rect -8726 691634 592650 691718
rect -8726 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 592650 691634
rect -8726 691366 592650 691398
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 682954 592650 682986
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect -8726 682634 592650 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect -8726 682366 592650 682398
rect -8726 678454 592650 678486
rect -8726 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 592650 678454
rect -8726 678134 592650 678218
rect -8726 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 592650 678134
rect -8726 677866 592650 677898
rect -8726 673954 592650 673986
rect -8726 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 592650 673954
rect -8726 673634 592650 673718
rect -8726 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 592650 673634
rect -8726 673366 592650 673398
rect -8726 669454 592650 669486
rect -8726 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 592650 669454
rect -8726 669134 592650 669218
rect -8726 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 592650 669134
rect -8726 668866 592650 668898
rect -8726 664954 592650 664986
rect -8726 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 592650 664954
rect -8726 664634 592650 664718
rect -8726 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 592650 664634
rect -8726 664366 592650 664398
rect -8726 660454 592650 660486
rect -8726 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 655954 592650 655986
rect -8726 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 592650 655954
rect -8726 655634 592650 655718
rect -8726 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 592650 655634
rect -8726 655366 592650 655398
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 646954 592650 646986
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect -8726 646634 592650 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect -8726 646366 592650 646398
rect -8726 642454 592650 642486
rect -8726 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 592650 642454
rect -8726 642134 592650 642218
rect -8726 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 592650 642134
rect -8726 641866 592650 641898
rect -8726 637954 592650 637986
rect -8726 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 592650 637954
rect -8726 637634 592650 637718
rect -8726 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 592650 637634
rect -8726 637366 592650 637398
rect -8726 633454 592650 633486
rect -8726 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 592650 633454
rect -8726 633134 592650 633218
rect -8726 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 592650 633134
rect -8726 632866 592650 632898
rect -8726 628954 592650 628986
rect -8726 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 592650 628954
rect -8726 628634 592650 628718
rect -8726 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 592650 628634
rect -8726 628366 592650 628398
rect -8726 624454 592650 624486
rect -8726 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 619954 592650 619986
rect -8726 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 592650 619954
rect -8726 619634 592650 619718
rect -8726 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 592650 619634
rect -8726 619366 592650 619398
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 610954 592650 610986
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect -8726 610634 592650 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect -8726 610366 592650 610398
rect -8726 606454 592650 606486
rect -8726 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 592650 606454
rect -8726 606134 592650 606218
rect -8726 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 592650 606134
rect -8726 605866 592650 605898
rect -8726 601954 592650 601986
rect -8726 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 592650 601954
rect -8726 601634 592650 601718
rect -8726 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 592650 601634
rect -8726 601366 592650 601398
rect -8726 597454 592650 597486
rect -8726 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 592650 597454
rect -8726 597134 592650 597218
rect -8726 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 592650 597134
rect -8726 596866 592650 596898
rect -8726 592954 592650 592986
rect -8726 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 592650 592954
rect -8726 592634 592650 592718
rect -8726 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 592650 592634
rect -8726 592366 592650 592398
rect -8726 588454 592650 588486
rect -8726 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 583954 592650 583986
rect -8726 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 592650 583954
rect -8726 583634 592650 583718
rect -8726 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 592650 583634
rect -8726 583366 592650 583398
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 574954 592650 574986
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect -8726 574634 592650 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect -8726 574366 592650 574398
rect -8726 570454 592650 570486
rect -8726 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 592650 570454
rect -8726 570134 592650 570218
rect -8726 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 592650 570134
rect -8726 569866 592650 569898
rect -8726 565954 592650 565986
rect -8726 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 592650 565954
rect -8726 565634 592650 565718
rect -8726 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 592650 565634
rect -8726 565366 592650 565398
rect -8726 561454 592650 561486
rect -8726 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 592650 561454
rect -8726 561134 592650 561218
rect -8726 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 592650 561134
rect -8726 560866 592650 560898
rect -8726 556954 592650 556986
rect -8726 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 592650 556954
rect -8726 556634 592650 556718
rect -8726 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 592650 556634
rect -8726 556366 592650 556398
rect -8726 552454 592650 552486
rect -8726 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 592650 552454
rect -8726 552134 592650 552218
rect -8726 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 547954 592650 547986
rect -8726 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 592650 547954
rect -8726 547634 592650 547718
rect -8726 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 592650 547634
rect -8726 547366 592650 547398
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 538954 592650 538986
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect -8726 538634 592650 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect -8726 538366 592650 538398
rect -8726 534454 592650 534486
rect -8726 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 529954 592650 529986
rect -8726 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 592650 529954
rect -8726 529634 592650 529718
rect -8726 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 592650 529634
rect -8726 529366 592650 529398
rect -8726 525454 592650 525486
rect -8726 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 592650 525454
rect -8726 525134 592650 525218
rect -8726 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 592650 525134
rect -8726 524866 592650 524898
rect -8726 520954 592650 520986
rect -8726 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 592650 520954
rect -8726 520634 592650 520718
rect -8726 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 592650 520634
rect -8726 520366 592650 520398
rect -8726 516454 592650 516486
rect -8726 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 511954 592650 511986
rect -8726 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 592650 511954
rect -8726 511634 592650 511718
rect -8726 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 592650 511634
rect -8726 511366 592650 511398
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 502954 592650 502986
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect -8726 502634 592650 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect -8726 502366 592650 502398
rect -8726 498454 592650 498486
rect -8726 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 592650 498454
rect -8726 498134 592650 498218
rect -8726 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 592650 498134
rect -8726 497866 592650 497898
rect -8726 493954 592650 493986
rect -8726 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 592650 493954
rect -8726 493634 592650 493718
rect -8726 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 592650 493634
rect -8726 493366 592650 493398
rect -8726 489454 592650 489486
rect -8726 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 592650 489454
rect -8726 489134 592650 489218
rect -8726 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 592650 489134
rect -8726 488866 592650 488898
rect -8726 484954 592650 484986
rect -8726 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 592650 484954
rect -8726 484634 592650 484718
rect -8726 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 592650 484634
rect -8726 484366 592650 484398
rect -8726 480454 592650 480486
rect -8726 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 475954 592650 475986
rect -8726 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 592650 475954
rect -8726 475634 592650 475718
rect -8726 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 592650 475634
rect -8726 475366 592650 475398
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 466954 592650 466986
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect -8726 466634 592650 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect -8726 466366 592650 466398
rect -8726 462454 592650 462486
rect -8726 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 592650 462454
rect -8726 462134 592650 462218
rect -8726 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 592650 462134
rect -8726 461866 592650 461898
rect -8726 457954 592650 457986
rect -8726 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 592650 457954
rect -8726 457634 592650 457718
rect -8726 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 592650 457634
rect -8726 457366 592650 457398
rect -8726 453454 592650 453486
rect -8726 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 592650 453454
rect -8726 453134 592650 453218
rect -8726 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 592650 453134
rect -8726 452866 592650 452898
rect -8726 448954 592650 448986
rect -8726 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 592650 448954
rect -8726 448634 592650 448718
rect -8726 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 592650 448634
rect -8726 448366 592650 448398
rect -8726 444454 592650 444486
rect -8726 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 439954 592650 439986
rect -8726 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 592650 439954
rect -8726 439634 592650 439718
rect -8726 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 592650 439634
rect -8726 439366 592650 439398
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 430954 592650 430986
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect -8726 430634 592650 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect -8726 430366 592650 430398
rect -8726 426454 592650 426486
rect -8726 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 592650 426454
rect -8726 426134 592650 426218
rect -8726 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 592650 426134
rect -8726 425866 592650 425898
rect -8726 421954 592650 421986
rect -8726 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 592650 421954
rect -8726 421634 592650 421718
rect -8726 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 592650 421634
rect -8726 421366 592650 421398
rect -8726 417454 592650 417486
rect -8726 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 592650 417454
rect -8726 417134 592650 417218
rect -8726 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 592650 417134
rect -8726 416866 592650 416898
rect -8726 412954 592650 412986
rect -8726 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 592650 412954
rect -8726 412634 592650 412718
rect -8726 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 592650 412634
rect -8726 412366 592650 412398
rect -8726 408454 592650 408486
rect -8726 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 403954 592650 403986
rect -8726 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 592650 403954
rect -8726 403634 592650 403718
rect -8726 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 592650 403634
rect -8726 403366 592650 403398
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 394954 592650 394986
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect -8726 394634 592650 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect -8726 394366 592650 394398
rect -8726 390454 592650 390486
rect -8726 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 592650 390454
rect -8726 390134 592650 390218
rect -8726 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 592650 390134
rect -8726 389866 592650 389898
rect -8726 385954 592650 385986
rect -8726 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 592650 385954
rect -8726 385634 592650 385718
rect -8726 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 592650 385634
rect -8726 385366 592650 385398
rect -8726 381454 592650 381486
rect -8726 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 592650 381454
rect -8726 381134 592650 381218
rect -8726 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 592650 381134
rect -8726 380866 592650 380898
rect -8726 376954 592650 376986
rect -8726 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 592650 376954
rect -8726 376634 592650 376718
rect -8726 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 592650 376634
rect -8726 376366 592650 376398
rect -8726 372454 592650 372486
rect -8726 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 367954 592650 367986
rect -8726 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 592650 367954
rect -8726 367634 592650 367718
rect -8726 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 592650 367634
rect -8726 367366 592650 367398
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 358954 592650 358986
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect -8726 358634 592650 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect -8726 358366 592650 358398
rect -8726 354454 592650 354486
rect -8726 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 349954 592650 349986
rect -8726 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 592650 349954
rect -8726 349634 592650 349718
rect -8726 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 592650 349634
rect -8726 349366 592650 349398
rect -8726 345454 592650 345486
rect -8726 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 592650 345454
rect -8726 345134 592650 345218
rect -8726 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 592650 345134
rect -8726 344866 592650 344898
rect -8726 340954 592650 340986
rect -8726 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 592650 340954
rect -8726 340634 592650 340718
rect -8726 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 592650 340634
rect -8726 340366 592650 340398
rect -8726 336454 592650 336486
rect -8726 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 331954 592650 331986
rect -8726 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 592650 331954
rect -8726 331634 592650 331718
rect -8726 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 592650 331634
rect -8726 331366 592650 331398
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 322954 592650 322986
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect -8726 322634 592650 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect -8726 322366 592650 322398
rect -8726 318454 592650 318486
rect -8726 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 592650 318454
rect -8726 318134 592650 318218
rect -8726 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 592650 318134
rect -8726 317866 592650 317898
rect -8726 313954 592650 313986
rect -8726 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 592650 313954
rect -8726 313634 592650 313718
rect -8726 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 592650 313634
rect -8726 313366 592650 313398
rect -8726 309454 592650 309486
rect -8726 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 592650 309454
rect -8726 309134 592650 309218
rect -8726 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 592650 309134
rect -8726 308866 592650 308898
rect -8726 304954 592650 304986
rect -8726 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 592650 304954
rect -8726 304634 592650 304718
rect -8726 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 592650 304634
rect -8726 304366 592650 304398
rect -8726 300454 592650 300486
rect -8726 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 295954 592650 295986
rect -8726 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 592650 295954
rect -8726 295634 592650 295718
rect -8726 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 592650 295634
rect -8726 295366 592650 295398
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 286954 592650 286986
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect -8726 286634 592650 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect -8726 286366 592650 286398
rect -8726 282454 592650 282486
rect -8726 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 592650 282454
rect -8726 282134 592650 282218
rect -8726 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 592650 282134
rect -8726 281866 592650 281898
rect -8726 277954 592650 277986
rect -8726 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 592650 277954
rect -8726 277634 592650 277718
rect -8726 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 592650 277634
rect -8726 277366 592650 277398
rect -8726 273454 592650 273486
rect -8726 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 592650 273454
rect -8726 273134 592650 273218
rect -8726 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 592650 273134
rect -8726 272866 592650 272898
rect -8726 268954 592650 268986
rect -8726 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 592650 268954
rect -8726 268634 592650 268718
rect -8726 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 592650 268634
rect -8726 268366 592650 268398
rect -8726 264454 592650 264486
rect -8726 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 259954 592650 259986
rect -8726 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 592650 259954
rect -8726 259634 592650 259718
rect -8726 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 592650 259634
rect -8726 259366 592650 259398
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 250954 592650 250986
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect -8726 250634 592650 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect -8726 250366 592650 250398
rect -8726 246454 592650 246486
rect -8726 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246303 424826 246454
rect 29382 246218 65342 246303
rect -8726 246134 65342 246218
rect -8726 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 246067 65342 246134
rect 65578 246067 65662 246303
rect 65898 246067 65982 246303
rect 66218 246067 66302 246303
rect 66538 246067 66622 246303
rect 66858 246067 66942 246303
rect 67178 246067 67262 246303
rect 67498 246067 67582 246303
rect 67818 246067 67902 246303
rect 68138 246067 68222 246303
rect 68458 246067 68542 246303
rect 68778 246067 68862 246303
rect 69098 246067 69182 246303
rect 69418 246067 69502 246303
rect 69738 246067 69822 246303
rect 70058 246218 424826 246303
rect 425062 246218 425146 246454
rect 425382 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 592650 246454
rect 70058 246134 592650 246218
rect 70058 246067 424826 246134
rect 29382 245898 424826 246067
rect 425062 245898 425146 246134
rect 425382 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 592650 246134
rect -8726 245866 592650 245898
rect -8726 241954 592650 241986
rect -8726 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241953 420326 241954
rect 24882 241718 65462 241953
rect -8726 241717 65462 241718
rect 65698 241717 65782 241953
rect 66018 241717 66102 241953
rect 66338 241717 66422 241953
rect 66658 241717 66742 241953
rect 66978 241717 67062 241953
rect 67298 241717 67382 241953
rect 67618 241717 67702 241953
rect 67938 241717 68022 241953
rect 68258 241717 68342 241953
rect 68578 241717 68662 241953
rect 68898 241717 68982 241953
rect 69218 241717 69302 241953
rect 69538 241717 69622 241953
rect 69858 241717 69942 241953
rect 70178 241717 70262 241953
rect 70498 241717 70582 241953
rect 70818 241717 70902 241953
rect 71138 241718 420326 241953
rect 420562 241718 420646 241954
rect 420882 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 592650 241954
rect 71138 241717 592650 241718
rect -8726 241634 592650 241717
rect -8726 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241633 420326 241634
rect 24882 241398 65462 241633
rect -8726 241397 65462 241398
rect 65698 241397 65782 241633
rect 66018 241397 66102 241633
rect 66338 241397 66422 241633
rect 66658 241397 66742 241633
rect 66978 241397 67062 241633
rect 67298 241397 67382 241633
rect 67618 241397 67702 241633
rect 67938 241397 68022 241633
rect 68258 241397 68342 241633
rect 68578 241397 68662 241633
rect 68898 241397 68982 241633
rect 69218 241397 69302 241633
rect 69538 241397 69622 241633
rect 69858 241397 69942 241633
rect 70178 241397 70262 241633
rect 70498 241397 70582 241633
rect 70818 241397 70902 241633
rect 71138 241398 420326 241633
rect 420562 241398 420646 241634
rect 420882 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 592650 241634
rect 71138 241397 592650 241398
rect -8726 241366 592650 241397
rect -8726 237454 592650 237486
rect -8726 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 592650 237454
rect -8726 237134 592650 237218
rect -8726 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 592650 237134
rect -8726 236866 592650 236898
rect -8726 232954 592650 232986
rect -8726 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 592650 232954
rect -8726 232634 592650 232718
rect -8726 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 592650 232634
rect -8726 232366 592650 232398
rect -8726 228454 592650 228486
rect -8726 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228453 406826 228454
rect 11382 228218 46826 228453
rect -8726 228217 46826 228218
rect 47062 228217 47146 228453
rect 47382 228217 82826 228453
rect 83062 228217 83146 228453
rect 83382 228217 118826 228453
rect 119062 228217 119146 228453
rect 119382 228217 190826 228453
rect 191062 228217 191146 228453
rect 191382 228217 226826 228453
rect 227062 228217 227146 228453
rect 227382 228217 262826 228453
rect 263062 228217 263146 228453
rect 263382 228217 298826 228453
rect 299062 228217 299146 228453
rect 299382 228217 334826 228453
rect 335062 228217 335146 228453
rect 335382 228217 370826 228453
rect 371062 228217 371146 228453
rect 371382 228218 406826 228453
rect 407062 228218 407146 228454
rect 407382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 592650 228454
rect 371382 228217 592650 228218
rect -8726 228134 592650 228217
rect -8726 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 228133 406826 228134
rect 11382 227898 46826 228133
rect -8726 227897 46826 227898
rect 47062 227897 47146 228133
rect 47382 227897 82826 228133
rect 83062 227897 83146 228133
rect 83382 227897 118826 228133
rect 119062 227897 119146 228133
rect 119382 227897 190826 228133
rect 191062 227897 191146 228133
rect 191382 227897 226826 228133
rect 227062 227897 227146 228133
rect 227382 227897 262826 228133
rect 263062 227897 263146 228133
rect 263382 227897 298826 228133
rect 299062 227897 299146 228133
rect 299382 227897 334826 228133
rect 335062 227897 335146 228133
rect 335382 227897 370826 228133
rect 371062 227897 371146 228133
rect 371382 227898 406826 228133
rect 407062 227898 407146 228134
rect 407382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 592650 228134
rect 371382 227897 592650 227898
rect -8726 227866 592650 227897
rect -8726 223954 592650 223986
rect -8726 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 592650 223954
rect -8726 223634 592650 223718
rect -8726 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 592650 223634
rect -8726 223366 592650 223398
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 214954 592650 214986
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect -8726 214634 592650 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect -8726 214366 592650 214398
rect -8726 210454 592650 210486
rect -8726 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 592650 210454
rect -8726 210134 592650 210218
rect -8726 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 592650 210134
rect -8726 209866 592650 209898
rect -8726 205954 592650 205986
rect -8726 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205861 204326 205954
rect 132882 205718 136036 205861
rect -8726 205634 136036 205718
rect -8726 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205625 136036 205634
rect 136272 205625 136356 205861
rect 136592 205625 136676 205861
rect 136912 205625 136996 205861
rect 137232 205625 137316 205861
rect 137552 205625 137636 205861
rect 137872 205625 137956 205861
rect 138192 205625 138276 205861
rect 138512 205625 138596 205861
rect 138832 205625 138916 205861
rect 139152 205625 139236 205861
rect 139472 205625 139556 205861
rect 139792 205625 139876 205861
rect 140112 205625 140196 205861
rect 140432 205625 140516 205861
rect 140752 205625 140836 205861
rect 141072 205625 141156 205861
rect 141392 205625 141476 205861
rect 141712 205625 141796 205861
rect 142032 205625 142116 205861
rect 142352 205625 142436 205861
rect 142672 205625 142756 205861
rect 142992 205625 143076 205861
rect 143312 205625 143396 205861
rect 143632 205625 143716 205861
rect 143952 205625 144036 205861
rect 144272 205625 144356 205861
rect 144592 205625 144676 205861
rect 144912 205625 144996 205861
rect 145232 205625 145316 205861
rect 145552 205625 145636 205861
rect 145872 205625 145956 205861
rect 146192 205625 146276 205861
rect 146512 205625 146596 205861
rect 146832 205625 146916 205861
rect 147152 205625 147236 205861
rect 147472 205625 147556 205861
rect 147792 205625 147876 205861
rect 148112 205625 148196 205861
rect 148432 205625 148516 205861
rect 148752 205625 148836 205861
rect 149072 205625 149156 205861
rect 149392 205625 149476 205861
rect 149712 205625 149796 205861
rect 150032 205625 150116 205861
rect 150352 205625 150436 205861
rect 150672 205625 150756 205861
rect 150992 205625 151076 205861
rect 151312 205625 151396 205861
rect 151632 205625 151716 205861
rect 151952 205625 152036 205861
rect 152272 205625 152356 205861
rect 152592 205625 152676 205861
rect 152912 205625 152996 205861
rect 153232 205625 153316 205861
rect 153552 205625 153636 205861
rect 153872 205625 153956 205861
rect 154192 205625 154276 205861
rect 154512 205625 154596 205861
rect 154832 205625 154916 205861
rect 155152 205625 155236 205861
rect 155472 205625 155556 205861
rect 155792 205625 155876 205861
rect 156112 205625 156196 205861
rect 156432 205625 156516 205861
rect 156752 205625 156836 205861
rect 157072 205625 157156 205861
rect 157392 205625 157476 205861
rect 157712 205625 157796 205861
rect 158032 205625 158116 205861
rect 158352 205625 158436 205861
rect 158672 205625 158756 205861
rect 158992 205625 159076 205861
rect 159312 205625 159396 205861
rect 159632 205625 159716 205861
rect 159952 205625 160036 205861
rect 160272 205625 160356 205861
rect 160592 205625 160676 205861
rect 160912 205625 160996 205861
rect 161232 205625 161316 205861
rect 161552 205625 161636 205861
rect 161872 205625 161956 205861
rect 162192 205625 162276 205861
rect 162512 205625 162596 205861
rect 162832 205625 162916 205861
rect 163152 205625 163236 205861
rect 163472 205625 163556 205861
rect 163792 205625 163876 205861
rect 164112 205625 164196 205861
rect 164432 205625 164516 205861
rect 164752 205625 164836 205861
rect 165072 205625 165156 205861
rect 165392 205718 204326 205861
rect 204562 205718 204646 205954
rect 204882 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 592650 205954
rect 165392 205634 592650 205718
rect 165392 205625 204326 205634
rect 132882 205398 204326 205625
rect 204562 205398 204646 205634
rect 204882 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 592650 205634
rect -8726 205366 592650 205398
rect -8726 201454 592650 201486
rect -8726 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201411 199826 201454
rect 128382 201218 137376 201411
rect -8726 201175 137376 201218
rect 137612 201175 137696 201411
rect 137932 201175 138016 201411
rect 138252 201175 138336 201411
rect 138572 201175 138656 201411
rect 138892 201175 138976 201411
rect 139212 201175 139296 201411
rect 139532 201175 139616 201411
rect 139852 201175 139936 201411
rect 140172 201175 140256 201411
rect 140492 201175 140576 201411
rect 140812 201175 140896 201411
rect 141132 201175 141216 201411
rect 141452 201175 141536 201411
rect 141772 201175 141856 201411
rect 142092 201175 142176 201411
rect 142412 201175 142496 201411
rect 142732 201175 142816 201411
rect 143052 201175 143136 201411
rect 143372 201175 143456 201411
rect 143692 201175 143776 201411
rect 144012 201175 144096 201411
rect 144332 201175 144416 201411
rect 144652 201175 144736 201411
rect 144972 201175 145056 201411
rect 145292 201175 145376 201411
rect 145612 201175 145696 201411
rect 145932 201175 146016 201411
rect 146252 201175 146336 201411
rect 146572 201175 146656 201411
rect 146892 201175 146976 201411
rect 147212 201175 147296 201411
rect 147532 201175 147616 201411
rect 147852 201175 147936 201411
rect 148172 201175 148256 201411
rect 148492 201175 148576 201411
rect 148812 201175 148896 201411
rect 149132 201175 149216 201411
rect 149452 201175 149536 201411
rect 149772 201175 149856 201411
rect 150092 201175 150176 201411
rect 150412 201175 150496 201411
rect 150732 201175 150816 201411
rect 151052 201175 151136 201411
rect 151372 201175 151456 201411
rect 151692 201175 151776 201411
rect 152012 201175 152096 201411
rect 152332 201175 152416 201411
rect 152652 201175 152736 201411
rect 152972 201175 153056 201411
rect 153292 201175 153376 201411
rect 153612 201175 153696 201411
rect 153932 201175 154016 201411
rect 154252 201175 154336 201411
rect 154572 201175 154656 201411
rect 154892 201175 154976 201411
rect 155212 201175 155296 201411
rect 155532 201175 155616 201411
rect 155852 201175 155936 201411
rect 156172 201175 156256 201411
rect 156492 201175 156576 201411
rect 156812 201175 156896 201411
rect 157132 201175 157216 201411
rect 157452 201175 157536 201411
rect 157772 201175 157856 201411
rect 158092 201175 158176 201411
rect 158412 201175 158496 201411
rect 158732 201175 158816 201411
rect 159052 201175 159136 201411
rect 159372 201175 159456 201411
rect 159692 201175 159776 201411
rect 160012 201175 160096 201411
rect 160332 201175 160416 201411
rect 160652 201175 160736 201411
rect 160972 201175 161056 201411
rect 161292 201175 161376 201411
rect 161612 201175 161696 201411
rect 161932 201175 162016 201411
rect 162252 201175 162336 201411
rect 162572 201175 162656 201411
rect 162892 201175 162976 201411
rect 163212 201175 163296 201411
rect 163532 201175 163616 201411
rect 163852 201175 163936 201411
rect 164172 201175 164256 201411
rect 164492 201175 164576 201411
rect 164812 201175 164896 201411
rect 165132 201175 165216 201411
rect 165452 201218 199826 201411
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 592650 201454
rect 165452 201175 592650 201218
rect -8726 201134 592650 201175
rect -8726 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 592650 201134
rect -8726 200866 592650 200898
rect -8726 196954 592650 196986
rect -8726 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 592650 196954
rect -8726 196634 592650 196718
rect -8726 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 592650 196634
rect -8726 196366 592650 196398
rect -8726 192454 592650 192486
rect -8726 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 187954 592650 187986
rect -8726 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 592650 187954
rect -8726 187634 592650 187718
rect -8726 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 592650 187634
rect -8726 187366 592650 187398
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 178954 592650 178986
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect -8726 178634 592650 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect -8726 178366 592650 178398
rect -8726 174454 592650 174486
rect -8726 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 137066 174454
rect 137302 174218 137386 174454
rect 137622 174218 137706 174454
rect 137942 174218 138026 174454
rect 138262 174218 138346 174454
rect 138582 174218 138666 174454
rect 138902 174218 138986 174454
rect 139222 174218 139306 174454
rect 139542 174218 139626 174454
rect 139862 174218 139946 174454
rect 140182 174218 140266 174454
rect 140502 174218 140586 174454
rect 140822 174218 140906 174454
rect 141142 174218 141226 174454
rect 141462 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 137066 174134
rect 137302 173898 137386 174134
rect 137622 173898 137706 174134
rect 137942 173898 138026 174134
rect 138262 173898 138346 174134
rect 138582 173898 138666 174134
rect 138902 173898 138986 174134
rect 139222 173898 139306 174134
rect 139542 173898 139626 174134
rect 139862 173898 139946 174134
rect 140182 173898 140266 174134
rect 140502 173898 140586 174134
rect 140822 173898 140906 174134
rect 141142 173898 141226 174134
rect 141462 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 169954 592650 169986
rect -8726 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 592650 169954
rect -8726 169634 592650 169718
rect -8726 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 592650 169634
rect -8726 169366 592650 169398
rect -8726 165454 592650 165486
rect -8726 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 592650 165454
rect -8726 165134 592650 165218
rect -8726 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 592650 165134
rect -8726 164866 592650 164898
rect -8726 160954 592650 160986
rect -8726 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 592650 160954
rect -8726 160634 592650 160718
rect -8726 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 592650 160634
rect -8726 160366 592650 160398
rect -8726 156454 592650 156486
rect -8726 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 151954 592650 151986
rect -8726 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 592650 151954
rect -8726 151634 592650 151718
rect -8726 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 592650 151634
rect -8726 151366 592650 151398
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 142954 592650 142986
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect -8726 142634 592650 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect -8726 142366 592650 142398
rect -8726 138454 592650 138486
rect -8726 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 592650 138454
rect -8726 138134 592650 138218
rect -8726 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 592650 138134
rect -8726 137866 592650 137898
rect -8726 133954 592650 133986
rect -8726 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 592650 133954
rect -8726 133634 592650 133718
rect -8726 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 592650 133634
rect -8726 133366 592650 133398
rect -8726 129454 592650 129486
rect -8726 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 592650 129454
rect -8726 129134 592650 129218
rect -8726 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 592650 129134
rect -8726 128866 592650 128898
rect -8726 124954 592650 124986
rect -8726 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 592650 124954
rect -8726 124634 592650 124718
rect -8726 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 592650 124634
rect -8726 124366 592650 124398
rect -8726 120454 592650 120486
rect -8726 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 115954 592650 115986
rect -8726 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 139610 115954
rect 139846 115718 170330 115954
rect 170566 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 592650 115954
rect -8726 115634 592650 115718
rect -8726 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 139610 115634
rect 139846 115398 170330 115634
rect 170566 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 592650 115634
rect -8726 115366 592650 115398
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 124250 111454
rect 124486 111218 154970 111454
rect 155206 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 124250 111134
rect 124486 110898 154970 111134
rect 155206 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 106954 592650 106986
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect -8726 106634 592650 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect -8726 106366 592650 106398
rect -8726 102454 592650 102486
rect -8726 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 592650 102454
rect -8726 102134 592650 102218
rect -8726 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 592650 102134
rect -8726 101866 592650 101898
rect -8726 97954 592650 97986
rect -8726 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 592650 97954
rect -8726 97634 592650 97718
rect -8726 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 592650 97634
rect -8726 97366 592650 97398
rect -8726 93454 592650 93486
rect -8726 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 592650 93454
rect -8726 93134 592650 93218
rect -8726 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 592650 93134
rect -8726 92866 592650 92898
rect -8726 88954 592650 88986
rect -8726 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 592650 88954
rect -8726 88634 592650 88718
rect -8726 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 592650 88634
rect -8726 88366 592650 88398
rect -8726 84454 592650 84486
rect -8726 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 79954 592650 79986
rect -8726 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 592650 79954
rect -8726 79634 592650 79718
rect -8726 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 592650 79634
rect -8726 79366 592650 79398
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 70954 592650 70986
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect -8726 70634 592650 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect -8726 70366 592650 70398
rect -8726 66454 592650 66486
rect -8726 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 592650 66454
rect -8726 66134 592650 66218
rect -8726 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 592650 66134
rect -8726 65866 592650 65898
rect -8726 61954 592650 61986
rect -8726 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 592650 61954
rect -8726 61634 592650 61718
rect -8726 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 592650 61634
rect -8726 61366 592650 61398
rect -8726 57454 592650 57486
rect -8726 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 592650 57454
rect -8726 57134 592650 57218
rect -8726 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 592650 57134
rect -8726 56866 592650 56898
rect -8726 52954 592650 52986
rect -8726 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 592650 52954
rect -8726 52634 592650 52718
rect -8726 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 592650 52634
rect -8726 52366 592650 52398
rect -8726 48454 592650 48486
rect -8726 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 43954 592650 43986
rect -8726 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 592650 43954
rect -8726 43634 592650 43718
rect -8726 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 592650 43634
rect -8726 43366 592650 43398
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 34954 592650 34986
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect -8726 34634 592650 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect -8726 34366 592650 34398
rect -8726 30454 592650 30486
rect -8726 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 592650 30454
rect -8726 30134 592650 30218
rect -8726 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 592650 30134
rect -8726 29866 592650 29898
rect -8726 25954 592650 25986
rect -8726 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 592650 25954
rect -8726 25634 592650 25718
rect -8726 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 592650 25634
rect -8726 25366 592650 25398
rect -8726 21454 592650 21486
rect -8726 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 592650 21454
rect -8726 21134 592650 21218
rect -8726 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 592650 21134
rect -8726 20866 592650 20898
rect -8726 16954 592650 16986
rect -8726 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 592650 16954
rect -8726 16634 592650 16718
rect -8726 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 592650 16634
rect -8726 16366 592650 16398
rect -8726 12454 592650 12486
rect -8726 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 592650 12134
rect -8726 11866 592650 11898
rect -8726 7954 592650 7986
rect -8726 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 592650 7954
rect -8726 7634 592650 7718
rect -8726 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 592650 7634
rect -8726 7366 592650 7398
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use PD_M1_M2  PD_M1_M2_macro0
timestamp 0
transform 1 0 16000 0 1 232484
box 30000 -2000 380500 14200
use rlbp_macro  rlbp_macro0
timestamp 0
transform 1 0 120000 0 1 80000
box 0 0 60000 60000
use SystemLevel  sl_macro0
timestamp 0
transform 1 0 148914 0 1 188300
box -13000 -15200 17500 18000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 248684 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 248684 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 78000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 248684 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 78000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 142000 182414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 248684 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 248684 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 248684 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 248684 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 248684 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 248684 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 248684 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 10794 -7654 11414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 -7654 47414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 248684 47414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 -7654 83414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 248684 83414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 -7654 119414 78000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 142000 119414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 248684 119414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 -7654 155414 78000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 248684 155414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 -7654 191414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 248684 191414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 -7654 227414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 248684 227414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 -7654 263414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 248684 263414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 -7654 299414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 248684 299414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 -7654 335414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 248684 335414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 -7654 371414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 248684 371414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 -7654 407414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 -7654 443414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 -7654 479414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 -7654 515414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 550794 -7654 551414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 11866 592650 12486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 47866 592650 48486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 83866 592650 84486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 119866 592650 120486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 155866 592650 156486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 191866 592650 192486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 227866 592650 228486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 263866 592650 264486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 299866 592650 300486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 335866 592650 336486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 371866 592650 372486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 407866 592650 408486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 443866 592650 444486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 479866 592650 480486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 515866 592650 516486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 551866 592650 552486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 587866 592650 588486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 623866 592650 624486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 659866 592650 660486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 695866 592650 696486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 19794 -7654 20414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 -7654 56414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 248684 56414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 -7654 92414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 248684 92414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 -7654 128414 78000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 142000 128414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 248684 128414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 -7654 164414 78000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 248684 164414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 -7654 200414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 248684 200414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 -7654 236414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 248684 236414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 -7654 272414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 248684 272414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 -7654 308414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 248684 308414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 -7654 344414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 248684 344414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 -7654 380414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 248684 380414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 -7654 416414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 451794 -7654 452414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 -7654 488414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 523794 -7654 524414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 559794 -7654 560414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 20866 592650 21486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 56866 592650 57486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 92866 592650 93486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 128866 592650 129486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 164866 592650 165486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 200866 592650 201486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 236866 592650 237486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 272866 592650 273486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 308866 592650 309486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 344866 592650 345486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 380866 592650 381486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 416866 592650 417486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 452866 592650 453486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 488866 592650 489486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 524866 592650 525486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 560866 592650 561486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 596866 592650 597486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 632866 592650 633486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 668866 592650 669486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 28794 -7654 29414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 -7654 65414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 248684 65414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 -7654 101414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 248684 101414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 -7654 137414 78000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 248684 137414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 -7654 173414 78000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 142000 173414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 248684 173414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 -7654 209414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 248684 209414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 -7654 245414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 248684 245414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 -7654 281414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 248684 281414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 -7654 317414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 248684 317414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 -7654 353414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 248684 353414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 -7654 389414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 248684 389414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 424794 -7654 425414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 460794 -7654 461414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 496794 -7654 497414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 532794 -7654 533414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 568794 -7654 569414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 29866 592650 30486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 65866 592650 66486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 101866 592650 102486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 137866 592650 138486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 173866 592650 174486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 209866 592650 210486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 245866 592650 246486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 281866 592650 282486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 317866 592650 318486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 353866 592650 354486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 389866 592650 390486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 425866 592650 426486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 461866 592650 462486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 497866 592650 498486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 533866 592650 534486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 569866 592650 570486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 605866 592650 606486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 641866 592650 642486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 677866 592650 678486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 24294 -7654 24914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 -7654 60914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 248684 60914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 -7654 96914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 248684 96914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 -7654 132914 78000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 142000 132914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 248684 132914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 -7654 168914 78000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 248684 168914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 -7654 204914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 248684 204914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 -7654 240914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 248684 240914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 -7654 276914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 248684 276914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 -7654 312914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 248684 312914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 -7654 348914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 248684 348914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 -7654 384914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 248684 384914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 -7654 420914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 456294 -7654 456914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 492294 -7654 492914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 528294 -7654 528914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 564294 -7654 564914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 25366 592650 25986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 61366 592650 61986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 97366 592650 97986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 133366 592650 133986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 169366 592650 169986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 205366 592650 205986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 241366 592650 241986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 277366 592650 277986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 313366 592650 313986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 349366 592650 349986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 385366 592650 385986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 421366 592650 421986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 457366 592650 457986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 493366 592650 493986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 529366 592650 529986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 565366 592650 565986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 601366 592650 601986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 637366 592650 637986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 673366 592650 673986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 33294 -7654 33914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 -7654 69914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 248684 69914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 -7654 105914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 248684 105914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 -7654 141914 78000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 248684 141914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 -7654 177914 78000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 142000 177914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 248684 177914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 -7654 213914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 248684 213914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 -7654 249914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 248684 249914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 -7654 285914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 248684 285914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 -7654 321914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 248684 321914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 -7654 357914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 248684 357914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 -7654 393914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 248684 393914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 -7654 429914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 465294 -7654 465914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 -7654 501914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 537294 -7654 537914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 573294 -7654 573914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 34366 592650 34986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 70366 592650 70986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 106366 592650 106986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 142366 592650 142986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 178366 592650 178986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 214366 592650 214986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 250366 592650 250986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 286366 592650 286986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 322366 592650 322986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 358366 592650 358986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 394366 592650 394986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 430366 592650 430986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 466366 592650 466986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 502366 592650 502986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 538366 592650 538986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 574366 592650 574986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 610366 592650 610986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 646366 592650 646986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 682366 592650 682986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 6294 -7654 6914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 42294 -7654 42914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 -7654 78914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 248684 78914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 -7654 114914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 248684 114914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 -7654 150914 78000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 248684 150914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 -7654 186914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 248684 186914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 -7654 222914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 248684 222914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 -7654 258914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 248684 258914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 -7654 294914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 248684 294914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 -7654 330914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 248684 330914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 -7654 366914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 248684 366914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 -7654 402914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 -7654 438914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 -7654 474914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 -7654 510914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 546294 -7654 546914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 582294 -7654 582914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 7366 592650 7986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 43366 592650 43986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 79366 592650 79986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 115366 592650 115986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 151366 592650 151986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 187366 592650 187986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 223366 592650 223986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 259366 592650 259986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 295366 592650 295986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 331366 592650 331986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 367366 592650 367986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 403366 592650 403986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 439366 592650 439986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 475366 592650 475986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 511366 592650 511986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 547366 592650 547986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 583366 592650 583986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 619366 592650 619986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 655366 592650 655986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 691366 592650 691986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 15294 -7654 15914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 -7654 51914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 248684 51914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 -7654 87914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 248684 87914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 -7654 123914 78000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 142000 123914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 248684 123914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 -7654 159914 78000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 248684 159914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 -7654 195914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 248684 195914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 -7654 231914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 248684 231914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 -7654 267914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 248684 267914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 -7654 303914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 248684 303914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 -7654 339914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 248684 339914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 -7654 375914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 248684 375914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 -7654 411914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 -7654 447914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 -7654 483914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 -7654 519914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 555294 -7654 555914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 16366 592650 16986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 52366 592650 52986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 88366 592650 88986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 124366 592650 124986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 160366 592650 160986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 196366 592650 196986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 232366 592650 232986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 268366 592650 268986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 304366 592650 304986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 340366 592650 340986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 376366 592650 376986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 412366 592650 412986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 448366 592650 448986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 484366 592650 484986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 520366 592650 520986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 556366 592650 556986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 592366 592650 592986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 628366 592650 628986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 664366 592650 664986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 700366 592650 700986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
