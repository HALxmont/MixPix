VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO PD1
  CLASS BLOCK ;
  FOREIGN PD1 ;
  ORIGIN -145.000 10.000 ;
  SIZE 1760.000 BY 105.000 ;
  PIN PD1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.640000 ;
    PORT
      LAYER nwell ;
        RECT 199.300 17.300 200.700 18.700 ;
      LAYER li1 ;
        RECT 199.500 17.500 200.500 18.500 ;
        RECT 199.750 6.150 200.250 17.500 ;
        RECT 199.750 5.650 205.400 6.150 ;
        RECT 204.900 1.500 205.400 5.650 ;
      LAYER met1 ;
        RECT 204.840 1.470 205.460 2.030 ;
        RECT 204.900 -6.280 205.400 1.470 ;
      LAYER via ;
        RECT 204.900 -6.250 205.400 -5.750 ;
      LAYER met2 ;
        RECT 202.500 -10.000 208.750 -5.000 ;
    END
  END PD1
  PIN PD2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.640000 ;
    PORT
      LAYER nwell ;
        RECT 349.300 17.300 350.700 18.700 ;
      LAYER li1 ;
        RECT 349.600 17.600 350.400 18.400 ;
        RECT 349.675 8.825 350.325 17.600 ;
        RECT 349.675 8.175 354.650 8.825 ;
        RECT 354.000 2.375 354.650 8.175 ;
      LAYER mcon ;
        RECT 354.030 2.405 354.620 2.995 ;
      LAYER met1 ;
        RECT 354.000 -2.250 354.650 3.055 ;
        RECT 355.250 -2.250 355.750 -2.220 ;
        RECT 354.000 -2.750 355.750 -2.250 ;
        RECT 355.250 -2.780 355.750 -2.750 ;
      LAYER via ;
        RECT 355.250 -2.750 355.750 -2.250 ;
      LAYER met2 ;
        RECT 355.220 -2.750 355.780 -2.250 ;
        RECT 355.250 -4.500 355.750 -2.750 ;
        RECT 355.000 -5.000 356.000 -4.500 ;
        RECT 352.500 -10.000 358.750 -5.000 ;
    END
  END PD2
  PIN PD3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.640000 ;
    PORT
      LAYER nwell ;
        RECT 499.300 17.300 500.700 18.700 ;
      LAYER li1 ;
        RECT 499.600 17.600 500.400 18.400 ;
        RECT 499.800 4.150 500.200 17.600 ;
        RECT 499.800 3.750 504.450 4.150 ;
      LAYER mcon ;
        RECT 504.050 3.750 504.450 4.150 ;
      LAYER met1 ;
        RECT 503.990 3.720 504.510 4.180 ;
        RECT 504.050 0.000 504.450 3.720 ;
        RECT 504.000 -1.750 504.450 0.000 ;
        RECT 505.250 -1.750 505.750 -1.720 ;
        RECT 504.000 -2.250 505.750 -1.750 ;
        RECT 505.250 -2.280 505.750 -2.250 ;
      LAYER via ;
        RECT 505.250 -2.250 505.750 -1.750 ;
      LAYER met2 ;
        RECT 505.220 -2.250 505.780 -1.750 ;
        RECT 505.250 -4.500 505.750 -2.250 ;
        RECT 505.000 -5.000 506.000 -4.500 ;
        RECT 502.500 -10.000 508.750 -5.000 ;
    END
  END PD3
  PIN PD4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.640000 ;
    PORT
      LAYER nwell ;
        RECT 649.300 17.300 650.700 18.700 ;
      LAYER li1 ;
        RECT 649.600 17.600 650.400 18.400 ;
        RECT 649.800 3.750 650.200 17.600 ;
      LAYER met1 ;
        RECT 649.740 4.150 650.260 4.180 ;
        RECT 649.740 3.750 654.450 4.150 ;
        RECT 649.740 3.720 650.260 3.750 ;
        RECT 654.050 0.000 654.450 3.750 ;
        RECT 654.000 -0.500 654.450 0.000 ;
        RECT 654.000 -1.000 655.750 -0.500 ;
        RECT 655.250 -4.030 655.750 -1.000 ;
      LAYER via ;
        RECT 655.250 -4.000 655.750 -3.500 ;
      LAYER met2 ;
        RECT 655.220 -4.000 655.780 -3.500 ;
        RECT 655.250 -4.500 655.750 -4.000 ;
        RECT 655.000 -5.000 656.000 -4.500 ;
        RECT 652.500 -10.000 658.750 -5.000 ;
    END
  END PD4
  PIN PD5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.640000 ;
    PORT
      LAYER nwell ;
        RECT 799.300 17.300 800.700 18.700 ;
      LAYER li1 ;
        RECT 799.600 17.600 800.400 18.400 ;
        RECT 799.800 4.400 800.200 17.600 ;
        RECT 799.800 4.000 805.700 4.400 ;
        RECT 805.300 2.600 805.700 4.000 ;
      LAYER met1 ;
        RECT 805.240 2.570 805.760 3.030 ;
        RECT 805.300 -0.450 805.700 2.570 ;
        RECT 805.200 -0.600 805.800 -0.450 ;
        RECT 805.250 -1.030 805.750 -0.600 ;
      LAYER via ;
        RECT 805.250 -1.000 805.750 -0.500 ;
      LAYER met2 ;
        RECT 805.220 -1.000 805.780 -0.500 ;
        RECT 805.250 -4.500 805.750 -1.000 ;
        RECT 805.000 -5.000 806.000 -4.500 ;
        RECT 802.500 -10.000 808.750 -5.000 ;
    END
  END PD5
  PIN PD6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.640000 ;
    PORT
      LAYER nwell ;
        RECT 949.300 17.300 950.700 18.700 ;
      LAYER li1 ;
        RECT 949.600 17.600 950.400 18.400 ;
        RECT 949.800 4.200 950.200 17.600 ;
        RECT 949.800 3.800 955.700 4.200 ;
        RECT 955.300 2.500 955.700 3.800 ;
      LAYER met1 ;
        RECT 955.240 2.470 955.760 2.930 ;
        RECT 955.300 -0.450 955.700 2.470 ;
        RECT 955.200 -0.600 955.800 -0.450 ;
        RECT 955.250 -1.030 955.750 -0.600 ;
      LAYER via ;
        RECT 955.250 -1.000 955.750 -0.500 ;
      LAYER met2 ;
        RECT 955.220 -1.000 955.780 -0.500 ;
        RECT 955.250 -4.500 955.750 -1.000 ;
        RECT 955.000 -5.000 956.000 -4.500 ;
        RECT 952.500 -10.000 958.750 -5.000 ;
    END
  END PD6
  PIN PD7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.640000 ;
    PORT
      LAYER nwell ;
        RECT 1099.300 17.300 1100.700 18.700 ;
      LAYER li1 ;
        RECT 1099.600 17.600 1100.400 18.400 ;
        RECT 1099.800 4.200 1100.200 17.600 ;
        RECT 1099.800 3.800 1105.700 4.200 ;
        RECT 1105.300 2.350 1105.700 3.800 ;
      LAYER met1 ;
        RECT 1105.240 2.320 1105.760 2.780 ;
        RECT 1105.300 -0.450 1105.700 2.320 ;
        RECT 1105.200 -1.050 1105.800 -0.450 ;
      LAYER via ;
        RECT 1105.250 -1.000 1105.750 -0.500 ;
      LAYER met2 ;
        RECT 1105.250 -4.500 1105.750 -0.470 ;
        RECT 1105.000 -5.000 1106.000 -4.500 ;
        RECT 1102.500 -10.000 1108.750 -5.000 ;
    END
  END PD7
  PIN PD8
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.640000 ;
    PORT
      LAYER nwell ;
        RECT 1249.300 17.300 1250.700 18.700 ;
      LAYER li1 ;
        RECT 1249.600 17.600 1250.400 18.400 ;
        RECT 1249.800 4.100 1250.200 17.600 ;
        RECT 1249.800 3.700 1255.650 4.100 ;
        RECT 1255.250 2.000 1255.650 3.700 ;
      LAYER met1 ;
        RECT 1255.190 1.970 1255.710 2.430 ;
        RECT 1255.250 -0.450 1255.650 1.970 ;
        RECT 1255.200 -1.050 1255.800 -0.450 ;
      LAYER via ;
        RECT 1255.250 -1.000 1255.750 -0.500 ;
      LAYER met2 ;
        RECT 1255.250 -4.500 1255.750 -0.470 ;
        RECT 1255.000 -5.000 1256.000 -4.500 ;
        RECT 1252.500 -10.000 1258.750 -5.000 ;
    END
  END PD8
  PIN PD9
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.640000 ;
    PORT
      LAYER nwell ;
        RECT 1399.300 17.300 1400.700 18.700 ;
      LAYER li1 ;
        RECT 1399.600 17.600 1400.400 18.400 ;
        RECT 1399.800 4.100 1400.200 17.600 ;
        RECT 1399.800 3.700 1405.650 4.100 ;
        RECT 1405.250 2.000 1405.650 3.700 ;
      LAYER met1 ;
        RECT 1405.190 1.970 1405.710 2.430 ;
        RECT 1405.250 -0.450 1405.650 1.970 ;
        RECT 1405.200 -1.050 1405.800 -0.450 ;
      LAYER via ;
        RECT 1405.250 -1.000 1405.750 -0.500 ;
      LAYER met2 ;
        RECT 1405.250 -4.500 1405.750 -0.470 ;
        RECT 1405.000 -5.000 1406.000 -4.500 ;
        RECT 1402.500 -10.000 1408.750 -5.000 ;
    END
  END PD9
  PIN PD10
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.640000 ;
    PORT
      LAYER nwell ;
        RECT 1549.300 17.300 1550.700 18.700 ;
      LAYER li1 ;
        RECT 1549.600 17.600 1550.400 18.400 ;
        RECT 1549.800 4.100 1550.200 17.600 ;
        RECT 1549.800 3.700 1555.650 4.100 ;
        RECT 1555.250 2.000 1555.650 3.700 ;
      LAYER met1 ;
        RECT 1555.190 1.970 1555.710 2.430 ;
        RECT 1555.250 -0.450 1555.650 1.970 ;
        RECT 1555.200 -1.050 1555.800 -0.450 ;
      LAYER via ;
        RECT 1555.250 -1.000 1555.750 -0.500 ;
      LAYER met2 ;
        RECT 1555.250 -4.500 1555.750 -0.470 ;
        RECT 1555.000 -5.000 1556.000 -4.500 ;
        RECT 1552.500 -10.000 1558.750 -5.000 ;
    END
  END PD10
  PIN PD11
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.640000 ;
    PORT
      LAYER nwell ;
        RECT 1699.300 17.300 1700.700 18.700 ;
      LAYER li1 ;
        RECT 1699.600 17.600 1700.400 18.400 ;
        RECT 1699.800 4.100 1700.200 17.600 ;
        RECT 1699.800 3.700 1705.650 4.100 ;
        RECT 1705.250 2.000 1705.650 3.700 ;
      LAYER met1 ;
        RECT 1705.190 1.970 1705.710 2.430 ;
        RECT 1705.250 -0.450 1705.650 1.970 ;
        RECT 1705.200 -1.050 1705.800 -0.450 ;
      LAYER via ;
        RECT 1705.250 -1.000 1705.750 -0.500 ;
      LAYER met2 ;
        RECT 1705.250 -4.500 1705.750 -0.470 ;
        RECT 1705.000 -5.000 1706.000 -4.500 ;
        RECT 1702.500 -10.000 1708.750 -5.000 ;
    END
  END PD11
  PIN PD12
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.640000 ;
    PORT
      LAYER nwell ;
        RECT 1849.300 17.300 1850.700 18.700 ;
      LAYER li1 ;
        RECT 1849.600 17.600 1850.400 18.400 ;
        RECT 1849.800 4.100 1850.200 17.600 ;
        RECT 1849.800 3.700 1855.650 4.100 ;
        RECT 1855.250 2.000 1855.650 3.700 ;
      LAYER met1 ;
        RECT 1855.190 1.970 1855.710 2.430 ;
        RECT 1855.250 -0.450 1855.650 1.970 ;
        RECT 1855.200 -1.050 1855.800 -0.450 ;
      LAYER via ;
        RECT 1855.250 -1.000 1855.750 -0.500 ;
      LAYER met2 ;
        RECT 1855.250 -4.500 1855.750 -0.470 ;
        RECT 1855.000 -5.000 1856.000 -4.500 ;
        RECT 1852.500 -10.000 1858.750 -5.000 ;
    END
  END PD12
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 246.500 67.000 270.500 71.000 ;
        RECT 246.500 63.000 270.470 67.000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 150.000 33.500 251.500 35.000 ;
        RECT 150.000 1.500 151.500 33.500 ;
        RECT 250.000 1.500 251.500 33.500 ;
        RECT 150.000 0.000 251.500 1.500 ;
        RECT 300.000 33.500 401.500 35.000 ;
        RECT 300.000 1.500 301.500 33.500 ;
        RECT 400.000 1.500 401.500 33.500 ;
        RECT 300.000 0.000 401.500 1.500 ;
        RECT 450.000 33.500 551.500 35.000 ;
        RECT 450.000 1.500 451.500 33.500 ;
        RECT 550.000 1.500 551.500 33.500 ;
        RECT 450.000 0.000 551.500 1.500 ;
        RECT 600.000 33.500 701.500 35.000 ;
        RECT 600.000 1.500 601.500 33.500 ;
        RECT 700.000 1.500 701.500 33.500 ;
        RECT 600.000 0.000 701.500 1.500 ;
        RECT 750.000 33.500 851.500 35.000 ;
        RECT 750.000 1.500 751.500 33.500 ;
        RECT 850.000 1.500 851.500 33.500 ;
        RECT 750.000 0.000 851.500 1.500 ;
        RECT 900.000 33.500 1001.500 35.000 ;
        RECT 900.000 1.500 901.500 33.500 ;
        RECT 1000.000 1.500 1001.500 33.500 ;
        RECT 900.000 0.000 1001.500 1.500 ;
        RECT 1050.000 33.500 1151.500 35.000 ;
        RECT 1050.000 1.500 1051.500 33.500 ;
        RECT 1150.000 1.500 1151.500 33.500 ;
        RECT 1050.000 0.000 1151.500 1.500 ;
        RECT 1200.000 33.500 1301.500 35.000 ;
        RECT 1200.000 1.500 1201.500 33.500 ;
        RECT 1300.000 1.500 1301.500 33.500 ;
        RECT 1200.000 0.000 1301.500 1.500 ;
        RECT 1350.000 33.500 1451.500 35.000 ;
        RECT 1350.000 1.500 1351.500 33.500 ;
        RECT 1450.000 1.500 1451.500 33.500 ;
        RECT 1350.000 0.000 1451.500 1.500 ;
        RECT 1500.000 33.500 1601.500 35.000 ;
        RECT 1500.000 1.500 1501.500 33.500 ;
        RECT 1600.000 1.500 1601.500 33.500 ;
        RECT 1500.000 0.000 1601.500 1.500 ;
        RECT 1650.000 33.500 1751.500 35.000 ;
        RECT 1650.000 1.500 1651.500 33.500 ;
        RECT 1750.000 1.500 1751.500 33.500 ;
        RECT 1650.000 0.000 1751.500 1.500 ;
        RECT 1800.000 33.500 1901.500 35.000 ;
        RECT 1800.000 1.500 1801.500 33.500 ;
        RECT 1900.000 1.500 1901.500 33.500 ;
        RECT 1800.000 0.000 1901.500 1.500 ;
      LAYER li1 ;
        RECT 286.000 38.000 290.000 93.000 ;
        RECT 150.500 34.000 1902.500 38.000 ;
        RECT 150.500 1.000 151.000 34.000 ;
        RECT 250.500 1.000 251.000 34.000 ;
        RECT 150.500 0.500 251.000 1.000 ;
        RECT 300.500 1.000 301.000 34.000 ;
        RECT 400.500 1.000 401.000 34.000 ;
        RECT 300.500 0.500 401.000 1.000 ;
        RECT 450.500 1.000 451.000 34.000 ;
        RECT 550.500 1.000 551.000 34.000 ;
        RECT 450.500 0.500 551.000 1.000 ;
        RECT 600.500 1.000 601.000 34.000 ;
        RECT 700.500 1.000 701.000 34.000 ;
        RECT 600.500 0.500 701.000 1.000 ;
        RECT 750.500 1.000 751.000 34.000 ;
        RECT 850.500 1.000 851.000 34.000 ;
        RECT 750.500 0.500 851.000 1.000 ;
        RECT 900.500 1.000 901.000 34.000 ;
        RECT 1000.500 1.000 1001.000 34.000 ;
        RECT 900.500 0.500 1001.000 1.000 ;
        RECT 1050.500 1.000 1051.000 34.000 ;
        RECT 1150.500 1.000 1151.000 34.000 ;
        RECT 1050.500 0.500 1151.000 1.000 ;
        RECT 1200.500 1.000 1201.000 34.000 ;
        RECT 1300.500 1.000 1301.000 34.000 ;
        RECT 1200.500 0.500 1301.000 1.000 ;
        RECT 1350.500 1.000 1351.000 34.000 ;
        RECT 1450.500 1.000 1451.000 34.000 ;
        RECT 1350.500 0.500 1451.000 1.000 ;
        RECT 1500.500 1.000 1501.000 34.000 ;
        RECT 1600.500 1.000 1601.000 34.000 ;
        RECT 1500.500 0.500 1601.000 1.000 ;
        RECT 1650.500 1.000 1651.000 34.000 ;
        RECT 1750.500 1.000 1751.000 34.000 ;
        RECT 1650.500 0.500 1751.000 1.000 ;
        RECT 1800.500 1.000 1801.000 34.000 ;
        RECT 1900.500 1.000 1901.000 34.000 ;
        RECT 1800.500 0.500 1901.000 1.000 ;
      LAYER mcon ;
        RECT 286.000 89.000 290.000 93.000 ;
      LAYER met1 ;
        RECT 285.940 93.000 290.060 93.030 ;
        RECT 282.970 89.000 290.060 93.000 ;
        RECT 285.940 88.970 290.060 89.000 ;
      LAYER via ;
        RECT 283.000 89.000 287.000 93.000 ;
      LAYER met2 ;
        RECT 283.000 93.000 287.000 93.030 ;
        RECT 279.955 89.000 287.000 93.000 ;
        RECT 283.000 88.970 287.000 89.000 ;
      LAYER via2 ;
        RECT 280.000 89.000 284.000 93.000 ;
      LAYER met3 ;
        RECT 279.945 88.975 284.025 93.025 ;
      LAYER via3 ;
        RECT 279.975 88.975 283.975 93.025 ;
      LAYER met4 ;
        RECT 251.000 89.000 295.000 95.000 ;
        RECT 279.970 88.970 283.980 89.000 ;
    END
  END VSS
  OBS
      LAYER nwell ;
        RECT 151.500 30.500 250.000 33.500 ;
        RECT 151.500 4.500 154.500 30.500 ;
        RECT 185.500 25.000 215.500 27.500 ;
        RECT 185.500 10.000 188.000 25.000 ;
        RECT 213.000 10.000 215.500 25.000 ;
        RECT 185.500 7.500 215.500 10.000 ;
        RECT 247.000 4.500 250.000 30.500 ;
        RECT 151.500 1.500 250.000 4.500 ;
        RECT 301.500 30.500 400.000 33.500 ;
        RECT 301.500 4.500 304.500 30.500 ;
        RECT 335.500 25.000 365.500 27.500 ;
        RECT 335.500 10.000 338.000 25.000 ;
        RECT 363.000 10.000 365.500 25.000 ;
        RECT 335.500 7.500 365.500 10.000 ;
        RECT 397.000 4.500 400.000 30.500 ;
        RECT 301.500 1.500 400.000 4.500 ;
        RECT 451.500 30.500 550.000 33.500 ;
        RECT 451.500 4.500 457.500 30.500 ;
        RECT 485.500 25.000 515.500 27.500 ;
        RECT 485.500 10.000 488.000 25.000 ;
        RECT 513.000 10.000 515.500 25.000 ;
        RECT 485.500 7.500 515.500 10.000 ;
        RECT 544.000 4.500 550.000 30.500 ;
        RECT 451.500 1.500 550.000 4.500 ;
        RECT 601.500 30.500 700.000 33.500 ;
        RECT 601.500 4.500 607.500 30.500 ;
        RECT 635.500 25.000 665.500 27.500 ;
        RECT 635.500 10.000 638.000 25.000 ;
        RECT 663.000 10.000 665.500 25.000 ;
        RECT 635.500 7.500 665.500 10.000 ;
        RECT 694.000 4.500 700.000 30.500 ;
        RECT 601.500 1.500 700.000 4.500 ;
        RECT 751.500 30.500 850.000 33.500 ;
        RECT 751.500 4.500 760.500 30.500 ;
        RECT 785.500 25.000 815.500 27.500 ;
        RECT 785.500 10.000 788.000 25.000 ;
        RECT 813.000 10.000 815.500 25.000 ;
        RECT 785.500 7.500 815.500 10.000 ;
        RECT 841.000 4.500 850.000 30.500 ;
        RECT 751.500 1.500 850.000 4.500 ;
        RECT 901.500 30.500 1000.000 33.500 ;
        RECT 901.500 4.500 910.500 30.500 ;
        RECT 935.500 25.000 965.500 27.500 ;
        RECT 935.500 10.000 938.000 25.000 ;
        RECT 963.000 10.000 965.500 25.000 ;
        RECT 935.500 7.500 965.500 10.000 ;
        RECT 991.000 4.500 1000.000 30.500 ;
        RECT 901.500 1.500 1000.000 4.500 ;
        RECT 1051.500 30.500 1150.000 33.500 ;
        RECT 1051.500 4.500 1063.500 30.500 ;
        RECT 1085.500 25.000 1115.500 27.500 ;
        RECT 1085.500 10.000 1088.000 25.000 ;
        RECT 1113.000 10.000 1115.500 25.000 ;
        RECT 1085.500 7.500 1115.500 10.000 ;
        RECT 1138.000 4.500 1150.000 30.500 ;
        RECT 1051.500 1.500 1150.000 4.500 ;
        RECT 1201.500 30.500 1300.000 33.500 ;
        RECT 1201.500 4.500 1213.500 30.500 ;
        RECT 1235.500 25.000 1265.500 27.500 ;
        RECT 1235.500 10.000 1238.000 25.000 ;
        RECT 1263.000 10.000 1265.500 25.000 ;
        RECT 1235.500 7.500 1265.500 10.000 ;
        RECT 1288.000 4.500 1300.000 30.500 ;
        RECT 1201.500 1.500 1300.000 4.500 ;
        RECT 1351.500 30.500 1450.000 33.500 ;
        RECT 1351.500 4.500 1366.500 30.500 ;
        RECT 1385.500 25.000 1415.500 27.500 ;
        RECT 1385.500 10.000 1388.000 25.000 ;
        RECT 1413.000 10.000 1415.500 25.000 ;
        RECT 1385.500 7.500 1415.500 10.000 ;
        RECT 1435.000 4.500 1450.000 30.500 ;
        RECT 1351.500 1.500 1450.000 4.500 ;
        RECT 1501.500 30.500 1600.000 33.500 ;
        RECT 1501.500 4.500 1516.500 30.500 ;
        RECT 1535.500 25.000 1565.500 27.500 ;
        RECT 1535.500 10.000 1538.000 25.000 ;
        RECT 1563.000 10.000 1565.500 25.000 ;
        RECT 1535.500 7.500 1565.500 10.000 ;
        RECT 1585.000 4.500 1600.000 30.500 ;
        RECT 1501.500 1.500 1600.000 4.500 ;
        RECT 1651.500 30.500 1750.000 33.500 ;
        RECT 1651.500 4.500 1669.500 30.500 ;
        RECT 1685.500 25.000 1715.500 27.500 ;
        RECT 1685.500 10.000 1688.000 25.000 ;
        RECT 1713.000 10.000 1715.500 25.000 ;
        RECT 1685.500 7.500 1715.500 10.000 ;
        RECT 1732.000 4.500 1750.000 30.500 ;
        RECT 1651.500 1.500 1750.000 4.500 ;
        RECT 1801.500 30.500 1900.000 33.500 ;
        RECT 1801.500 4.500 1819.500 30.500 ;
        RECT 1835.500 25.000 1865.500 27.500 ;
        RECT 1835.500 10.000 1838.000 25.000 ;
        RECT 1863.000 10.000 1865.500 25.000 ;
        RECT 1835.500 7.500 1865.500 10.000 ;
        RECT 1882.000 4.500 1900.000 30.500 ;
        RECT 1801.500 1.500 1900.000 4.500 ;
      LAYER li1 ;
        RECT 152.500 2.500 153.500 32.500 ;
        RECT 196.500 31.500 203.500 32.500 ;
        RECT 186.500 14.500 187.500 21.500 ;
        RECT 213.500 14.500 214.500 21.500 ;
        RECT 196.500 2.500 203.500 3.500 ;
        RECT 248.000 2.500 249.000 32.500 ;
        RECT 302.500 2.500 303.500 32.500 ;
        RECT 346.500 31.500 353.500 32.500 ;
        RECT 336.500 14.500 337.500 21.500 ;
        RECT 363.500 14.500 364.500 21.500 ;
        RECT 346.500 2.500 353.500 3.500 ;
        RECT 398.000 2.500 399.000 32.500 ;
        RECT 452.500 2.500 453.500 32.500 ;
        RECT 496.500 31.500 503.500 32.500 ;
        RECT 486.500 14.500 487.500 21.500 ;
        RECT 513.500 14.500 514.500 21.500 ;
        RECT 496.500 2.500 503.500 3.500 ;
        RECT 548.000 2.500 549.000 32.500 ;
        RECT 602.500 2.500 603.500 32.500 ;
        RECT 646.500 31.500 653.500 32.500 ;
        RECT 636.500 14.500 637.500 21.500 ;
        RECT 663.500 14.500 664.500 21.500 ;
        RECT 646.500 2.500 653.500 3.500 ;
        RECT 698.000 2.500 699.000 32.500 ;
        RECT 752.500 2.500 753.500 32.500 ;
        RECT 796.500 31.500 803.500 32.500 ;
        RECT 786.500 14.500 787.500 21.500 ;
        RECT 813.500 14.500 814.500 21.500 ;
        RECT 796.500 2.500 803.500 3.500 ;
        RECT 848.000 2.500 849.000 32.500 ;
        RECT 902.500 2.500 903.500 32.500 ;
        RECT 946.500 31.500 953.500 32.500 ;
        RECT 936.500 14.500 937.500 21.500 ;
        RECT 963.500 14.500 964.500 21.500 ;
        RECT 946.500 2.500 953.500 3.500 ;
        RECT 998.000 2.500 999.000 32.500 ;
        RECT 1052.500 2.500 1053.500 32.500 ;
        RECT 1096.500 31.500 1103.500 32.500 ;
        RECT 1086.500 14.500 1087.500 21.500 ;
        RECT 1113.500 14.500 1114.500 21.500 ;
        RECT 1096.500 2.500 1103.500 3.500 ;
        RECT 1148.000 2.500 1149.000 32.500 ;
        RECT 1202.500 2.500 1203.500 32.500 ;
        RECT 1246.500 31.500 1253.500 32.500 ;
        RECT 1236.500 14.500 1237.500 21.500 ;
        RECT 1263.500 14.500 1264.500 21.500 ;
        RECT 1246.500 2.500 1253.500 3.500 ;
        RECT 1298.000 2.500 1299.000 32.500 ;
        RECT 1352.500 2.500 1353.500 32.500 ;
        RECT 1396.500 31.500 1403.500 32.500 ;
        RECT 1386.500 14.500 1387.500 21.500 ;
        RECT 1413.500 14.500 1414.500 21.500 ;
        RECT 1396.500 2.500 1403.500 3.500 ;
        RECT 1448.000 2.500 1449.000 32.500 ;
        RECT 1502.500 2.500 1503.500 32.500 ;
        RECT 1546.500 31.500 1553.500 32.500 ;
        RECT 1536.500 14.500 1537.500 21.500 ;
        RECT 1563.500 14.500 1564.500 21.500 ;
        RECT 1546.500 2.500 1553.500 3.500 ;
        RECT 1598.000 2.500 1599.000 32.500 ;
        RECT 1652.500 2.500 1653.500 32.500 ;
        RECT 1696.500 31.500 1703.500 32.500 ;
        RECT 1686.500 14.500 1687.500 21.500 ;
        RECT 1713.500 14.500 1714.500 21.500 ;
        RECT 1696.500 2.500 1703.500 3.500 ;
        RECT 1748.000 2.500 1749.000 32.500 ;
        RECT 1802.500 2.500 1803.500 32.500 ;
        RECT 1846.500 31.500 1853.500 32.500 ;
        RECT 1836.500 14.500 1837.500 21.500 ;
        RECT 1863.500 14.500 1864.500 21.500 ;
        RECT 1846.500 2.500 1853.500 3.500 ;
        RECT 1898.000 2.500 1899.000 32.500 ;
      LAYER met1 ;
        RECT 154.500 4.500 247.000 30.500 ;
        RECT 304.500 4.500 397.000 30.500 ;
        RECT 457.500 4.500 544.000 30.500 ;
        RECT 607.500 4.500 694.000 30.500 ;
        RECT 760.500 4.500 841.000 30.500 ;
        RECT 910.500 4.500 991.000 30.500 ;
        RECT 1063.500 4.500 1138.000 30.500 ;
        RECT 1213.500 4.500 1288.000 30.500 ;
        RECT 1363.500 4.500 1438.000 30.500 ;
        RECT 1513.500 4.500 1588.000 30.500 ;
        RECT 1663.500 4.500 1738.000 30.500 ;
        RECT 1813.500 4.500 1888.000 30.500 ;
      LAYER met2 ;
        RECT 150.000 0.000 251.500 35.500 ;
        RECT 300.000 0.000 402.000 36.000 ;
        RECT 450.000 0.000 552.000 36.000 ;
        RECT 600.000 0.000 702.000 36.000 ;
        RECT 750.000 0.000 852.000 36.000 ;
        RECT 900.000 0.000 1002.000 36.000 ;
        RECT 1050.000 0.000 1152.000 36.000 ;
        RECT 1200.000 0.000 1302.000 36.000 ;
        RECT 1350.000 0.000 1452.000 36.000 ;
        RECT 1500.000 0.000 1602.000 36.000 ;
        RECT 1650.000 0.000 1752.000 36.000 ;
        RECT 1800.000 0.000 1902.000 36.000 ;
      LAYER met3 ;
        RECT 150.000 0.000 251.500 35.500 ;
        RECT 300.000 0.000 402.000 36.000 ;
        RECT 450.000 0.000 552.000 36.000 ;
        RECT 600.000 0.000 702.000 36.000 ;
        RECT 750.000 0.000 852.000 36.000 ;
        RECT 900.000 0.000 1002.000 36.000 ;
        RECT 1050.000 0.000 1152.000 36.000 ;
        RECT 1200.000 0.000 1302.000 36.000 ;
        RECT 1350.000 0.000 1452.000 36.000 ;
        RECT 1500.000 0.000 1602.000 36.000 ;
        RECT 1650.000 0.000 1752.000 36.000 ;
        RECT 1800.000 0.000 1902.000 36.000 ;
      LAYER met4 ;
        RECT 150.000 0.000 251.500 35.500 ;
        RECT 300.000 0.000 402.000 36.000 ;
        RECT 450.000 0.000 552.000 36.000 ;
        RECT 600.000 0.000 702.000 36.000 ;
        RECT 750.000 0.000 852.000 36.000 ;
        RECT 900.000 0.000 1002.000 36.000 ;
        RECT 1050.000 0.000 1152.000 36.000 ;
        RECT 1200.000 0.000 1302.000 36.000 ;
        RECT 1350.000 0.000 1452.000 36.000 ;
        RECT 1500.000 0.000 1602.000 36.000 ;
        RECT 1650.000 0.000 1752.000 36.000 ;
        RECT 1800.000 0.000 1902.000 36.000 ;
      LAYER met5 ;
        RECT 150.000 0.000 251.500 35.500 ;
        RECT 300.000 0.000 402.000 36.000 ;
        RECT 450.000 0.000 552.000 36.000 ;
        RECT 600.000 0.000 702.000 36.000 ;
        RECT 750.000 0.000 852.000 36.000 ;
        RECT 900.000 0.000 1002.000 36.000 ;
        RECT 1050.000 0.000 1152.000 36.000 ;
        RECT 1200.000 0.000 1302.000 36.000 ;
        RECT 1350.000 0.000 1452.000 36.000 ;
        RECT 1500.000 0.000 1602.000 36.000 ;
        RECT 1650.000 0.000 1752.000 36.000 ;
        RECT 1800.000 0.000 1902.000 36.000 ;
  END
END PD1
END LIBRARY

