magic
tech sky130B
magscale 1 2
timestamp 1667857198
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 137830 700816 137836 700868
rect 137888 700856 137894 700868
rect 157978 700856 157984 700868
rect 137888 700828 157984 700856
rect 137888 700816 137894 700828
rect 157978 700816 157984 700828
rect 158036 700816 158042 700868
rect 155954 700748 155960 700800
rect 156012 700788 156018 700800
rect 202782 700788 202788 700800
rect 156012 700760 202788 700788
rect 156012 700748 156018 700760
rect 202782 700748 202788 700760
rect 202840 700748 202846 700800
rect 89162 700680 89168 700732
rect 89220 700720 89226 700732
rect 160738 700720 160744 700732
rect 89220 700692 160744 700720
rect 89220 700680 89226 700692
rect 160738 700680 160744 700692
rect 160796 700680 160802 700732
rect 154574 700612 154580 700664
rect 154632 700652 154638 700664
rect 267642 700652 267648 700664
rect 154632 700624 267648 700652
rect 154632 700612 154638 700624
rect 267642 700612 267648 700624
rect 267700 700612 267706 700664
rect 24302 700544 24308 700596
rect 24360 700584 24366 700596
rect 162210 700584 162216 700596
rect 24360 700556 162216 700584
rect 24360 700544 24366 700556
rect 162210 700544 162216 700556
rect 162268 700544 162274 700596
rect 8110 700476 8116 700528
rect 8168 700516 8174 700528
rect 162118 700516 162124 700528
rect 8168 700488 162124 700516
rect 8168 700476 8174 700488
rect 162118 700476 162124 700488
rect 162176 700476 162182 700528
rect 153838 700408 153844 700460
rect 153896 700448 153902 700460
rect 332502 700448 332508 700460
rect 153896 700420 332508 700448
rect 153896 700408 153902 700420
rect 332502 700408 332508 700420
rect 332560 700408 332566 700460
rect 152458 700340 152464 700392
rect 152516 700380 152522 700392
rect 413646 700380 413652 700392
rect 152516 700352 413652 700380
rect 152516 700340 152522 700352
rect 413646 700340 413652 700352
rect 413704 700340 413710 700392
rect 148318 700272 148324 700324
rect 148376 700312 148382 700324
rect 543458 700312 543464 700324
rect 148376 700284 543464 700312
rect 148376 700272 148382 700284
rect 543458 700272 543464 700284
rect 543516 700272 543522 700324
rect 559650 700312 559656 700324
rect 547846 700284 559656 700312
rect 542998 700204 543004 700256
rect 543056 700244 543062 700256
rect 547846 700244 547874 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 543056 700216 547874 700244
rect 543056 700204 543062 700216
rect 105446 699660 105452 699712
rect 105504 699700 105510 699712
rect 106918 699700 106924 699712
rect 105504 699672 106924 699700
rect 105504 699660 105510 699672
rect 106918 699660 106924 699672
rect 106976 699660 106982 699712
rect 396718 699660 396724 699712
rect 396776 699700 396782 699712
rect 397454 699700 397460 699712
rect 396776 699672 397460 699700
rect 396776 699660 396782 699672
rect 397454 699660 397460 699672
rect 397512 699660 397518 699712
rect 428458 699660 428464 699712
rect 428516 699700 428522 699712
rect 429838 699700 429844 699712
rect 428516 699672 429844 699700
rect 428516 699660 428522 699672
rect 429838 699660 429844 699672
rect 429896 699660 429902 699712
rect 146938 696940 146944 696992
rect 146996 696980 147002 696992
rect 580166 696980 580172 696992
rect 146996 696952 580172 696980
rect 146996 696940 147002 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 3418 683204 3424 683256
rect 3476 683244 3482 683256
rect 161474 683244 161480 683256
rect 3476 683216 161480 683244
rect 3476 683204 3482 683216
rect 161474 683204 161480 683216
rect 161532 683204 161538 683256
rect 147030 683136 147036 683188
rect 147088 683176 147094 683188
rect 580166 683176 580172 683188
rect 147088 683148 580172 683176
rect 147088 683136 147094 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 163498 670732 163504 670744
rect 3568 670704 163504 670732
rect 3568 670692 3574 670704
rect 163498 670692 163504 670704
rect 163556 670692 163562 670744
rect 185578 670692 185584 670744
rect 185636 670732 185642 670744
rect 580166 670732 580172 670744
rect 185636 670704 580172 670732
rect 185636 670692 185642 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 149054 660288 149060 660340
rect 149112 660328 149118 660340
rect 462314 660328 462320 660340
rect 149112 660300 462320 660328
rect 149112 660288 149118 660300
rect 462314 660288 462320 660300
rect 462372 660288 462378 660340
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 163590 656928 163596 656940
rect 3476 656900 163596 656928
rect 3476 656888 3482 656900
rect 163590 656888 163596 656900
rect 163648 656888 163654 656940
rect 184198 643084 184204 643136
rect 184256 643124 184262 643136
rect 580166 643124 580172 643136
rect 184256 643096 580172 643124
rect 184256 643084 184262 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 164234 632108 164240 632120
rect 3476 632080 164240 632108
rect 3476 632068 3482 632080
rect 164234 632068 164240 632080
rect 164292 632068 164298 632120
rect 203518 630640 203524 630692
rect 203576 630680 203582 630692
rect 580166 630680 580172 630692
rect 203576 630652 580172 630680
rect 203576 630640 203582 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 3142 618264 3148 618316
rect 3200 618304 3206 618316
rect 164878 618304 164884 618316
rect 3200 618276 164884 618304
rect 3200 618264 3206 618276
rect 164878 618264 164884 618276
rect 164936 618264 164942 618316
rect 143534 616836 143540 616888
rect 143592 616876 143598 616888
rect 580166 616876 580172 616888
rect 143592 616848 580172 616876
rect 143592 616836 143598 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3234 605820 3240 605872
rect 3292 605860 3298 605872
rect 164970 605860 164976 605872
rect 3292 605832 164976 605860
rect 3292 605820 3298 605832
rect 164970 605820 164976 605832
rect 165028 605820 165034 605872
rect 142154 590656 142160 590708
rect 142212 590696 142218 590708
rect 579798 590696 579804 590708
rect 142212 590668 579804 590696
rect 142212 590656 142218 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 165614 579680 165620 579692
rect 3384 579652 165620 579680
rect 3384 579640 3390 579652
rect 165614 579640 165620 579652
rect 165672 579640 165678 579692
rect 144178 576852 144184 576904
rect 144236 576892 144242 576904
rect 580166 576892 580172 576904
rect 144236 576864 580172 576892
rect 144236 576852 144242 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 3418 565836 3424 565888
rect 3476 565876 3482 565888
rect 167638 565876 167644 565888
rect 3476 565848 167644 565876
rect 3476 565836 3482 565848
rect 167638 565836 167644 565848
rect 167696 565836 167702 565888
rect 142798 563048 142804 563100
rect 142856 563088 142862 563100
rect 579798 563088 579804 563100
rect 142856 563060 579804 563088
rect 142856 563048 142862 563060
rect 579798 563048 579804 563060
rect 579856 563048 579862 563100
rect 3418 553392 3424 553444
rect 3476 553432 3482 553444
rect 166258 553432 166264 553444
rect 3476 553404 166264 553432
rect 3476 553392 3482 553404
rect 166258 553392 166264 553404
rect 166316 553392 166322 553444
rect 178678 536800 178684 536852
rect 178736 536840 178742 536852
rect 580166 536840 580172 536852
rect 178736 536812 580172 536840
rect 178736 536800 178742 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 3418 527144 3424 527196
rect 3476 527184 3482 527196
rect 166994 527184 167000 527196
rect 3476 527156 167000 527184
rect 3476 527144 3482 527156
rect 166994 527144 167000 527156
rect 167052 527144 167058 527196
rect 142890 524424 142896 524476
rect 142948 524464 142954 524476
rect 580166 524464 580172 524476
rect 142948 524436 580172 524464
rect 142948 524424 142954 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3418 514768 3424 514820
rect 3476 514808 3482 514820
rect 8938 514808 8944 514820
rect 3476 514780 8944 514808
rect 3476 514768 3482 514780
rect 8938 514768 8944 514780
rect 8996 514768 9002 514820
rect 181438 510620 181444 510672
rect 181496 510660 181502 510672
rect 580166 510660 580172 510672
rect 181496 510632 580172 510660
rect 181496 510620 181502 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 3050 500964 3056 501016
rect 3108 501004 3114 501016
rect 167270 501004 167276 501016
rect 3108 500976 167276 501004
rect 3108 500964 3114 500976
rect 167270 500964 167276 500976
rect 167328 500964 167334 501016
rect 139394 484372 139400 484424
rect 139452 484412 139458 484424
rect 580166 484412 580172 484424
rect 139452 484384 580172 484412
rect 139452 484372 139458 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 139670 470568 139676 470620
rect 139728 470608 139734 470620
rect 579982 470608 579988 470620
rect 139728 470580 579988 470608
rect 139728 470568 139734 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 3510 462340 3516 462392
rect 3568 462380 3574 462392
rect 170398 462380 170404 462392
rect 3568 462352 170404 462380
rect 3568 462340 3574 462352
rect 170398 462340 170404 462352
rect 170456 462340 170462 462392
rect 180058 456764 180064 456816
rect 180116 456804 180122 456816
rect 580166 456804 580172 456816
rect 180116 456776 580172 456804
rect 180116 456764 180122 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 170490 448576 170496 448588
rect 3200 448548 170496 448576
rect 3200 448536 3206 448548
rect 170490 448536 170496 448548
rect 170548 448536 170554 448588
rect 158622 447788 158628 447840
rect 158680 447828 158686 447840
rect 169754 447828 169760 447840
rect 158680 447800 169760 447828
rect 158680 447788 158686 447800
rect 169754 447788 169760 447800
rect 169812 447788 169818 447840
rect 138658 430584 138664 430636
rect 138716 430624 138722 430636
rect 580166 430624 580172 430636
rect 138716 430596 580172 430624
rect 138716 430584 138722 430596
rect 580166 430584 580172 430596
rect 580224 430584 580230 430636
rect 3510 422288 3516 422340
rect 3568 422328 3574 422340
rect 169754 422328 169760 422340
rect 3568 422300 169760 422328
rect 3568 422288 3574 422300
rect 169754 422288 169760 422300
rect 169812 422288 169818 422340
rect 138750 418140 138756 418192
rect 138808 418180 138814 418192
rect 580166 418180 580172 418192
rect 138808 418152 580172 418180
rect 138808 418140 138814 418152
rect 580166 418140 580172 418152
rect 580224 418140 580230 418192
rect 2866 409844 2872 409896
rect 2924 409884 2930 409896
rect 171778 409884 171784 409896
rect 2924 409856 171784 409884
rect 2924 409844 2930 409856
rect 171778 409844 171784 409856
rect 171836 409844 171842 409896
rect 199378 404336 199384 404388
rect 199436 404376 199442 404388
rect 580166 404376 580172 404388
rect 199436 404348 580172 404376
rect 199436 404336 199442 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 3510 397468 3516 397520
rect 3568 397508 3574 397520
rect 171870 397508 171876 397520
rect 3568 397480 171876 397508
rect 3568 397468 3574 397480
rect 171870 397468 171876 397480
rect 171928 397468 171934 397520
rect 182818 378156 182824 378208
rect 182876 378196 182882 378208
rect 580166 378196 580172 378208
rect 182876 378168 580172 378196
rect 182876 378156 182882 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 2774 371288 2780 371340
rect 2832 371328 2838 371340
rect 4798 371328 4804 371340
rect 2832 371300 4804 371328
rect 2832 371288 2838 371300
rect 4798 371288 4804 371300
rect 4856 371288 4862 371340
rect 3142 357416 3148 357468
rect 3200 357456 3206 357468
rect 10318 357456 10324 357468
rect 3200 357428 10324 357456
rect 3200 357416 3206 357428
rect 10318 357416 10324 357428
rect 10376 357416 10382 357468
rect 135254 351908 135260 351960
rect 135312 351948 135318 351960
rect 580166 351948 580172 351960
rect 135312 351920 580172 351948
rect 135312 351908 135318 351920
rect 580166 351908 580172 351920
rect 580224 351908 580230 351960
rect 3510 345176 3516 345228
rect 3568 345216 3574 345228
rect 7558 345216 7564 345228
rect 3568 345188 7564 345216
rect 3568 345176 3574 345188
rect 7558 345176 7564 345188
rect 7616 345176 7622 345228
rect 134518 324300 134524 324352
rect 134576 324340 134582 324352
rect 580166 324340 580172 324352
rect 134576 324312 580172 324340
rect 134576 324300 134582 324312
rect 580166 324300 580172 324312
rect 580224 324300 580230 324352
rect 3326 318792 3332 318844
rect 3384 318832 3390 318844
rect 173894 318832 173900 318844
rect 3384 318804 173900 318832
rect 3384 318792 3390 318804
rect 173894 318792 173900 318804
rect 173952 318792 173958 318844
rect 135898 311856 135904 311908
rect 135956 311896 135962 311908
rect 579982 311896 579988 311908
rect 135956 311868 579988 311896
rect 135956 311856 135962 311868
rect 579982 311856 579988 311868
rect 580040 311856 580046 311908
rect 3510 304988 3516 305040
rect 3568 305028 3574 305040
rect 175918 305028 175924 305040
rect 3568 305000 175924 305028
rect 3568 304988 3574 305000
rect 175918 304988 175924 305000
rect 175976 304988 175982 305040
rect 134610 298120 134616 298172
rect 134668 298160 134674 298172
rect 580166 298160 580172 298172
rect 134668 298132 580172 298160
rect 134668 298120 134674 298132
rect 580166 298120 580172 298132
rect 580224 298120 580230 298172
rect 3510 292544 3516 292596
rect 3568 292584 3574 292596
rect 174538 292584 174544 292596
rect 3568 292556 174544 292584
rect 3568 292544 3574 292556
rect 174538 292544 174544 292556
rect 174596 292544 174602 292596
rect 10318 289076 10324 289128
rect 10376 289116 10382 289128
rect 173158 289116 173164 289128
rect 10376 289088 173164 289116
rect 10376 289076 10382 289088
rect 173158 289076 173164 289088
rect 173216 289076 173222 289128
rect 145558 287648 145564 287700
rect 145616 287688 145622 287700
rect 203518 287688 203524 287700
rect 145616 287660 203524 287688
rect 145616 287648 145622 287660
rect 203518 287648 203524 287660
rect 203576 287648 203582 287700
rect 137278 286288 137284 286340
rect 137336 286328 137342 286340
rect 182818 286328 182824 286340
rect 137336 286300 182824 286328
rect 137336 286288 137342 286300
rect 182818 286288 182824 286300
rect 182876 286288 182882 286340
rect 150434 284928 150440 284980
rect 150492 284968 150498 284980
rect 396718 284968 396724 284980
rect 150492 284940 396724 284968
rect 150492 284928 150498 284940
rect 396718 284928 396724 284940
rect 396776 284928 396782 284980
rect 147674 283568 147680 283620
rect 147732 283608 147738 283620
rect 527174 283608 527180 283620
rect 147732 283580 527180 283608
rect 147732 283568 147738 283580
rect 527174 283568 527180 283580
rect 527232 283568 527238 283620
rect 145650 282140 145656 282192
rect 145708 282180 145714 282192
rect 184198 282180 184204 282192
rect 145708 282152 184204 282180
rect 145708 282140 145714 282152
rect 184198 282140 184204 282152
rect 184256 282140 184262 282192
rect 140774 280780 140780 280832
rect 140832 280820 140838 280832
rect 178678 280820 178684 280832
rect 140832 280792 178684 280820
rect 140832 280780 140838 280792
rect 178678 280780 178684 280792
rect 178736 280780 178742 280832
rect 40034 279420 40040 279472
rect 40092 279460 40098 279472
rect 160094 279460 160100 279472
rect 40092 279432 160100 279460
rect 40092 279420 40098 279432
rect 160094 279420 160100 279432
rect 160152 279420 160158 279472
rect 189074 277992 189080 278044
rect 189132 278032 189138 278044
rect 234614 278032 234620 278044
rect 189132 278004 234620 278032
rect 189132 277992 189138 278004
rect 234614 277992 234620 278004
rect 234672 277992 234678 278044
rect 156046 277380 156052 277432
rect 156104 277420 156110 277432
rect 189074 277420 189080 277432
rect 156104 277392 189080 277420
rect 156104 277380 156110 277392
rect 189074 277380 189080 277392
rect 189132 277380 189138 277432
rect 204714 276632 204720 276684
rect 204772 276672 204778 276684
rect 299474 276672 299480 276684
rect 204772 276644 299480 276672
rect 204772 276632 204778 276644
rect 299474 276632 299480 276644
rect 299532 276632 299538 276684
rect 153286 276020 153292 276072
rect 153344 276060 153350 276072
rect 204438 276060 204444 276072
rect 153344 276032 204444 276060
rect 153344 276020 153350 276032
rect 204438 276020 204444 276032
rect 204496 276060 204502 276072
rect 204714 276060 204720 276072
rect 204496 276032 204720 276060
rect 204496 276020 204502 276032
rect 204714 276020 204720 276032
rect 204772 276020 204778 276072
rect 8938 273980 8944 274032
rect 8996 274020 9002 274032
rect 169018 274020 169024 274032
rect 8996 273992 169024 274020
rect 8996 273980 9002 273992
rect 169018 273980 169024 273992
rect 169076 273980 169082 274032
rect 151078 273912 151084 273964
rect 151136 273952 151142 273964
rect 428458 273952 428464 273964
rect 151136 273924 428464 273952
rect 151136 273912 151142 273924
rect 428458 273912 428464 273924
rect 428516 273912 428522 273964
rect 133138 271872 133144 271924
rect 133196 271912 133202 271924
rect 580166 271912 580172 271924
rect 133196 271884 580172 271912
rect 133196 271872 133202 271884
rect 580166 271872 580172 271884
rect 580224 271872 580230 271924
rect 7558 271192 7564 271244
rect 7616 271232 7622 271244
rect 172514 271232 172520 271244
rect 7616 271204 172520 271232
rect 7616 271192 7622 271204
rect 172514 271192 172520 271204
rect 172572 271192 172578 271244
rect 149146 271124 149152 271176
rect 149204 271164 149210 271176
rect 494054 271164 494060 271176
rect 149204 271136 494060 271164
rect 149204 271124 149210 271136
rect 494054 271124 494060 271136
rect 494112 271124 494118 271176
rect 71774 269832 71780 269884
rect 71832 269872 71838 269884
rect 158806 269872 158812 269884
rect 71832 269844 158812 269872
rect 71832 269832 71838 269844
rect 158806 269832 158812 269844
rect 158864 269832 158870 269884
rect 147766 269764 147772 269816
rect 147824 269804 147830 269816
rect 542998 269804 543004 269816
rect 147824 269776 543004 269804
rect 147824 269764 147830 269776
rect 542998 269764 543004 269776
rect 543056 269764 543062 269816
rect 146202 268404 146208 268456
rect 146260 268444 146266 268456
rect 185578 268444 185584 268456
rect 146260 268416 185584 268444
rect 146260 268404 146266 268416
rect 185578 268404 185584 268416
rect 185636 268404 185642 268456
rect 4798 268336 4804 268388
rect 4856 268376 4862 268388
rect 172698 268376 172704 268388
rect 4856 268348 172704 268376
rect 4856 268336 4862 268348
rect 172698 268336 172704 268348
rect 172756 268336 172762 268388
rect 137830 266976 137836 267028
rect 137888 267016 137894 267028
rect 199378 267016 199384 267028
rect 137888 266988 199384 267016
rect 137888 266976 137894 266988
rect 199378 266976 199384 266988
rect 199436 266976 199442 267028
rect 3050 266364 3056 266416
rect 3108 266404 3114 266416
rect 175918 266404 175924 266416
rect 3108 266376 175924 266404
rect 3108 266364 3114 266376
rect 175918 266364 175924 266376
rect 175976 266364 175982 266416
rect 164878 265820 164884 265872
rect 164936 265860 164942 265872
rect 165154 265860 165160 265872
rect 164936 265832 165160 265860
rect 164936 265820 164942 265832
rect 165154 265820 165160 265832
rect 165212 265820 165218 265872
rect 141418 265684 141424 265736
rect 141476 265724 141482 265736
rect 181438 265724 181444 265736
rect 141476 265696 181444 265724
rect 141476 265684 141482 265696
rect 181438 265684 181444 265696
rect 181496 265684 181502 265736
rect 3418 265616 3424 265668
rect 3476 265656 3482 265668
rect 169110 265656 169116 265668
rect 3476 265628 169116 265656
rect 3476 265616 3482 265628
rect 169110 265616 169116 265628
rect 169168 265616 169174 265668
rect 174538 265548 174544 265600
rect 174596 265588 174602 265600
rect 174596 265560 180794 265588
rect 174596 265548 174602 265560
rect 180766 265520 180794 265560
rect 195974 265520 195980 265532
rect 180766 265492 195980 265520
rect 195974 265480 195980 265492
rect 196032 265480 196038 265532
rect 166258 265412 166264 265464
rect 166316 265452 166322 265464
rect 192110 265452 192116 265464
rect 166316 265424 192116 265452
rect 166316 265412 166322 265424
rect 192110 265412 192116 265424
rect 192168 265412 192174 265464
rect 171778 265344 171784 265396
rect 171836 265384 171842 265396
rect 197630 265384 197636 265396
rect 171836 265356 197636 265384
rect 171836 265344 171842 265356
rect 197630 265344 197636 265356
rect 197688 265344 197694 265396
rect 173434 265276 173440 265328
rect 173492 265316 173498 265328
rect 199194 265316 199200 265328
rect 173492 265288 199200 265316
rect 173492 265276 173498 265288
rect 199194 265276 199200 265288
rect 199252 265276 199258 265328
rect 170398 265208 170404 265260
rect 170456 265248 170462 265260
rect 170674 265248 170680 265260
rect 170456 265220 170680 265248
rect 170456 265208 170462 265220
rect 170674 265208 170680 265220
rect 170732 265248 170738 265260
rect 199102 265248 199108 265260
rect 170732 265220 199108 265248
rect 170732 265208 170738 265220
rect 199102 265208 199108 265220
rect 199160 265208 199166 265260
rect 113082 265140 113088 265192
rect 113140 265180 113146 265192
rect 138750 265180 138756 265192
rect 113140 265152 138756 265180
rect 113140 265140 113146 265152
rect 138750 265140 138756 265152
rect 138808 265140 138814 265192
rect 162210 265140 162216 265192
rect 162268 265180 162274 265192
rect 195238 265180 195244 265192
rect 162268 265152 195244 265180
rect 162268 265140 162274 265152
rect 195238 265140 195244 265152
rect 195296 265140 195302 265192
rect 116578 265072 116584 265124
rect 116636 265112 116642 265124
rect 143626 265112 143632 265124
rect 116636 265084 143632 265112
rect 116636 265072 116642 265084
rect 143626 265072 143632 265084
rect 143684 265112 143690 265124
rect 144178 265112 144184 265124
rect 143684 265084 144184 265112
rect 143684 265072 143690 265084
rect 144178 265072 144184 265084
rect 144236 265072 144242 265124
rect 170214 265072 170220 265124
rect 170272 265112 170278 265124
rect 170490 265112 170496 265124
rect 170272 265084 170496 265112
rect 170272 265072 170278 265084
rect 170490 265072 170496 265084
rect 170548 265112 170554 265124
rect 203242 265112 203248 265124
rect 170548 265084 203248 265112
rect 170548 265072 170554 265084
rect 203242 265072 203248 265084
rect 203300 265072 203306 265124
rect 112806 265004 112812 265056
rect 112864 265044 112870 265056
rect 145558 265044 145564 265056
rect 112864 265016 145564 265044
rect 112864 265004 112870 265016
rect 145558 265004 145564 265016
rect 145616 265004 145622 265056
rect 160830 265004 160836 265056
rect 160888 265044 160894 265056
rect 194870 265044 194876 265056
rect 160888 265016 194876 265044
rect 160888 265004 160894 265016
rect 194870 265004 194876 265016
rect 194928 265004 194934 265056
rect 119614 264936 119620 264988
rect 119672 264976 119678 264988
rect 152182 264976 152188 264988
rect 119672 264948 152188 264976
rect 119672 264936 119678 264948
rect 152182 264936 152188 264948
rect 152240 264976 152246 264988
rect 152458 264976 152464 264988
rect 152240 264948 152464 264976
rect 152240 264936 152246 264948
rect 152458 264936 152464 264948
rect 152516 264936 152522 264988
rect 165154 264936 165160 264988
rect 165212 264976 165218 264988
rect 203150 264976 203156 264988
rect 165212 264948 203156 264976
rect 165212 264936 165218 264948
rect 203150 264936 203156 264948
rect 203208 264936 203214 264988
rect 106918 264188 106924 264240
rect 106976 264228 106982 264240
rect 118694 264228 118700 264240
rect 106976 264200 118700 264228
rect 106976 264188 106982 264200
rect 118694 264188 118700 264200
rect 118752 264188 118758 264240
rect 139394 264188 139400 264240
rect 139452 264228 139458 264240
rect 180058 264228 180064 264240
rect 139452 264200 180064 264228
rect 139452 264188 139458 264200
rect 180058 264188 180064 264200
rect 180116 264188 180122 264240
rect 120994 263916 121000 263968
rect 121052 263956 121058 263968
rect 134242 263956 134248 263968
rect 121052 263928 134248 263956
rect 121052 263916 121058 263928
rect 134242 263916 134248 263928
rect 134300 263956 134306 263968
rect 134610 263956 134616 263968
rect 134300 263928 134616 263956
rect 134300 263916 134306 263928
rect 134610 263916 134616 263928
rect 134668 263916 134674 263968
rect 119522 263848 119528 263900
rect 119580 263888 119586 263900
rect 137830 263888 137836 263900
rect 119580 263860 137836 263888
rect 119580 263848 119586 263860
rect 137830 263848 137836 263860
rect 137888 263848 137894 263900
rect 120902 263780 120908 263832
rect 120960 263820 120966 263832
rect 139394 263820 139400 263832
rect 120960 263792 139400 263820
rect 120960 263780 120966 263792
rect 139394 263780 139400 263792
rect 139452 263780 139458 263832
rect 117958 263712 117964 263764
rect 118016 263752 118022 263764
rect 137186 263752 137192 263764
rect 118016 263724 137192 263752
rect 118016 263712 118022 263724
rect 137186 263712 137192 263724
rect 137244 263712 137250 263764
rect 172698 263712 172704 263764
rect 172756 263752 172762 263764
rect 190638 263752 190644 263764
rect 172756 263724 190644 263752
rect 172756 263712 172762 263724
rect 190638 263712 190644 263724
rect 190696 263712 190702 263764
rect 119706 263644 119712 263696
rect 119764 263684 119770 263696
rect 141142 263684 141148 263696
rect 119764 263656 141148 263684
rect 119764 263644 119770 263656
rect 141142 263644 141148 263656
rect 141200 263684 141206 263696
rect 141418 263684 141424 263696
rect 141200 263656 141424 263684
rect 141200 263644 141206 263656
rect 141418 263644 141424 263656
rect 141476 263644 141482 263696
rect 157886 263644 157892 263696
rect 157944 263684 157950 263696
rect 158622 263684 158628 263696
rect 157944 263656 158628 263684
rect 157944 263644 157950 263656
rect 158622 263644 158628 263656
rect 158680 263684 158686 263696
rect 188246 263684 188252 263696
rect 158680 263656 188252 263684
rect 158680 263644 158686 263656
rect 188246 263644 188252 263656
rect 188304 263644 188310 263696
rect 118694 263576 118700 263628
rect 118752 263616 118758 263628
rect 119982 263616 119988 263628
rect 118752 263588 119988 263616
rect 118752 263576 118758 263588
rect 119982 263576 119988 263588
rect 120040 263616 120046 263628
rect 159082 263616 159088 263628
rect 120040 263588 159088 263616
rect 120040 263576 120046 263588
rect 159082 263576 159088 263588
rect 159140 263576 159146 263628
rect 175734 263576 175740 263628
rect 175792 263616 175798 263628
rect 197722 263616 197728 263628
rect 175792 263588 197728 263616
rect 175792 263576 175798 263588
rect 197722 263576 197728 263588
rect 197780 263576 197786 263628
rect 137462 263508 137468 263560
rect 137520 263548 137526 263560
rect 580258 263548 580264 263560
rect 137520 263520 580264 263548
rect 137520 263508 137526 263520
rect 580258 263508 580264 263520
rect 580316 263508 580322 263560
rect 189994 263440 190000 263492
rect 190052 263480 190058 263492
rect 282914 263480 282920 263492
rect 190052 263452 282920 263480
rect 190052 263440 190058 263452
rect 282914 263440 282920 263452
rect 282972 263440 282978 263492
rect 171686 263372 171692 263424
rect 171744 263412 171750 263424
rect 171870 263412 171876 263424
rect 171744 263384 171876 263412
rect 171744 263372 171750 263384
rect 171870 263372 171876 263384
rect 171928 263372 171934 263424
rect 163406 263236 163412 263288
rect 163464 263276 163470 263288
rect 163590 263276 163596 263288
rect 163464 263248 163596 263276
rect 163464 263236 163470 263248
rect 163590 263236 163596 263248
rect 163648 263236 163654 263288
rect 116854 263100 116860 263152
rect 116912 263140 116918 263152
rect 129274 263140 129280 263152
rect 116912 263112 129280 263140
rect 116912 263100 116918 263112
rect 129274 263100 129280 263112
rect 129332 263100 129338 263152
rect 171686 263100 171692 263152
rect 171744 263140 171750 263152
rect 196618 263140 196624 263152
rect 171744 263112 196624 263140
rect 171744 263100 171750 263112
rect 196618 263100 196624 263112
rect 196676 263100 196682 263152
rect 3418 263032 3424 263084
rect 3476 263072 3482 263084
rect 178402 263072 178408 263084
rect 3476 263044 178408 263072
rect 3476 263032 3482 263044
rect 178402 263032 178408 263044
rect 178460 263032 178466 263084
rect 180150 263032 180156 263084
rect 180208 263072 180214 263084
rect 194962 263072 194968 263084
rect 180208 263044 194968 263072
rect 180208 263032 180214 263044
rect 194962 263032 194968 263044
rect 195020 263032 195026 263084
rect 117038 262964 117044 263016
rect 117096 263004 117102 263016
rect 125962 263004 125968 263016
rect 117096 262976 125968 263004
rect 117096 262964 117102 262976
rect 125962 262964 125968 262976
rect 126020 262964 126026 263016
rect 132310 262964 132316 263016
rect 132368 263004 132374 263016
rect 580350 263004 580356 263016
rect 132368 262976 580356 263004
rect 132368 262964 132374 262976
rect 580350 262964 580356 262976
rect 580408 262964 580414 263016
rect 116670 262896 116676 262948
rect 116728 262936 116734 262948
rect 127526 262936 127532 262948
rect 116728 262908 127532 262936
rect 116728 262896 116734 262908
rect 127526 262896 127532 262908
rect 127584 262896 127590 262948
rect 580442 262936 580448 262948
rect 132466 262908 580448 262936
rect 115382 262828 115388 262880
rect 115440 262868 115446 262880
rect 131758 262868 131764 262880
rect 115440 262840 131764 262868
rect 115440 262828 115446 262840
rect 131758 262828 131764 262840
rect 131816 262868 131822 262880
rect 132466 262868 132494 262908
rect 580442 262896 580448 262908
rect 580500 262896 580506 262948
rect 218054 262868 218060 262880
rect 131816 262840 132494 262868
rect 200086 262840 218060 262868
rect 131816 262828 131822 262840
rect 115474 262760 115480 262812
rect 115532 262800 115538 262812
rect 134518 262800 134524 262812
rect 115532 262772 134524 262800
rect 115532 262760 115538 262772
rect 134518 262760 134524 262772
rect 134576 262800 134582 262812
rect 134794 262800 134800 262812
rect 134576 262772 134800 262800
rect 134576 262760 134582 262772
rect 134794 262760 134800 262772
rect 134852 262760 134858 262812
rect 153194 262760 153200 262812
rect 153252 262800 153258 262812
rect 158714 262800 158720 262812
rect 153252 262772 158720 262800
rect 153252 262760 153258 262772
rect 158714 262760 158720 262772
rect 158772 262760 158778 262812
rect 164970 262760 164976 262812
rect 165028 262800 165034 262812
rect 193582 262800 193588 262812
rect 165028 262772 193588 262800
rect 165028 262760 165034 262772
rect 193582 262760 193588 262772
rect 193640 262760 193646 262812
rect 118326 262692 118332 262744
rect 118384 262732 118390 262744
rect 122834 262732 122840 262744
rect 118384 262704 122840 262732
rect 118384 262692 118390 262704
rect 122834 262692 122840 262704
rect 122892 262692 122898 262744
rect 127526 262692 127532 262744
rect 127584 262732 127590 262744
rect 133138 262732 133144 262744
rect 127584 262704 133144 262732
rect 127584 262692 127590 262704
rect 133138 262692 133144 262704
rect 133196 262692 133202 262744
rect 163406 262692 163412 262744
rect 163464 262732 163470 262744
rect 192478 262732 192484 262744
rect 163464 262704 192484 262732
rect 163464 262692 163470 262704
rect 192478 262692 192484 262704
rect 192536 262692 192542 262744
rect 118234 262624 118240 262676
rect 118292 262664 118298 262676
rect 127618 262664 127624 262676
rect 118292 262636 127624 262664
rect 118292 262624 118298 262636
rect 127618 262624 127624 262636
rect 127676 262624 127682 262676
rect 157978 262624 157984 262676
rect 158036 262664 158042 262676
rect 192202 262664 192208 262676
rect 158036 262636 192208 262664
rect 158036 262624 158042 262636
rect 192202 262624 192208 262636
rect 192260 262624 192266 262676
rect 114002 262556 114008 262608
rect 114060 262596 114066 262608
rect 129826 262596 129832 262608
rect 114060 262568 129832 262596
rect 114060 262556 114066 262568
rect 129826 262556 129832 262568
rect 129884 262556 129890 262608
rect 155862 262556 155868 262608
rect 155920 262596 155926 262608
rect 189258 262596 189264 262608
rect 155920 262568 189264 262596
rect 155920 262556 155926 262568
rect 189258 262556 189264 262568
rect 189316 262596 189322 262608
rect 189994 262596 190000 262608
rect 189316 262568 190000 262596
rect 189316 262556 189322 262568
rect 189994 262556 190000 262568
rect 190052 262556 190058 262608
rect 119798 262488 119804 262540
rect 119856 262528 119862 262540
rect 153286 262528 153292 262540
rect 119856 262500 153292 262528
rect 119856 262488 119862 262500
rect 153286 262488 153292 262500
rect 153344 262528 153350 262540
rect 153838 262528 153844 262540
rect 153344 262500 153844 262528
rect 153344 262488 153350 262500
rect 153838 262488 153844 262500
rect 153896 262488 153902 262540
rect 157150 262488 157156 262540
rect 157208 262528 157214 262540
rect 192386 262528 192392 262540
rect 157208 262500 192392 262528
rect 157208 262488 157214 262500
rect 192386 262488 192392 262500
rect 192444 262528 192450 262540
rect 200086 262528 200114 262840
rect 218054 262828 218060 262840
rect 218112 262828 218118 262880
rect 192444 262500 200114 262528
rect 192444 262488 192450 262500
rect 3510 262420 3516 262472
rect 3568 262460 3574 262472
rect 176746 262460 176752 262472
rect 3568 262432 176752 262460
rect 3568 262420 3574 262432
rect 176746 262420 176752 262432
rect 176804 262420 176810 262472
rect 179230 262420 179236 262472
rect 179288 262460 179294 262472
rect 192662 262460 192668 262472
rect 179288 262432 192668 262460
rect 179288 262420 179294 262432
rect 192662 262420 192668 262432
rect 192720 262420 192726 262472
rect 122834 262352 122840 262404
rect 122892 262392 122898 262404
rect 131114 262392 131120 262404
rect 122892 262364 131120 262392
rect 122892 262352 122898 262364
rect 131114 262352 131120 262364
rect 131172 262352 131178 262404
rect 182910 262352 182916 262404
rect 182968 262392 182974 262404
rect 190454 262392 190460 262404
rect 182968 262364 190460 262392
rect 182968 262352 182974 262364
rect 190454 262352 190460 262364
rect 190512 262352 190518 262404
rect 181254 262284 181260 262336
rect 181312 262324 181318 262336
rect 190546 262324 190552 262336
rect 181312 262296 190552 262324
rect 181312 262284 181318 262296
rect 190546 262284 190552 262296
rect 190604 262284 190610 262336
rect 116486 262216 116492 262268
rect 116544 262256 116550 262268
rect 122742 262256 122748 262268
rect 116544 262228 122748 262256
rect 116544 262216 116550 262228
rect 122742 262216 122748 262228
rect 122800 262216 122806 262268
rect 184566 262216 184572 262268
rect 184624 262256 184630 262268
rect 189166 262256 189172 262268
rect 184624 262228 189172 262256
rect 184624 262216 184630 262228
rect 189166 262216 189172 262228
rect 189224 262216 189230 262268
rect 158714 261604 158720 261656
rect 158772 261644 158778 261656
rect 193674 261644 193680 261656
rect 158772 261616 193680 261644
rect 158772 261604 158778 261616
rect 193674 261604 193680 261616
rect 193732 261604 193738 261656
rect 129826 261536 129832 261588
rect 129884 261576 129890 261588
rect 189810 261576 189816 261588
rect 129884 261548 189816 261576
rect 129884 261536 129890 261548
rect 189810 261536 189816 261548
rect 189868 261536 189874 261588
rect 176746 261468 176752 261520
rect 176804 261508 176810 261520
rect 199286 261508 199292 261520
rect 176804 261480 199292 261508
rect 176804 261468 176810 261480
rect 199286 261468 199292 261480
rect 199344 261468 199350 261520
rect 131114 261400 131120 261452
rect 131172 261440 131178 261452
rect 471238 261440 471244 261452
rect 131172 261412 471244 261440
rect 131172 261400 131178 261412
rect 471238 261400 471244 261412
rect 471296 261400 471302 261452
rect 181806 261332 181812 261384
rect 181864 261372 181870 261384
rect 193490 261372 193496 261384
rect 181864 261344 193496 261372
rect 181864 261332 181870 261344
rect 193490 261332 193496 261344
rect 193548 261332 193554 261384
rect 177298 261264 177304 261316
rect 177356 261304 177362 261316
rect 193766 261304 193772 261316
rect 177356 261276 193772 261304
rect 177356 261264 177362 261276
rect 193766 261264 193772 261276
rect 193824 261264 193830 261316
rect 178402 261196 178408 261248
rect 178460 261236 178466 261248
rect 197906 261236 197912 261248
rect 178460 261208 197912 261236
rect 178460 261196 178466 261208
rect 197906 261196 197912 261208
rect 197964 261196 197970 261248
rect 112898 261128 112904 261180
rect 112956 261168 112962 261180
rect 128722 261168 128728 261180
rect 112956 261140 128728 261168
rect 112956 261128 112962 261140
rect 128722 261128 128728 261140
rect 128780 261128 128786 261180
rect 176194 261128 176200 261180
rect 176252 261168 176258 261180
rect 195054 261168 195060 261180
rect 176252 261140 195060 261168
rect 176252 261128 176258 261140
rect 195054 261128 195060 261140
rect 195112 261128 195118 261180
rect 116762 261060 116768 261112
rect 116820 261100 116826 261112
rect 133230 261100 133236 261112
rect 116820 261072 133236 261100
rect 116820 261060 116826 261072
rect 133230 261060 133236 261072
rect 133288 261060 133294 261112
rect 184014 261060 184020 261112
rect 184072 261100 184078 261112
rect 196434 261100 196440 261112
rect 184072 261072 196440 261100
rect 184072 261060 184078 261072
rect 196434 261060 196440 261072
rect 196492 261060 196498 261112
rect 111058 260992 111064 261044
rect 111116 261032 111122 261044
rect 127066 261032 127072 261044
rect 111116 261004 127072 261032
rect 111116 260992 111122 261004
rect 127066 260992 127072 261004
rect 127124 260992 127130 261044
rect 180518 260992 180524 261044
rect 180576 261032 180582 261044
rect 197998 261032 198004 261044
rect 180576 261004 198004 261032
rect 180576 260992 180582 261004
rect 197998 260992 198004 261004
rect 198056 260992 198062 261044
rect 4798 260924 4804 260976
rect 4856 260964 4862 260976
rect 176194 260964 176200 260976
rect 4856 260936 176200 260964
rect 4856 260924 4862 260936
rect 176194 260924 176200 260936
rect 176252 260924 176258 260976
rect 184750 260924 184756 260976
rect 184808 260964 184814 260976
rect 197078 260964 197084 260976
rect 184808 260936 197084 260964
rect 184808 260924 184814 260936
rect 197078 260924 197084 260936
rect 197136 260924 197142 260976
rect 112622 260856 112628 260908
rect 112680 260896 112686 260908
rect 130378 260896 130384 260908
rect 112680 260868 130384 260896
rect 112680 260856 112686 260868
rect 130378 260856 130384 260868
rect 130436 260856 130442 260908
rect 181990 260856 181996 260908
rect 182048 260896 182054 260908
rect 197814 260896 197820 260908
rect 182048 260868 197820 260896
rect 182048 260856 182054 260868
rect 197814 260856 197820 260868
rect 197872 260856 197878 260908
rect 119890 260788 119896 260840
rect 119948 260828 119954 260840
rect 124306 260828 124312 260840
rect 119948 260800 124312 260828
rect 119948 260788 119954 260800
rect 124306 260788 124312 260800
rect 124364 260788 124370 260840
rect 119246 260720 119252 260772
rect 119304 260760 119310 260772
rect 122834 260760 122840 260772
rect 119304 260732 122840 260760
rect 119304 260720 119310 260732
rect 122834 260720 122840 260732
rect 122892 260720 122898 260772
rect 122742 260652 122748 260704
rect 122800 260692 122806 260704
rect 123202 260692 123208 260704
rect 122800 260664 123208 260692
rect 122800 260652 122806 260664
rect 123202 260652 123208 260664
rect 123260 260652 123266 260704
rect 180794 260516 180800 260568
rect 180852 260556 180858 260568
rect 189534 260556 189540 260568
rect 180852 260528 189540 260556
rect 180852 260516 180858 260528
rect 189534 260516 189540 260528
rect 189592 260516 189598 260568
rect 173894 260448 173900 260500
rect 173952 260488 173958 260500
rect 185578 260488 185584 260500
rect 173952 260460 185584 260488
rect 173952 260448 173958 260460
rect 185578 260448 185584 260460
rect 185636 260448 185642 260500
rect 133230 260380 133236 260432
rect 133288 260420 133294 260432
rect 485038 260420 485044 260432
rect 133288 260392 485044 260420
rect 133288 260380 133294 260392
rect 485038 260380 485044 260392
rect 485096 260380 485102 260432
rect 7558 260312 7564 260364
rect 7616 260352 7622 260364
rect 177298 260352 177304 260364
rect 7616 260324 177304 260352
rect 7616 260312 7622 260324
rect 177298 260312 177304 260324
rect 177356 260312 177362 260364
rect 192294 260352 192300 260364
rect 180766 260324 192300 260352
rect 114186 260244 114192 260296
rect 114244 260284 114250 260296
rect 126514 260284 126520 260296
rect 114244 260256 126520 260284
rect 114244 260244 114250 260256
rect 126514 260244 126520 260256
rect 126572 260244 126578 260296
rect 132466 260256 139532 260284
rect 118142 260176 118148 260228
rect 118200 260216 118206 260228
rect 132466 260216 132494 260256
rect 139504 260228 139532 260256
rect 164234 260244 164240 260296
rect 164292 260284 164298 260296
rect 175826 260284 175832 260296
rect 164292 260256 175832 260284
rect 164292 260244 164298 260256
rect 175826 260244 175832 260256
rect 175884 260244 175890 260296
rect 118200 260188 132494 260216
rect 118200 260176 118206 260188
rect 135254 260176 135260 260228
rect 135312 260216 135318 260228
rect 136220 260216 136226 260228
rect 135312 260188 136226 260216
rect 135312 260176 135318 260188
rect 136220 260176 136226 260188
rect 136278 260176 136284 260228
rect 139486 260176 139492 260228
rect 139544 260216 139550 260228
rect 140084 260216 140090 260228
rect 139544 260188 140090 260216
rect 139544 260176 139550 260188
rect 140084 260176 140090 260188
rect 140142 260176 140148 260228
rect 143534 260176 143540 260228
rect 143592 260216 143598 260228
rect 144500 260216 144506 260228
rect 143592 260188 144506 260216
rect 143592 260176 143598 260188
rect 144500 260176 144506 260188
rect 144558 260176 144564 260228
rect 155954 260176 155960 260228
rect 156012 260216 156018 260228
rect 156644 260216 156650 260228
rect 156012 260188 156650 260216
rect 156012 260176 156018 260188
rect 156644 260176 156650 260188
rect 156702 260176 156708 260228
rect 167270 260176 167276 260228
rect 167328 260216 167334 260228
rect 168236 260216 168242 260228
rect 167328 260188 168242 260216
rect 167328 260176 167334 260188
rect 168236 260176 168242 260188
rect 168294 260176 168300 260228
rect 169754 260176 169760 260228
rect 169812 260216 169818 260228
rect 170996 260216 171002 260228
rect 169812 260188 171002 260216
rect 169812 260176 169818 260188
rect 170996 260176 171002 260188
rect 171054 260176 171060 260228
rect 172514 260176 172520 260228
rect 172572 260216 172578 260228
rect 173204 260216 173210 260228
rect 172572 260188 173210 260216
rect 172572 260176 172578 260188
rect 173204 260176 173210 260188
rect 173262 260176 173268 260228
rect 175918 260176 175924 260228
rect 175976 260216 175982 260228
rect 180766 260216 180794 260324
rect 192294 260312 192300 260324
rect 192352 260312 192358 260364
rect 185578 260244 185584 260296
rect 185636 260284 185642 260296
rect 193858 260284 193864 260296
rect 185636 260256 193864 260284
rect 185636 260244 185642 260256
rect 193858 260244 193864 260256
rect 193916 260244 193922 260296
rect 191006 260216 191012 260228
rect 175976 260188 180794 260216
rect 180904 260188 191012 260216
rect 175976 260176 175982 260188
rect 113726 260108 113732 260160
rect 113784 260148 113790 260160
rect 139670 260148 139676 260160
rect 113784 260120 139676 260148
rect 113784 260108 113790 260120
rect 139670 260108 139676 260120
rect 139728 260148 139734 260160
rect 140636 260148 140642 260160
rect 139728 260120 140642 260148
rect 139728 260108 139734 260120
rect 140636 260108 140642 260120
rect 140694 260108 140700 260160
rect 166994 260108 167000 260160
rect 167052 260148 167058 260160
rect 167684 260148 167690 260160
rect 167052 260120 167690 260148
rect 167052 260108 167058 260120
rect 167684 260108 167690 260120
rect 167742 260148 167748 260160
rect 180794 260148 180800 260160
rect 167742 260120 180800 260148
rect 167742 260108 167748 260120
rect 180794 260108 180800 260120
rect 180852 260108 180858 260160
rect 118050 260040 118056 260092
rect 118108 260080 118114 260092
rect 135070 260080 135076 260092
rect 118108 260052 135076 260080
rect 118108 260040 118114 260052
rect 135070 260040 135076 260052
rect 135128 260040 135134 260092
rect 169340 260040 169346 260092
rect 169398 260080 169404 260092
rect 180904 260080 180932 260188
rect 191006 260176 191012 260188
rect 191064 260176 191070 260228
rect 189718 260148 189724 260160
rect 169398 260052 180932 260080
rect 183296 260120 189724 260148
rect 169398 260040 169404 260052
rect 112438 259972 112444 260024
rect 112496 260012 112502 260024
rect 132034 260012 132040 260024
rect 112496 259984 132040 260012
rect 112496 259972 112502 259984
rect 132034 259972 132040 259984
rect 132092 259972 132098 260024
rect 183296 260012 183324 260120
rect 189718 260108 189724 260120
rect 189776 260108 189782 260160
rect 189626 260080 189632 260092
rect 171520 259984 183324 260012
rect 183388 260052 189632 260080
rect 120626 259904 120632 259956
rect 120684 259944 120690 259956
rect 142154 259944 142160 259956
rect 120684 259916 142160 259944
rect 120684 259904 120690 259916
rect 142154 259904 142160 259916
rect 142212 259944 142218 259956
rect 143074 259944 143080 259956
rect 142212 259916 143080 259944
rect 142212 259904 142218 259916
rect 143074 259904 143080 259916
rect 143132 259904 143138 259956
rect 168374 259904 168380 259956
rect 168432 259944 168438 259956
rect 171520 259944 171548 259984
rect 183278 259944 183284 259956
rect 168432 259916 171548 259944
rect 171612 259916 183284 259944
rect 168432 259904 168438 259916
rect 119338 259836 119344 259888
rect 119396 259876 119402 259888
rect 143534 259876 143540 259888
rect 119396 259848 143540 259876
rect 119396 259836 119402 259848
rect 143534 259836 143540 259848
rect 143592 259836 143598 259888
rect 166166 259836 166172 259888
rect 166224 259876 166230 259888
rect 171612 259876 171640 259916
rect 183278 259904 183284 259916
rect 183336 259904 183342 259956
rect 166224 259848 171640 259876
rect 166224 259836 166230 259848
rect 175826 259836 175832 259888
rect 175884 259876 175890 259888
rect 183388 259876 183416 260052
rect 189626 260040 189632 260052
rect 189684 260040 189690 260092
rect 190914 260080 190920 260092
rect 190426 260052 190920 260080
rect 183462 259972 183468 260024
rect 183520 260012 183526 260024
rect 190426 260012 190454 260052
rect 190914 260040 190920 260052
rect 190972 260040 190978 260092
rect 183520 259984 190454 260012
rect 183520 259972 183526 259984
rect 192570 259944 192576 259956
rect 190426 259916 192576 259944
rect 175884 259848 183416 259876
rect 175884 259836 175890 259848
rect 183462 259836 183468 259888
rect 183520 259876 183526 259888
rect 190426 259876 190454 259916
rect 192570 259904 192576 259916
rect 192628 259904 192634 259956
rect 183520 259848 190454 259876
rect 183520 259836 183526 259848
rect 117866 259768 117872 259820
rect 117924 259808 117930 259820
rect 150434 259808 150440 259820
rect 117924 259780 150440 259808
rect 117924 259768 117930 259780
rect 150434 259768 150440 259780
rect 150492 259808 150498 259820
rect 151354 259808 151360 259820
rect 150492 259780 151360 259808
rect 150492 259768 150498 259780
rect 151354 259768 151360 259780
rect 151412 259768 151418 259820
rect 171134 259768 171140 259820
rect 171192 259808 171198 259820
rect 201862 259808 201868 259820
rect 171192 259780 201868 259808
rect 171192 259768 171198 259780
rect 201862 259768 201868 259780
rect 201920 259768 201926 259820
rect 115014 259700 115020 259752
rect 115072 259740 115078 259752
rect 149054 259740 149060 259752
rect 115072 259712 149060 259740
rect 115072 259700 115078 259712
rect 149054 259700 149060 259712
rect 149112 259740 149118 259752
rect 149698 259740 149704 259752
rect 149112 259712 149704 259740
rect 149112 259700 149118 259712
rect 149698 259700 149704 259712
rect 149756 259700 149762 259752
rect 156966 259700 156972 259752
rect 157024 259740 157030 259752
rect 185762 259740 185768 259752
rect 157024 259712 185768 259740
rect 157024 259700 157030 259712
rect 185762 259700 185768 259712
rect 185820 259700 185826 259752
rect 113818 259632 113824 259684
rect 113876 259672 113882 259684
rect 123754 259672 123760 259684
rect 113876 259644 123760 259672
rect 113876 259632 113882 259644
rect 123754 259632 123760 259644
rect 123812 259632 123818 259684
rect 134334 259632 134340 259684
rect 134392 259672 134398 259684
rect 187694 259672 187700 259684
rect 134392 259644 187700 259672
rect 134392 259632 134398 259644
rect 187694 259632 187700 259644
rect 187752 259632 187758 259684
rect 117774 259564 117780 259616
rect 117832 259604 117838 259616
rect 178034 259604 178040 259616
rect 117832 259576 178040 259604
rect 117832 259564 117838 259576
rect 178034 259564 178040 259576
rect 178092 259604 178098 259616
rect 196710 259604 196716 259616
rect 178092 259576 196716 259604
rect 178092 259564 178098 259576
rect 196710 259564 196716 259576
rect 196768 259564 196774 259616
rect 114094 259496 114100 259548
rect 114152 259536 114158 259548
rect 124858 259536 124864 259548
rect 114152 259508 124864 259536
rect 114152 259496 114158 259508
rect 124858 259496 124864 259508
rect 124916 259496 124922 259548
rect 173342 259496 173348 259548
rect 173400 259536 173406 259548
rect 201954 259536 201960 259548
rect 173400 259508 201960 259536
rect 173400 259496 173406 259508
rect 201954 259496 201960 259508
rect 202012 259496 202018 259548
rect 115198 259428 115204 259480
rect 115256 259468 115262 259480
rect 128354 259468 128360 259480
rect 115256 259440 128360 259468
rect 115256 259428 115262 259440
rect 128354 259428 128360 259440
rect 128412 259428 128418 259480
rect 185762 259428 185768 259480
rect 185820 259468 185826 259480
rect 190730 259468 190736 259480
rect 185820 259440 190736 259468
rect 185820 259428 185826 259440
rect 190730 259428 190736 259440
rect 190788 259428 190794 259480
rect 187694 259360 187700 259412
rect 187752 259400 187758 259412
rect 580166 259400 580172 259412
rect 187752 259372 580172 259400
rect 187752 259360 187758 259372
rect 580166 259360 580172 259372
rect 580224 259360 580230 259412
rect 485038 245556 485044 245608
rect 485096 245596 485102 245608
rect 580166 245596 580172 245608
rect 485096 245568 580172 245596
rect 485096 245556 485102 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 2774 241204 2780 241256
rect 2832 241244 2838 241256
rect 4798 241244 4804 241256
rect 2832 241216 4804 241244
rect 2832 241204 2838 241216
rect 4798 241204 4804 241216
rect 4856 241204 4862 241256
rect 3510 215092 3516 215144
rect 3568 215132 3574 215144
rect 7558 215132 7564 215144
rect 3568 215104 7564 215132
rect 3568 215092 3574 215104
rect 7558 215092 7564 215104
rect 7616 215092 7622 215144
rect 471238 206932 471244 206984
rect 471296 206972 471302 206984
rect 579798 206972 579804 206984
rect 471296 206944 579804 206972
rect 471296 206932 471302 206944
rect 579798 206932 579804 206944
rect 579856 206932 579862 206984
rect 146266 200892 149054 200920
rect 126256 200824 131114 200852
rect 126256 200728 126284 200824
rect 126238 200676 126244 200728
rect 126296 200676 126302 200728
rect 131086 200716 131114 200824
rect 132218 200716 132224 200728
rect 131086 200688 132224 200716
rect 132218 200676 132224 200688
rect 132276 200676 132282 200728
rect 128998 200648 129004 200660
rect 122806 200620 129004 200648
rect 107286 200540 107292 200592
rect 107344 200580 107350 200592
rect 122806 200580 122834 200620
rect 128998 200608 129004 200620
rect 129056 200608 129062 200660
rect 132144 200620 142154 200648
rect 107344 200552 122834 200580
rect 107344 200540 107350 200552
rect 128538 200540 128544 200592
rect 128596 200580 128602 200592
rect 131942 200580 131948 200592
rect 128596 200552 131948 200580
rect 128596 200540 128602 200552
rect 131942 200540 131948 200552
rect 132000 200540 132006 200592
rect 104802 200472 104808 200524
rect 104860 200512 104866 200524
rect 131574 200512 131580 200524
rect 104860 200484 131580 200512
rect 104860 200472 104866 200484
rect 131574 200472 131580 200484
rect 131632 200472 131638 200524
rect 132144 200444 132172 200620
rect 132218 200540 132224 200592
rect 132276 200580 132282 200592
rect 142126 200580 142154 200620
rect 143506 200620 144914 200648
rect 143506 200580 143534 200620
rect 132276 200552 140774 200580
rect 142126 200552 143534 200580
rect 144886 200580 144914 200620
rect 146266 200580 146294 200892
rect 149026 200852 149054 200892
rect 151878 200892 180104 200920
rect 149026 200824 149882 200852
rect 144886 200552 146294 200580
rect 132276 200540 132282 200552
rect 140746 200512 140774 200552
rect 140746 200484 143534 200512
rect 131086 200416 132172 200444
rect 121362 200336 121368 200388
rect 121420 200376 121426 200388
rect 131086 200376 131114 200416
rect 132218 200404 132224 200456
rect 132276 200444 132282 200456
rect 132276 200416 141004 200444
rect 132276 200404 132282 200416
rect 121420 200348 131114 200376
rect 121420 200336 121426 200348
rect 132034 200336 132040 200388
rect 132092 200376 132098 200388
rect 132092 200348 140912 200376
rect 132092 200336 132098 200348
rect 130286 200268 130292 200320
rect 130344 200308 130350 200320
rect 130344 200280 136542 200308
rect 130344 200268 130350 200280
rect 110230 200200 110236 200252
rect 110288 200240 110294 200252
rect 110288 200212 125594 200240
rect 110288 200200 110294 200212
rect 125566 199968 125594 200212
rect 127618 200200 127624 200252
rect 127676 200240 127682 200252
rect 132218 200240 132224 200252
rect 127676 200212 132224 200240
rect 127676 200200 127682 200212
rect 132218 200200 132224 200212
rect 132276 200200 132282 200252
rect 130470 200132 130476 200184
rect 130528 200172 130534 200184
rect 132034 200172 132040 200184
rect 130528 200144 132040 200172
rect 130528 200132 130534 200144
rect 132034 200132 132040 200144
rect 132092 200132 132098 200184
rect 131482 200064 131488 200116
rect 131540 200104 131546 200116
rect 136514 200104 136542 200280
rect 131540 200076 136358 200104
rect 136514 200076 139670 200104
rect 131540 200064 131546 200076
rect 130378 199996 130384 200048
rect 130436 200036 130442 200048
rect 131850 200036 131856 200048
rect 130436 200008 131856 200036
rect 130436 199996 130442 200008
rect 131850 199996 131856 200008
rect 131908 199996 131914 200048
rect 132218 199968 132224 199980
rect 125566 199940 132224 199968
rect 132218 199928 132224 199940
rect 132276 199928 132282 199980
rect 133846 199940 134518 199968
rect 119890 199860 119896 199912
rect 119948 199900 119954 199912
rect 125134 199900 125140 199912
rect 119948 199872 125140 199900
rect 119948 199860 119954 199872
rect 125134 199860 125140 199872
rect 125192 199860 125198 199912
rect 128354 199860 128360 199912
rect 128412 199900 128418 199912
rect 132632 199900 132638 199912
rect 128412 199872 132638 199900
rect 128412 199860 128418 199872
rect 132632 199860 132638 199872
rect 132690 199860 132696 199912
rect 132908 199860 132914 199912
rect 132966 199860 132972 199912
rect 133736 199860 133742 199912
rect 133794 199860 133800 199912
rect 127526 199792 127532 199844
rect 127584 199832 127590 199844
rect 132926 199832 132954 199860
rect 127584 199804 132954 199832
rect 127584 199792 127590 199804
rect 128998 199724 129004 199776
rect 129056 199764 129062 199776
rect 132954 199764 132960 199776
rect 129056 199736 132960 199764
rect 129056 199724 129062 199736
rect 132954 199724 132960 199736
rect 133012 199724 133018 199776
rect 111702 199656 111708 199708
rect 111760 199696 111766 199708
rect 130470 199696 130476 199708
rect 111760 199668 130476 199696
rect 111760 199656 111766 199668
rect 130470 199656 130476 199668
rect 130528 199656 130534 199708
rect 130562 199656 130568 199708
rect 130620 199696 130626 199708
rect 132310 199696 132316 199708
rect 130620 199668 132316 199696
rect 130620 199656 130626 199668
rect 132310 199656 132316 199668
rect 132368 199656 132374 199708
rect 133754 199696 133782 199860
rect 132420 199668 133782 199696
rect 109862 199588 109868 199640
rect 109920 199628 109926 199640
rect 130378 199628 130384 199640
rect 109920 199600 130384 199628
rect 109920 199588 109926 199600
rect 130378 199588 130384 199600
rect 130436 199588 130442 199640
rect 114462 199520 114468 199572
rect 114520 199560 114526 199572
rect 132310 199560 132316 199572
rect 114520 199532 132316 199560
rect 114520 199520 114526 199532
rect 132310 199520 132316 199532
rect 132368 199520 132374 199572
rect 114370 199452 114376 199504
rect 114428 199492 114434 199504
rect 114428 199464 126974 199492
rect 114428 199452 114434 199464
rect 126946 199424 126974 199464
rect 132218 199452 132224 199504
rect 132276 199492 132282 199504
rect 132420 199492 132448 199668
rect 133846 199640 133874 199940
rect 134490 199912 134518 199940
rect 136330 199912 136358 200076
rect 137250 200008 138566 200036
rect 137250 199912 137278 200008
rect 137480 199940 138474 199968
rect 133920 199860 133926 199912
rect 133978 199860 133984 199912
rect 134012 199860 134018 199912
rect 134070 199900 134076 199912
rect 134070 199860 134104 199900
rect 134196 199860 134202 199912
rect 134254 199860 134260 199912
rect 134288 199860 134294 199912
rect 134346 199860 134352 199912
rect 134472 199860 134478 199912
rect 134530 199860 134536 199912
rect 134564 199860 134570 199912
rect 134622 199860 134628 199912
rect 134656 199860 134662 199912
rect 134714 199860 134720 199912
rect 134840 199860 134846 199912
rect 134898 199860 134904 199912
rect 134932 199860 134938 199912
rect 134990 199860 134996 199912
rect 135116 199860 135122 199912
rect 135174 199860 135180 199912
rect 135300 199860 135306 199912
rect 135358 199860 135364 199912
rect 135484 199860 135490 199912
rect 135542 199900 135548 199912
rect 135542 199872 135622 199900
rect 135542 199860 135548 199872
rect 133782 199588 133788 199640
rect 133840 199600 133874 199640
rect 133840 199588 133846 199600
rect 132276 199464 132448 199492
rect 133938 199504 133966 199860
rect 134076 199640 134104 199860
rect 134214 199832 134242 199860
rect 134168 199804 134242 199832
rect 134168 199640 134196 199804
rect 134306 199708 134334 199860
rect 134242 199656 134248 199708
rect 134300 199668 134334 199708
rect 134582 199696 134610 199860
rect 134444 199668 134610 199696
rect 134300 199656 134306 199668
rect 134058 199588 134064 199640
rect 134116 199588 134122 199640
rect 134150 199588 134156 199640
rect 134208 199588 134214 199640
rect 134444 199628 134472 199668
rect 134260 199600 134472 199628
rect 133938 199464 133972 199504
rect 132276 199452 132282 199464
rect 133966 199452 133972 199464
rect 134024 199452 134030 199504
rect 132862 199424 132868 199436
rect 126946 199396 132868 199424
rect 132862 199384 132868 199396
rect 132920 199384 132926 199436
rect 132954 199384 132960 199436
rect 133012 199424 133018 199436
rect 133874 199424 133880 199436
rect 133012 199396 133880 199424
rect 133012 199384 133018 199396
rect 133874 199384 133880 199396
rect 133932 199384 133938 199436
rect 134260 199424 134288 199600
rect 134518 199588 134524 199640
rect 134576 199628 134582 199640
rect 134674 199628 134702 199860
rect 134858 199832 134886 199860
rect 134812 199804 134886 199832
rect 134812 199708 134840 199804
rect 134950 199776 134978 199860
rect 134886 199724 134892 199776
rect 134944 199736 134978 199776
rect 134944 199724 134950 199736
rect 134794 199656 134800 199708
rect 134852 199656 134858 199708
rect 134576 199600 134702 199628
rect 135134 199640 135162 199860
rect 135134 199600 135168 199640
rect 134576 199588 134582 199600
rect 135162 199588 135168 199600
rect 135220 199588 135226 199640
rect 135318 199628 135346 199860
rect 135318 199600 135392 199628
rect 135364 199572 135392 199600
rect 134334 199520 134340 199572
rect 134392 199560 134398 199572
rect 135254 199560 135260 199572
rect 134392 199532 135260 199560
rect 134392 199520 134398 199532
rect 135254 199520 135260 199532
rect 135312 199520 135318 199572
rect 135346 199520 135352 199572
rect 135404 199520 135410 199572
rect 135438 199520 135444 199572
rect 135496 199560 135502 199572
rect 135594 199560 135622 199872
rect 135668 199860 135674 199912
rect 135726 199860 135732 199912
rect 136036 199860 136042 199912
rect 136094 199860 136100 199912
rect 136220 199860 136226 199912
rect 136278 199860 136284 199912
rect 136312 199860 136318 199912
rect 136370 199860 136376 199912
rect 136680 199860 136686 199912
rect 136738 199900 136744 199912
rect 136738 199860 136772 199900
rect 137048 199860 137054 199912
rect 137106 199860 137112 199912
rect 137232 199860 137238 199912
rect 137290 199860 137296 199912
rect 137324 199860 137330 199912
rect 137382 199860 137388 199912
rect 135496 199532 135622 199560
rect 135686 199572 135714 199860
rect 135686 199532 135720 199572
rect 135496 199520 135502 199532
rect 135714 199520 135720 199532
rect 135772 199520 135778 199572
rect 136054 199504 136082 199860
rect 136238 199640 136266 199860
rect 136744 199640 136772 199860
rect 137066 199708 137094 199860
rect 137342 199776 137370 199860
rect 137278 199724 137284 199776
rect 137336 199736 137370 199776
rect 137336 199724 137342 199736
rect 137066 199668 137100 199708
rect 137094 199656 137100 199668
rect 137152 199656 137158 199708
rect 137480 199640 137508 199940
rect 138446 199912 138474 199940
rect 137600 199900 137606 199912
rect 137572 199860 137606 199900
rect 137658 199860 137664 199912
rect 137692 199860 137698 199912
rect 137750 199860 137756 199912
rect 137784 199860 137790 199912
rect 137842 199860 137848 199912
rect 137876 199860 137882 199912
rect 137934 199860 137940 199912
rect 138060 199860 138066 199912
rect 138118 199860 138124 199912
rect 138152 199860 138158 199912
rect 138210 199860 138216 199912
rect 138244 199860 138250 199912
rect 138302 199900 138308 199912
rect 138302 199860 138336 199900
rect 138428 199860 138434 199912
rect 138486 199860 138492 199912
rect 137572 199640 137600 199860
rect 137710 199832 137738 199860
rect 137664 199804 137738 199832
rect 137664 199776 137692 199804
rect 137802 199776 137830 199860
rect 137646 199724 137652 199776
rect 137704 199724 137710 199776
rect 137738 199724 137744 199776
rect 137796 199736 137830 199776
rect 137796 199724 137802 199736
rect 137894 199708 137922 199860
rect 138078 199776 138106 199860
rect 138170 199832 138198 199860
rect 138170 199804 138244 199832
rect 138216 199776 138244 199804
rect 138078 199736 138112 199776
rect 138106 199724 138112 199736
rect 138164 199724 138170 199776
rect 138198 199724 138204 199776
rect 138256 199724 138262 199776
rect 137830 199656 137836 199708
rect 137888 199668 137922 199708
rect 137888 199656 137894 199668
rect 136238 199600 136272 199640
rect 136266 199588 136272 199600
rect 136324 199588 136330 199640
rect 136726 199588 136732 199640
rect 136784 199588 136790 199640
rect 137462 199588 137468 199640
rect 137520 199588 137526 199640
rect 137554 199588 137560 199640
rect 137612 199588 137618 199640
rect 136634 199520 136640 199572
rect 136692 199560 136698 199572
rect 138308 199560 138336 199860
rect 138382 199724 138388 199776
rect 138440 199764 138446 199776
rect 138538 199764 138566 200008
rect 139642 199912 139670 200076
rect 140884 200036 140912 200348
rect 140976 200104 141004 200416
rect 143506 200172 143534 200484
rect 143506 200144 145006 200172
rect 140976 200076 144914 200104
rect 140884 200008 142430 200036
rect 140102 199940 140314 199968
rect 138612 199860 138618 199912
rect 138670 199860 138676 199912
rect 138980 199860 138986 199912
rect 139038 199860 139044 199912
rect 139348 199860 139354 199912
rect 139406 199860 139412 199912
rect 139440 199860 139446 199912
rect 139498 199900 139504 199912
rect 139498 199860 139532 199900
rect 139624 199860 139630 199912
rect 139682 199860 139688 199912
rect 139716 199860 139722 199912
rect 139774 199860 139780 199912
rect 138440 199736 138566 199764
rect 138440 199724 138446 199736
rect 138630 199708 138658 199860
rect 138998 199764 139026 199860
rect 138566 199656 138572 199708
rect 138624 199668 138658 199708
rect 138952 199736 139026 199764
rect 138624 199656 138630 199668
rect 138952 199640 138980 199736
rect 138934 199588 138940 199640
rect 138992 199588 138998 199640
rect 139366 199560 139394 199860
rect 139504 199708 139532 199860
rect 139486 199656 139492 199708
rect 139544 199656 139550 199708
rect 136692 199532 138336 199560
rect 138400 199532 139394 199560
rect 139734 199572 139762 199860
rect 139808 199792 139814 199844
rect 139866 199832 139872 199844
rect 139992 199832 139998 199844
rect 139866 199792 139900 199832
rect 139872 199708 139900 199792
rect 139964 199792 139998 199832
rect 140050 199792 140056 199844
rect 139964 199708 139992 199792
rect 139854 199656 139860 199708
rect 139912 199656 139918 199708
rect 139946 199656 139952 199708
rect 140004 199656 140010 199708
rect 140102 199572 140130 199940
rect 140286 199912 140314 199940
rect 141758 199940 141970 199968
rect 141758 199912 141786 199940
rect 140268 199860 140274 199912
rect 140326 199860 140332 199912
rect 140452 199860 140458 199912
rect 140510 199860 140516 199912
rect 140544 199860 140550 199912
rect 140602 199860 140608 199912
rect 140820 199900 140826 199912
rect 140792 199860 140826 199900
rect 140878 199860 140884 199912
rect 141004 199860 141010 199912
rect 141062 199860 141068 199912
rect 141096 199860 141102 199912
rect 141154 199860 141160 199912
rect 141280 199860 141286 199912
rect 141338 199860 141344 199912
rect 141372 199860 141378 199912
rect 141430 199860 141436 199912
rect 141740 199860 141746 199912
rect 141798 199860 141804 199912
rect 141832 199860 141838 199912
rect 141890 199860 141896 199912
rect 140176 199656 140182 199708
rect 140234 199696 140240 199708
rect 140234 199656 140268 199696
rect 139734 199532 139768 199572
rect 136692 199520 136698 199532
rect 134628 199464 135852 199492
rect 134628 199436 134656 199464
rect 134426 199424 134432 199436
rect 134260 199396 134432 199424
rect 134426 199384 134432 199396
rect 134484 199384 134490 199436
rect 134610 199384 134616 199436
rect 134668 199384 134674 199436
rect 135824 199424 135852 199464
rect 135990 199452 135996 199504
rect 136048 199464 136082 199504
rect 136048 199452 136054 199464
rect 138014 199452 138020 199504
rect 138072 199492 138078 199504
rect 138400 199492 138428 199532
rect 139762 199520 139768 199532
rect 139820 199520 139826 199572
rect 140102 199532 140136 199572
rect 140130 199520 140136 199532
rect 140188 199520 140194 199572
rect 138072 199464 138428 199492
rect 138072 199452 138078 199464
rect 138750 199452 138756 199504
rect 138808 199492 138814 199504
rect 139026 199492 139032 199504
rect 138808 199464 139032 199492
rect 138808 199452 138814 199464
rect 139026 199452 139032 199464
rect 139084 199452 139090 199504
rect 139118 199452 139124 199504
rect 139176 199492 139182 199504
rect 140240 199492 140268 199656
rect 140470 199628 140498 199860
rect 140562 199832 140590 199860
rect 140562 199804 140728 199832
rect 140590 199628 140596 199640
rect 140470 199600 140596 199628
rect 140590 199588 140596 199600
rect 140648 199588 140654 199640
rect 140406 199520 140412 199572
rect 140464 199560 140470 199572
rect 140700 199560 140728 199804
rect 140792 199640 140820 199860
rect 140866 199724 140872 199776
rect 140924 199764 140930 199776
rect 141022 199764 141050 199860
rect 140924 199736 141050 199764
rect 141114 199776 141142 199860
rect 141114 199736 141148 199776
rect 140924 199724 140930 199736
rect 141142 199724 141148 199736
rect 141200 199724 141206 199776
rect 141298 199696 141326 199860
rect 141160 199668 141326 199696
rect 140774 199588 140780 199640
rect 140832 199588 140838 199640
rect 140464 199532 140728 199560
rect 140464 199520 140470 199532
rect 139176 199464 140268 199492
rect 141160 199492 141188 199668
rect 141234 199520 141240 199572
rect 141292 199560 141298 199572
rect 141390 199560 141418 199860
rect 141464 199724 141470 199776
rect 141522 199764 141528 199776
rect 141522 199724 141556 199764
rect 141528 199640 141556 199724
rect 141850 199696 141878 199860
rect 141620 199668 141878 199696
rect 141510 199588 141516 199640
rect 141568 199588 141574 199640
rect 141292 199532 141418 199560
rect 141292 199520 141298 199532
rect 141326 199492 141332 199504
rect 141160 199464 141332 199492
rect 139176 199452 139182 199464
rect 141326 199452 141332 199464
rect 141384 199452 141390 199504
rect 141418 199452 141424 199504
rect 141476 199492 141482 199504
rect 141620 199492 141648 199668
rect 141476 199464 141648 199492
rect 141476 199452 141482 199464
rect 141786 199452 141792 199504
rect 141844 199492 141850 199504
rect 141942 199492 141970 199940
rect 142402 199912 142430 200008
rect 142016 199860 142022 199912
rect 142074 199860 142080 199912
rect 142384 199860 142390 199912
rect 142442 199860 142448 199912
rect 143212 199860 143218 199912
rect 143270 199860 143276 199912
rect 144500 199900 144506 199912
rect 144380 199872 144506 199900
rect 142034 199708 142062 199860
rect 142936 199792 142942 199844
rect 142994 199792 143000 199844
rect 142016 199656 142022 199708
rect 142074 199656 142080 199708
rect 142954 199572 142982 199792
rect 143230 199572 143258 199860
rect 143764 199832 143770 199844
rect 143460 199804 143770 199832
rect 142954 199532 142988 199572
rect 142982 199520 142988 199532
rect 143040 199520 143046 199572
rect 143230 199532 143264 199572
rect 143258 199520 143264 199532
rect 143316 199520 143322 199572
rect 141844 199464 141970 199492
rect 143460 199492 143488 199804
rect 143764 199792 143770 199804
rect 143822 199792 143828 199844
rect 143856 199792 143862 199844
rect 143914 199792 143920 199844
rect 143948 199792 143954 199844
rect 144006 199792 144012 199844
rect 144132 199832 144138 199844
rect 144104 199792 144138 199832
rect 144190 199792 144196 199844
rect 143874 199764 143902 199792
rect 143690 199736 143902 199764
rect 143580 199696 143586 199708
rect 143552 199656 143586 199696
rect 143638 199656 143644 199708
rect 143552 199572 143580 199656
rect 143690 199572 143718 199736
rect 143966 199708 143994 199792
rect 144104 199708 144132 199792
rect 143902 199656 143908 199708
rect 143960 199668 143994 199708
rect 143960 199656 143966 199668
rect 144086 199656 144092 199708
rect 144144 199656 144150 199708
rect 144380 199640 144408 199872
rect 144500 199860 144506 199872
rect 144558 199860 144564 199912
rect 144592 199860 144598 199912
rect 144650 199860 144656 199912
rect 144684 199860 144690 199912
rect 144742 199860 144748 199912
rect 144776 199860 144782 199912
rect 144834 199860 144840 199912
rect 144610 199832 144638 199860
rect 144564 199804 144638 199832
rect 144564 199708 144592 199804
rect 144702 199764 144730 199860
rect 144656 199736 144730 199764
rect 144656 199708 144684 199736
rect 144794 199708 144822 199860
rect 144546 199656 144552 199708
rect 144604 199656 144610 199708
rect 144638 199656 144644 199708
rect 144696 199656 144702 199708
rect 144730 199656 144736 199708
rect 144788 199668 144822 199708
rect 144886 199696 144914 200076
rect 144978 199912 145006 200144
rect 145162 200008 147674 200036
rect 144960 199860 144966 199912
rect 145018 199860 145024 199912
rect 145052 199860 145058 199912
rect 145110 199860 145116 199912
rect 145070 199776 145098 199860
rect 145006 199724 145012 199776
rect 145064 199736 145098 199776
rect 145064 199724 145070 199736
rect 145162 199696 145190 200008
rect 145346 199940 145834 199968
rect 145346 199776 145374 199940
rect 145696 199860 145702 199912
rect 145754 199860 145760 199912
rect 145328 199724 145334 199776
rect 145386 199724 145392 199776
rect 144886 199668 145190 199696
rect 144788 199656 144794 199668
rect 144362 199588 144368 199640
rect 144420 199588 144426 199640
rect 144822 199588 144828 199640
rect 144880 199628 144886 199640
rect 145714 199628 145742 199860
rect 144880 199600 145742 199628
rect 144880 199588 144886 199600
rect 143534 199520 143540 199572
rect 143592 199520 143598 199572
rect 143626 199520 143632 199572
rect 143684 199532 143718 199572
rect 143684 199520 143690 199532
rect 145282 199520 145288 199572
rect 145340 199560 145346 199572
rect 145806 199560 145834 199940
rect 146174 199940 146386 199968
rect 146174 199912 146202 199940
rect 145880 199860 145886 199912
rect 145938 199860 145944 199912
rect 146064 199900 146070 199912
rect 146036 199860 146070 199900
rect 146122 199860 146128 199912
rect 146156 199860 146162 199912
rect 146214 199860 146220 199912
rect 146248 199860 146254 199912
rect 146306 199860 146312 199912
rect 145340 199532 145834 199560
rect 145340 199520 145346 199532
rect 143810 199492 143816 199504
rect 143460 199464 143816 199492
rect 141844 199452 141850 199464
rect 143810 199452 143816 199464
rect 143868 199452 143874 199504
rect 137002 199424 137008 199436
rect 135824 199396 137008 199424
rect 137002 199384 137008 199396
rect 137060 199384 137066 199436
rect 137186 199384 137192 199436
rect 137244 199424 137250 199436
rect 144270 199424 144276 199436
rect 137244 199396 144276 199424
rect 137244 199384 137250 199396
rect 144270 199384 144276 199396
rect 144328 199384 144334 199436
rect 145650 199384 145656 199436
rect 145708 199424 145714 199436
rect 145898 199424 145926 199860
rect 146036 199640 146064 199860
rect 146266 199776 146294 199860
rect 146202 199724 146208 199776
rect 146260 199736 146294 199776
rect 146260 199724 146266 199736
rect 146018 199588 146024 199640
rect 146076 199588 146082 199640
rect 146358 199504 146386 199940
rect 146432 199860 146438 199912
rect 146490 199860 146496 199912
rect 146800 199860 146806 199912
rect 146858 199860 146864 199912
rect 146984 199860 146990 199912
rect 147042 199860 147048 199912
rect 147536 199860 147542 199912
rect 147594 199860 147600 199912
rect 146450 199776 146478 199860
rect 146450 199736 146484 199776
rect 146478 199724 146484 199736
rect 146536 199724 146542 199776
rect 146818 199696 146846 199860
rect 146294 199452 146300 199504
rect 146352 199464 146386 199504
rect 146450 199668 146846 199696
rect 146352 199452 146358 199464
rect 145708 199396 145926 199424
rect 145708 199384 145714 199396
rect 146110 199384 146116 199436
rect 146168 199424 146174 199436
rect 146450 199424 146478 199668
rect 146754 199588 146760 199640
rect 146812 199628 146818 199640
rect 147002 199628 147030 199860
rect 147554 199776 147582 199860
rect 147646 199832 147674 200008
rect 148888 199940 149146 199968
rect 147812 199832 147818 199844
rect 147646 199804 147818 199832
rect 147812 199792 147818 199804
rect 147870 199792 147876 199844
rect 148456 199792 148462 199844
rect 148514 199792 148520 199844
rect 148640 199832 148646 199844
rect 148612 199792 148646 199832
rect 148698 199792 148704 199844
rect 147490 199724 147496 199776
rect 147548 199736 147582 199776
rect 147548 199724 147554 199736
rect 147582 199656 147588 199708
rect 147640 199696 147646 199708
rect 148364 199696 148370 199708
rect 147640 199668 148370 199696
rect 147640 199656 147646 199668
rect 148364 199656 148370 199668
rect 148422 199656 148428 199708
rect 146812 199600 147030 199628
rect 146812 199588 146818 199600
rect 147306 199588 147312 199640
rect 147364 199628 147370 199640
rect 147364 199600 147674 199628
rect 147364 199588 147370 199600
rect 147646 199560 147674 199600
rect 148474 199560 148502 199792
rect 148612 199708 148640 199792
rect 148594 199656 148600 199708
rect 148652 199656 148658 199708
rect 147646 199532 148502 199560
rect 148888 199492 148916 199940
rect 149118 199912 149146 199940
rect 149854 199912 149882 200824
rect 151878 199968 151906 200892
rect 149946 199940 151078 199968
rect 149100 199860 149106 199912
rect 149158 199860 149164 199912
rect 149192 199860 149198 199912
rect 149250 199860 149256 199912
rect 149468 199860 149474 199912
rect 149526 199860 149532 199912
rect 149836 199860 149842 199912
rect 149894 199860 149900 199912
rect 149210 199708 149238 199860
rect 149146 199656 149152 199708
rect 149204 199668 149238 199708
rect 149486 199696 149514 199860
rect 149652 199792 149658 199844
rect 149710 199832 149716 199844
rect 149710 199792 149744 199832
rect 149486 199668 149652 199696
rect 149204 199656 149210 199668
rect 149624 199640 149652 199668
rect 149606 199588 149612 199640
rect 149664 199588 149670 199640
rect 149422 199520 149428 199572
rect 149480 199560 149486 199572
rect 149716 199560 149744 199792
rect 149480 199532 149744 199560
rect 149480 199520 149486 199532
rect 149054 199492 149060 199504
rect 148888 199464 149060 199492
rect 149054 199452 149060 199464
rect 149112 199452 149118 199504
rect 146168 199396 146478 199424
rect 146168 199384 146174 199396
rect 148318 199384 148324 199436
rect 148376 199424 148382 199436
rect 149946 199424 149974 199940
rect 151050 199912 151078 199940
rect 151786 199940 151906 199968
rect 151970 200824 155586 200852
rect 150020 199860 150026 199912
rect 150078 199860 150084 199912
rect 150204 199860 150210 199912
rect 150262 199860 150268 199912
rect 150480 199860 150486 199912
rect 150538 199860 150544 199912
rect 150572 199860 150578 199912
rect 150630 199860 150636 199912
rect 150664 199860 150670 199912
rect 150722 199860 150728 199912
rect 150940 199860 150946 199912
rect 150998 199860 151004 199912
rect 151032 199860 151038 199912
rect 151090 199860 151096 199912
rect 151216 199860 151222 199912
rect 151274 199860 151280 199912
rect 151308 199860 151314 199912
rect 151366 199860 151372 199912
rect 151400 199860 151406 199912
rect 151458 199860 151464 199912
rect 151676 199860 151682 199912
rect 151734 199860 151740 199912
rect 150038 199572 150066 199860
rect 150222 199832 150250 199860
rect 150176 199804 150250 199832
rect 150176 199640 150204 199804
rect 150296 199792 150302 199844
rect 150354 199792 150360 199844
rect 150498 199832 150526 199860
rect 150452 199804 150526 199832
rect 150314 199708 150342 199792
rect 150452 199776 150480 199804
rect 150590 199776 150618 199860
rect 150434 199724 150440 199776
rect 150492 199724 150498 199776
rect 150526 199724 150532 199776
rect 150584 199736 150618 199776
rect 150682 199764 150710 199860
rect 150848 199832 150854 199844
rect 150820 199792 150854 199832
rect 150906 199792 150912 199844
rect 150682 199736 150756 199764
rect 150584 199724 150590 199736
rect 150728 199708 150756 199736
rect 150820 199708 150848 199792
rect 150250 199656 150256 199708
rect 150308 199668 150342 199708
rect 150308 199656 150314 199668
rect 150710 199656 150716 199708
rect 150768 199656 150774 199708
rect 150802 199656 150808 199708
rect 150860 199656 150866 199708
rect 150158 199588 150164 199640
rect 150216 199588 150222 199640
rect 150038 199532 150072 199572
rect 150066 199520 150072 199532
rect 150124 199520 150130 199572
rect 150958 199560 150986 199860
rect 151234 199764 151262 199860
rect 151096 199736 151262 199764
rect 151096 199640 151124 199736
rect 151078 199588 151084 199640
rect 151136 199588 151142 199640
rect 151170 199588 151176 199640
rect 151228 199628 151234 199640
rect 151326 199628 151354 199860
rect 151418 199776 151446 199860
rect 151418 199736 151452 199776
rect 151446 199724 151452 199736
rect 151504 199724 151510 199776
rect 151694 199640 151722 199860
rect 151228 199600 151354 199628
rect 151228 199588 151234 199600
rect 151630 199588 151636 199640
rect 151688 199600 151722 199640
rect 151688 199588 151694 199600
rect 151262 199560 151268 199572
rect 150958 199532 151268 199560
rect 151262 199520 151268 199532
rect 151320 199520 151326 199572
rect 151786 199492 151814 199940
rect 151860 199860 151866 199912
rect 151918 199860 151924 199912
rect 151878 199708 151906 199860
rect 151970 199764 151998 200824
rect 152062 200756 155034 200784
rect 152062 199912 152090 200756
rect 152568 199940 153470 199968
rect 152044 199860 152050 199912
rect 152102 199860 152108 199912
rect 152136 199860 152142 199912
rect 152194 199860 152200 199912
rect 152228 199860 152234 199912
rect 152286 199860 152292 199912
rect 152154 199764 152182 199860
rect 151970 199736 152044 199764
rect 151878 199668 151912 199708
rect 151906 199656 151912 199668
rect 151964 199656 151970 199708
rect 152016 199560 152044 199736
rect 152108 199736 152182 199764
rect 152108 199708 152136 199736
rect 152246 199708 152274 199860
rect 152412 199792 152418 199844
rect 152470 199792 152476 199844
rect 152090 199656 152096 199708
rect 152148 199656 152154 199708
rect 152182 199656 152188 199708
rect 152240 199668 152274 199708
rect 152240 199656 152246 199668
rect 152430 199640 152458 199792
rect 152366 199588 152372 199640
rect 152424 199600 152458 199640
rect 152424 199588 152430 199600
rect 152568 199560 152596 199940
rect 153442 199912 153470 199940
rect 152688 199860 152694 199912
rect 152746 199860 152752 199912
rect 152780 199860 152786 199912
rect 152838 199860 152844 199912
rect 152964 199860 152970 199912
rect 153022 199860 153028 199912
rect 153056 199860 153062 199912
rect 153114 199860 153120 199912
rect 153148 199860 153154 199912
rect 153206 199900 153212 199912
rect 153206 199860 153240 199900
rect 153332 199860 153338 199912
rect 153390 199860 153396 199912
rect 153424 199860 153430 199912
rect 153482 199860 153488 199912
rect 153608 199860 153614 199912
rect 153666 199860 153672 199912
rect 153700 199860 153706 199912
rect 153758 199860 153764 199912
rect 153976 199900 153982 199912
rect 153810 199872 153982 199900
rect 152706 199832 152734 199860
rect 152660 199804 152734 199832
rect 152660 199628 152688 199804
rect 152798 199776 152826 199860
rect 152734 199724 152740 199776
rect 152792 199736 152826 199776
rect 152982 199776 153010 199860
rect 153074 199832 153102 199860
rect 153074 199804 153148 199832
rect 153120 199776 153148 199804
rect 153212 199776 153240 199860
rect 153350 199776 153378 199860
rect 153626 199832 153654 199860
rect 153580 199804 153654 199832
rect 153580 199776 153608 199804
rect 152982 199736 153016 199776
rect 152792 199724 152798 199736
rect 153010 199724 153016 199736
rect 153068 199724 153074 199776
rect 153102 199724 153108 199776
rect 153160 199724 153166 199776
rect 153194 199724 153200 199776
rect 153252 199724 153258 199776
rect 153350 199736 153384 199776
rect 153378 199724 153384 199736
rect 153436 199724 153442 199776
rect 153562 199724 153568 199776
rect 153620 199724 153626 199776
rect 153470 199656 153476 199708
rect 153528 199696 153534 199708
rect 153718 199696 153746 199860
rect 153528 199668 153746 199696
rect 153528 199656 153534 199668
rect 152918 199628 152924 199640
rect 152660 199600 152924 199628
rect 152918 199588 152924 199600
rect 152976 199588 152982 199640
rect 153654 199588 153660 199640
rect 153712 199628 153718 199640
rect 153810 199628 153838 199872
rect 153976 199860 153982 199872
rect 154034 199860 154040 199912
rect 154068 199860 154074 199912
rect 154126 199860 154132 199912
rect 154160 199860 154166 199912
rect 154218 199860 154224 199912
rect 154252 199860 154258 199912
rect 154310 199860 154316 199912
rect 154436 199860 154442 199912
rect 154494 199860 154500 199912
rect 154086 199708 154114 199860
rect 154022 199656 154028 199708
rect 154080 199668 154114 199708
rect 154080 199656 154086 199668
rect 153712 199600 153838 199628
rect 154178 199640 154206 199860
rect 154270 199696 154298 199860
rect 154270 199668 154344 199696
rect 154178 199600 154212 199640
rect 153712 199588 153718 199600
rect 154206 199588 154212 199600
rect 154264 199588 154270 199640
rect 152016 199532 152596 199560
rect 154114 199520 154120 199572
rect 154172 199560 154178 199572
rect 154316 199560 154344 199668
rect 154454 199572 154482 199860
rect 154620 199832 154626 199844
rect 154546 199804 154626 199832
rect 154546 199640 154574 199804
rect 154620 199792 154626 199804
rect 154678 199792 154684 199844
rect 154712 199792 154718 199844
rect 154770 199792 154776 199844
rect 155006 199832 155034 200756
rect 155080 199860 155086 199912
rect 155138 199900 155144 199912
rect 155138 199872 155264 199900
rect 155138 199860 155144 199872
rect 155006 199804 155080 199832
rect 154528 199588 154534 199640
rect 154586 199588 154592 199640
rect 154172 199532 154344 199560
rect 154172 199520 154178 199532
rect 154390 199520 154396 199572
rect 154448 199532 154482 199572
rect 154730 199560 154758 199792
rect 154942 199560 154948 199572
rect 154730 199532 154948 199560
rect 154448 199520 154454 199532
rect 154942 199520 154948 199532
rect 155000 199520 155006 199572
rect 154666 199492 154672 199504
rect 151786 199464 154672 199492
rect 154666 199452 154672 199464
rect 154724 199452 154730 199504
rect 154850 199452 154856 199504
rect 154908 199492 154914 199504
rect 155052 199492 155080 199804
rect 154908 199464 155080 199492
rect 155236 199492 155264 199872
rect 155356 199832 155362 199844
rect 155328 199792 155362 199832
rect 155414 199792 155420 199844
rect 155328 199572 155356 199792
rect 155558 199696 155586 200824
rect 160066 200824 177804 200852
rect 160066 200104 160094 200824
rect 177776 200728 177804 200824
rect 179386 200756 180012 200784
rect 172578 200688 173710 200716
rect 172578 200648 172606 200688
rect 170232 200620 172422 200648
rect 165816 200416 168374 200444
rect 165816 200376 165844 200416
rect 159238 200076 160094 200104
rect 162826 200348 165844 200376
rect 168346 200376 168374 200416
rect 168346 200348 168788 200376
rect 158686 200008 159174 200036
rect 156294 199940 157196 199968
rect 156294 199844 156322 199940
rect 156552 199860 156558 199912
rect 156610 199860 156616 199912
rect 155632 199792 155638 199844
rect 155690 199832 155696 199844
rect 155690 199792 155724 199832
rect 155816 199792 155822 199844
rect 155874 199832 155880 199844
rect 155874 199792 155908 199832
rect 156000 199792 156006 199844
rect 156058 199792 156064 199844
rect 156184 199792 156190 199844
rect 156242 199792 156248 199844
rect 156276 199792 156282 199844
rect 156334 199792 156340 199844
rect 155696 199708 155724 199792
rect 155880 199708 155908 199792
rect 156018 199708 156046 199792
rect 156202 199708 156230 199792
rect 156570 199764 156598 199860
rect 156920 199764 156926 199776
rect 156524 199736 156598 199764
rect 155558 199668 155632 199696
rect 155604 199640 155632 199668
rect 155678 199656 155684 199708
rect 155736 199656 155742 199708
rect 155862 199656 155868 199708
rect 155920 199656 155926 199708
rect 156018 199668 156052 199708
rect 156046 199656 156052 199668
rect 156104 199656 156110 199708
rect 156202 199668 156236 199708
rect 156230 199656 156236 199668
rect 156288 199656 156294 199708
rect 156524 199640 156552 199736
rect 156892 199724 156926 199764
rect 156978 199724 156984 199776
rect 156892 199640 156920 199724
rect 157168 199640 157196 199940
rect 157398 199940 157610 199968
rect 157398 199844 157426 199940
rect 157472 199860 157478 199912
rect 157530 199860 157536 199912
rect 157288 199792 157294 199844
rect 157346 199792 157352 199844
rect 157380 199792 157386 199844
rect 157438 199792 157444 199844
rect 157306 199640 157334 199792
rect 157490 199708 157518 199860
rect 157426 199656 157432 199708
rect 157484 199668 157518 199708
rect 157484 199656 157490 199668
rect 155586 199588 155592 199640
rect 155644 199588 155650 199640
rect 156506 199588 156512 199640
rect 156564 199588 156570 199640
rect 156874 199588 156880 199640
rect 156932 199588 156938 199640
rect 157150 199588 157156 199640
rect 157208 199588 157214 199640
rect 157306 199600 157340 199640
rect 157334 199588 157340 199600
rect 157392 199588 157398 199640
rect 155310 199520 155316 199572
rect 155368 199520 155374 199572
rect 157582 199560 157610 199940
rect 158686 199912 158714 200008
rect 157656 199860 157662 199912
rect 157714 199860 157720 199912
rect 158116 199860 158122 199912
rect 158174 199860 158180 199912
rect 158484 199860 158490 199912
rect 158542 199860 158548 199912
rect 158668 199860 158674 199912
rect 158726 199860 158732 199912
rect 157674 199708 157702 199860
rect 158134 199832 158162 199860
rect 157858 199804 158162 199832
rect 157674 199668 157708 199708
rect 157702 199656 157708 199668
rect 157760 199656 157766 199708
rect 157536 199532 157610 199560
rect 157858 199572 157886 199804
rect 157932 199724 157938 199776
rect 157990 199764 157996 199776
rect 158116 199764 158122 199776
rect 157990 199724 158024 199764
rect 157858 199532 157892 199572
rect 157536 199504 157564 199532
rect 157886 199520 157892 199532
rect 157944 199520 157950 199572
rect 157242 199492 157248 199504
rect 155236 199464 157248 199492
rect 154908 199452 154914 199464
rect 157242 199452 157248 199464
rect 157300 199452 157306 199504
rect 157518 199452 157524 199504
rect 157576 199452 157582 199504
rect 157610 199452 157616 199504
rect 157668 199492 157674 199504
rect 157996 199492 158024 199724
rect 158088 199724 158122 199764
rect 158174 199724 158180 199776
rect 158088 199572 158116 199724
rect 158502 199696 158530 199860
rect 158576 199792 158582 199844
rect 158634 199832 158640 199844
rect 158634 199792 158668 199832
rect 159036 199792 159042 199844
rect 159094 199792 159100 199844
rect 158456 199668 158530 199696
rect 158456 199640 158484 199668
rect 158438 199588 158444 199640
rect 158496 199588 158502 199640
rect 158530 199588 158536 199640
rect 158588 199628 158594 199640
rect 158640 199628 158668 199792
rect 158588 199600 158668 199628
rect 159054 199640 159082 199792
rect 159146 199696 159174 200008
rect 159238 199912 159266 200076
rect 159698 200008 160278 200036
rect 159698 199912 159726 200008
rect 159220 199860 159226 199912
rect 159278 199860 159284 199912
rect 159312 199860 159318 199912
rect 159370 199860 159376 199912
rect 159404 199860 159410 199912
rect 159462 199860 159468 199912
rect 159588 199860 159594 199912
rect 159646 199860 159652 199912
rect 159680 199860 159686 199912
rect 159738 199860 159744 199912
rect 160140 199860 160146 199912
rect 160198 199860 160204 199912
rect 159330 199776 159358 199860
rect 159266 199724 159272 199776
rect 159324 199736 159358 199776
rect 159324 199724 159330 199736
rect 159422 199708 159450 199860
rect 159146 199668 159312 199696
rect 159054 199600 159088 199640
rect 158588 199588 158594 199600
rect 159082 199588 159088 199600
rect 159140 199588 159146 199640
rect 159284 199628 159312 199668
rect 159358 199656 159364 199708
rect 159416 199668 159450 199708
rect 159606 199708 159634 199860
rect 160048 199832 160054 199844
rect 159744 199804 160054 199832
rect 159606 199668 159640 199708
rect 159416 199656 159422 199668
rect 159634 199656 159640 199668
rect 159692 199656 159698 199708
rect 159744 199640 159772 199804
rect 160048 199792 160054 199804
rect 160106 199792 160112 199844
rect 159542 199628 159548 199640
rect 159284 199600 159548 199628
rect 159542 199588 159548 199600
rect 159600 199588 159606 199640
rect 159726 199588 159732 199640
rect 159784 199588 159790 199640
rect 160158 199628 160186 199860
rect 159836 199600 160186 199628
rect 158070 199520 158076 199572
rect 158128 199520 158134 199572
rect 159450 199520 159456 199572
rect 159508 199560 159514 199572
rect 159836 199560 159864 199600
rect 160250 199572 160278 200008
rect 159508 199532 159864 199560
rect 159508 199520 159514 199532
rect 160186 199520 160192 199572
rect 160244 199532 160278 199572
rect 160388 200008 162670 200036
rect 160388 199560 160416 200008
rect 160802 199940 161290 199968
rect 160600 199860 160606 199912
rect 160658 199860 160664 199912
rect 160692 199860 160698 199912
rect 160750 199860 160756 199912
rect 160618 199832 160646 199860
rect 160480 199804 160646 199832
rect 160480 199628 160508 199804
rect 160554 199656 160560 199708
rect 160612 199696 160618 199708
rect 160710 199696 160738 199860
rect 160612 199668 160738 199696
rect 160802 199696 160830 199940
rect 161262 199912 161290 199940
rect 162642 199912 162670 200008
rect 160894 199872 161106 199900
rect 160894 199844 160922 199872
rect 160876 199792 160882 199844
rect 160934 199792 160940 199844
rect 160968 199792 160974 199844
rect 161026 199792 161032 199844
rect 160986 199708 161014 199792
rect 160802 199668 160876 199696
rect 160612 199656 160618 199668
rect 160738 199628 160744 199640
rect 160480 199600 160744 199628
rect 160738 199588 160744 199600
rect 160796 199588 160802 199640
rect 160646 199560 160652 199572
rect 160388 199532 160652 199560
rect 160244 199520 160250 199532
rect 160646 199520 160652 199532
rect 160704 199520 160710 199572
rect 160848 199560 160876 199668
rect 160922 199656 160928 199708
rect 160980 199668 161014 199708
rect 160980 199656 160986 199668
rect 161078 199628 161106 199872
rect 161152 199860 161158 199912
rect 161210 199860 161216 199912
rect 161244 199860 161250 199912
rect 161302 199860 161308 199912
rect 161428 199860 161434 199912
rect 161486 199860 161492 199912
rect 161520 199860 161526 199912
rect 161578 199860 161584 199912
rect 161704 199860 161710 199912
rect 161762 199860 161768 199912
rect 161796 199860 161802 199912
rect 161854 199860 161860 199912
rect 161888 199860 161894 199912
rect 161946 199860 161952 199912
rect 162164 199860 162170 199912
rect 162222 199860 162228 199912
rect 162348 199860 162354 199912
rect 162406 199860 162412 199912
rect 162440 199860 162446 199912
rect 162498 199860 162504 199912
rect 162532 199860 162538 199912
rect 162590 199860 162596 199912
rect 162624 199860 162630 199912
rect 162682 199860 162688 199912
rect 161170 199776 161198 199860
rect 161446 199832 161474 199860
rect 161400 199804 161474 199832
rect 161170 199736 161204 199776
rect 161198 199724 161204 199736
rect 161256 199724 161262 199776
rect 161400 199708 161428 199804
rect 161538 199776 161566 199860
rect 161722 199832 161750 199860
rect 161676 199804 161750 199832
rect 161676 199776 161704 199804
rect 161814 199776 161842 199860
rect 161474 199724 161480 199776
rect 161532 199736 161566 199776
rect 161532 199724 161538 199736
rect 161658 199724 161664 199776
rect 161716 199724 161722 199776
rect 161750 199724 161756 199776
rect 161808 199736 161842 199776
rect 161808 199724 161814 199736
rect 161906 199708 161934 199860
rect 162182 199708 162210 199860
rect 162366 199832 162394 199860
rect 162320 199804 162394 199832
rect 162320 199776 162348 199804
rect 162458 199776 162486 199860
rect 162302 199724 162308 199776
rect 162360 199724 162366 199776
rect 162394 199724 162400 199776
rect 162452 199736 162486 199776
rect 162452 199724 162458 199736
rect 161382 199656 161388 199708
rect 161440 199656 161446 199708
rect 161842 199656 161848 199708
rect 161900 199668 161934 199708
rect 161900 199656 161906 199668
rect 162118 199656 162124 199708
rect 162176 199668 162210 199708
rect 162550 199708 162578 199860
rect 162550 199668 162584 199708
rect 162176 199656 162182 199668
rect 162578 199656 162584 199668
rect 162636 199656 162642 199708
rect 161474 199628 161480 199640
rect 161078 199600 161480 199628
rect 161474 199588 161480 199600
rect 161532 199588 161538 199640
rect 161566 199588 161572 199640
rect 161624 199628 161630 199640
rect 162826 199628 162854 200348
rect 168760 200308 168788 200348
rect 161624 199600 162854 199628
rect 162918 200280 168696 200308
rect 168760 200280 169202 200308
rect 161624 199588 161630 199600
rect 161198 199560 161204 199572
rect 160848 199532 161204 199560
rect 161198 199520 161204 199532
rect 161256 199520 161262 199572
rect 157668 199464 158024 199492
rect 157668 199452 157674 199464
rect 162394 199452 162400 199504
rect 162452 199492 162458 199504
rect 162918 199492 162946 200280
rect 163102 200212 168052 200240
rect 162992 199860 162998 199912
rect 163050 199860 163056 199912
rect 162452 199464 162946 199492
rect 162452 199452 162458 199464
rect 148376 199396 149974 199424
rect 148376 199384 148382 199396
rect 156230 199384 156236 199436
rect 156288 199424 156294 199436
rect 160186 199424 160192 199436
rect 156288 199396 160192 199424
rect 156288 199384 156294 199396
rect 160186 199384 160192 199396
rect 160244 199384 160250 199436
rect 161382 199384 161388 199436
rect 161440 199424 161446 199436
rect 163010 199424 163038 199860
rect 161440 199396 163038 199424
rect 161440 199384 161446 199396
rect 118602 199316 118608 199368
rect 118660 199356 118666 199368
rect 145098 199356 145104 199368
rect 118660 199328 135254 199356
rect 118660 199316 118666 199328
rect 118418 199248 118424 199300
rect 118476 199288 118482 199300
rect 135070 199288 135076 199300
rect 118476 199260 135076 199288
rect 118476 199248 118482 199260
rect 135070 199248 135076 199260
rect 135128 199248 135134 199300
rect 135226 199288 135254 199328
rect 135318 199328 145104 199356
rect 135318 199288 135346 199328
rect 145098 199316 145104 199328
rect 145156 199316 145162 199368
rect 145190 199316 145196 199368
rect 145248 199356 145254 199368
rect 148410 199356 148416 199368
rect 145248 199328 148416 199356
rect 145248 199316 145254 199328
rect 148410 199316 148416 199328
rect 148468 199316 148474 199368
rect 150618 199316 150624 199368
rect 150676 199356 150682 199368
rect 150676 199328 154666 199356
rect 150676 199316 150682 199328
rect 135226 199260 135346 199288
rect 135714 199248 135720 199300
rect 135772 199288 135778 199300
rect 146202 199288 146208 199300
rect 135772 199260 146208 199288
rect 135772 199248 135778 199260
rect 146202 199248 146208 199260
rect 146260 199248 146266 199300
rect 149514 199248 149520 199300
rect 149572 199288 149578 199300
rect 154638 199288 154666 199328
rect 155466 199328 159404 199356
rect 155466 199288 155494 199328
rect 149572 199260 154574 199288
rect 154638 199260 155494 199288
rect 149572 199248 149578 199260
rect 117222 199180 117228 199232
rect 117280 199220 117286 199232
rect 145374 199220 145380 199232
rect 117280 199192 145380 199220
rect 117280 199180 117286 199192
rect 145374 199180 145380 199192
rect 145432 199180 145438 199232
rect 115750 199112 115756 199164
rect 115808 199152 115814 199164
rect 145926 199152 145932 199164
rect 115808 199124 145932 199152
rect 115808 199112 115814 199124
rect 145926 199112 145932 199124
rect 145984 199112 145990 199164
rect 154546 199152 154574 199260
rect 157794 199248 157800 199300
rect 157852 199288 157858 199300
rect 158714 199288 158720 199300
rect 157852 199260 158720 199288
rect 157852 199248 157858 199260
rect 158714 199248 158720 199260
rect 158772 199248 158778 199300
rect 159376 199288 159404 199328
rect 159542 199316 159548 199368
rect 159600 199356 159606 199368
rect 162026 199356 162032 199368
rect 159600 199328 162032 199356
rect 159600 199316 159606 199328
rect 162026 199316 162032 199328
rect 162084 199316 162090 199368
rect 162486 199316 162492 199368
rect 162544 199356 162550 199368
rect 163102 199356 163130 200212
rect 163194 200144 166948 200172
rect 163194 199504 163222 200144
rect 163516 200076 166028 200104
rect 163268 199860 163274 199912
rect 163326 199860 163332 199912
rect 163360 199860 163366 199912
rect 163418 199860 163424 199912
rect 163286 199776 163314 199860
rect 163268 199724 163274 199776
rect 163326 199724 163332 199776
rect 163378 199764 163406 199860
rect 163378 199736 163452 199764
rect 163424 199640 163452 199736
rect 163268 199588 163274 199640
rect 163326 199628 163332 199640
rect 163326 199588 163360 199628
rect 163406 199588 163412 199640
rect 163464 199588 163470 199640
rect 163194 199464 163228 199504
rect 163222 199452 163228 199464
rect 163280 199452 163286 199504
rect 163332 199436 163360 199588
rect 163314 199384 163320 199436
rect 163372 199384 163378 199436
rect 162544 199328 163130 199356
rect 162544 199316 162550 199328
rect 163516 199288 163544 200076
rect 163700 200008 164510 200036
rect 163700 199572 163728 200008
rect 163912 199860 163918 199912
rect 163970 199900 163976 199912
rect 163970 199872 164234 199900
rect 163970 199860 163976 199872
rect 163820 199792 163826 199844
rect 163878 199792 163884 199844
rect 163838 199708 163866 199792
rect 164206 199764 164234 199872
rect 164280 199860 164286 199912
rect 164338 199900 164344 199912
rect 164338 199860 164372 199900
rect 164344 199776 164372 199860
rect 164206 199736 164280 199764
rect 163838 199668 163872 199708
rect 163866 199656 163872 199668
rect 163924 199656 163930 199708
rect 164252 199640 164280 199736
rect 164326 199724 164332 199776
rect 164384 199724 164390 199776
rect 164482 199640 164510 200008
rect 164850 200008 165614 200036
rect 164556 199860 164562 199912
rect 164614 199860 164620 199912
rect 164574 199832 164602 199860
rect 164850 199844 164878 200008
rect 164574 199804 164786 199832
rect 164234 199588 164240 199640
rect 164292 199588 164298 199640
rect 164418 199588 164424 199640
rect 164476 199600 164510 199640
rect 164476 199588 164482 199600
rect 163682 199520 163688 199572
rect 163740 199520 163746 199572
rect 163958 199520 163964 199572
rect 164016 199560 164022 199572
rect 164602 199560 164608 199572
rect 164016 199532 164608 199560
rect 164016 199520 164022 199532
rect 164602 199520 164608 199532
rect 164660 199520 164666 199572
rect 164758 199504 164786 199804
rect 164832 199792 164838 199844
rect 164890 199792 164896 199844
rect 164924 199792 164930 199844
rect 164982 199792 164988 199844
rect 165016 199792 165022 199844
rect 165074 199792 165080 199844
rect 165292 199792 165298 199844
rect 165350 199792 165356 199844
rect 164942 199504 164970 199792
rect 165034 199628 165062 199792
rect 165154 199628 165160 199640
rect 165034 199600 165160 199628
rect 165154 199588 165160 199600
rect 165212 199588 165218 199640
rect 165310 199504 165338 199792
rect 165586 199640 165614 200008
rect 165660 199724 165666 199776
rect 165718 199724 165724 199776
rect 165678 199696 165706 199724
rect 165678 199668 165936 199696
rect 165586 199600 165620 199640
rect 165614 199588 165620 199600
rect 165672 199588 165678 199640
rect 165706 199520 165712 199572
rect 165764 199560 165770 199572
rect 165908 199560 165936 199668
rect 165764 199532 165936 199560
rect 165764 199520 165770 199532
rect 164510 199492 164516 199504
rect 163700 199464 164516 199492
rect 163590 199384 163596 199436
rect 163648 199424 163654 199436
rect 163700 199424 163728 199464
rect 164510 199452 164516 199464
rect 164568 199452 164574 199504
rect 164758 199464 164792 199504
rect 164786 199452 164792 199464
rect 164844 199452 164850 199504
rect 164942 199464 164976 199504
rect 164970 199452 164976 199464
rect 165028 199452 165034 199504
rect 165310 199464 165344 199504
rect 165338 199452 165344 199464
rect 165396 199452 165402 199504
rect 166000 199492 166028 200076
rect 166396 199900 166402 199912
rect 166368 199860 166402 199900
rect 166454 199860 166460 199912
rect 166488 199860 166494 199912
rect 166546 199860 166552 199912
rect 166580 199860 166586 199912
rect 166638 199860 166644 199912
rect 166672 199860 166678 199912
rect 166730 199860 166736 199912
rect 166764 199860 166770 199912
rect 166822 199860 166828 199912
rect 166368 199776 166396 199860
rect 166506 199832 166534 199860
rect 166460 199804 166534 199832
rect 166350 199724 166356 199776
rect 166408 199724 166414 199776
rect 166460 199708 166488 199804
rect 166598 199776 166626 199860
rect 166534 199724 166540 199776
rect 166592 199736 166626 199776
rect 166592 199724 166598 199736
rect 166690 199708 166718 199860
rect 166442 199656 166448 199708
rect 166500 199656 166506 199708
rect 166626 199656 166632 199708
rect 166684 199668 166718 199708
rect 166684 199656 166690 199668
rect 166782 199572 166810 199860
rect 166920 199640 166948 200144
rect 167040 199860 167046 199912
rect 167098 199860 167104 199912
rect 167500 199860 167506 199912
rect 167558 199860 167564 199912
rect 167592 199860 167598 199912
rect 167650 199860 167656 199912
rect 166902 199588 166908 199640
rect 166960 199588 166966 199640
rect 166718 199520 166724 199572
rect 166776 199532 166810 199572
rect 167058 199560 167086 199860
rect 167316 199832 167322 199844
rect 167288 199792 167322 199832
rect 167374 199792 167380 199844
rect 167288 199640 167316 199792
rect 167518 199764 167546 199860
rect 167472 199736 167546 199764
rect 167270 199588 167276 199640
rect 167328 199588 167334 199640
rect 167362 199560 167368 199572
rect 167058 199532 167368 199560
rect 166776 199520 166782 199532
rect 167362 199520 167368 199532
rect 167420 199520 167426 199572
rect 166258 199492 166264 199504
rect 166000 199464 166264 199492
rect 166258 199452 166264 199464
rect 166316 199452 166322 199504
rect 167472 199492 167500 199736
rect 167610 199708 167638 199860
rect 167546 199656 167552 199708
rect 167604 199668 167638 199708
rect 167604 199656 167610 199668
rect 167776 199656 167782 199708
rect 167834 199656 167840 199708
rect 167794 199572 167822 199656
rect 167730 199520 167736 199572
rect 167788 199532 167822 199572
rect 168024 199560 168052 200212
rect 168144 199860 168150 199912
rect 168202 199860 168208 199912
rect 168236 199860 168242 199912
rect 168294 199900 168300 199912
rect 168294 199860 168328 199900
rect 168162 199708 168190 199860
rect 168162 199668 168196 199708
rect 168190 199656 168196 199668
rect 168248 199656 168254 199708
rect 168098 199588 168104 199640
rect 168156 199628 168162 199640
rect 168300 199628 168328 199860
rect 168512 199724 168518 199776
rect 168570 199724 168576 199776
rect 168420 199656 168426 199708
rect 168478 199656 168484 199708
rect 168156 199600 168328 199628
rect 168156 199588 168162 199600
rect 168438 199572 168466 199656
rect 168530 199640 168558 199724
rect 168668 199640 168696 200280
rect 168788 199860 168794 199912
rect 168846 199860 168852 199912
rect 168880 199860 168886 199912
rect 168938 199860 168944 199912
rect 168806 199708 168834 199860
rect 168898 199776 168926 199860
rect 169064 199792 169070 199844
rect 169122 199792 169128 199844
rect 168898 199736 168932 199776
rect 168926 199724 168932 199736
rect 168984 199724 168990 199776
rect 169082 199708 169110 199792
rect 168806 199668 168840 199708
rect 168834 199656 168840 199668
rect 168892 199656 168898 199708
rect 169018 199656 169024 199708
rect 169076 199668 169110 199708
rect 169076 199656 169082 199668
rect 169174 199640 169202 200280
rect 170232 200104 170260 200620
rect 172394 200580 172422 200620
rect 172486 200620 172606 200648
rect 172486 200580 172514 200620
rect 172394 200552 172514 200580
rect 170140 200076 170260 200104
rect 170554 200484 171778 200512
rect 170140 199968 170168 200076
rect 170554 199968 170582 200484
rect 171750 200308 171778 200484
rect 173682 200444 173710 200688
rect 177758 200676 177764 200728
rect 177816 200676 177822 200728
rect 178862 200676 178868 200728
rect 178920 200716 178926 200728
rect 179386 200716 179414 200756
rect 179984 200728 180012 200756
rect 178920 200688 179414 200716
rect 178920 200676 178926 200688
rect 179966 200676 179972 200728
rect 180024 200676 180030 200728
rect 178678 200608 178684 200660
rect 178736 200648 178742 200660
rect 180076 200648 180104 200892
rect 189074 200784 189080 200796
rect 180260 200756 189080 200784
rect 180260 200728 180288 200756
rect 189074 200744 189080 200756
rect 189132 200744 189138 200796
rect 180242 200676 180248 200728
rect 180300 200676 180306 200728
rect 178736 200620 180104 200648
rect 178736 200608 178742 200620
rect 177850 200540 177856 200592
rect 177908 200580 177914 200592
rect 178770 200580 178776 200592
rect 177908 200552 178776 200580
rect 177908 200540 177914 200552
rect 178770 200540 178776 200552
rect 178828 200540 178834 200592
rect 199010 200444 199016 200456
rect 173682 200416 199016 200444
rect 199010 200404 199016 200416
rect 199068 200404 199074 200456
rect 177758 200336 177764 200388
rect 177816 200376 177822 200388
rect 193306 200376 193312 200388
rect 177816 200348 193312 200376
rect 177816 200336 177822 200348
rect 193306 200336 193312 200348
rect 193364 200336 193370 200388
rect 187694 200308 187700 200320
rect 171750 200280 187700 200308
rect 187694 200268 187700 200280
rect 187752 200268 187758 200320
rect 186682 200240 186688 200252
rect 171612 200212 186688 200240
rect 171612 199968 171640 200212
rect 186682 200200 186688 200212
rect 186740 200200 186746 200252
rect 213914 200172 213920 200184
rect 170140 199940 170306 199968
rect 169248 199792 169254 199844
rect 169306 199792 169312 199844
rect 169432 199792 169438 199844
rect 169490 199792 169496 199844
rect 169524 199792 169530 199844
rect 169582 199792 169588 199844
rect 170168 199832 170174 199844
rect 169680 199804 170174 199832
rect 168530 199600 168564 199640
rect 168558 199588 168564 199600
rect 168616 199588 168622 199640
rect 168650 199588 168656 199640
rect 168708 199588 168714 199640
rect 169110 199588 169116 199640
rect 169168 199600 169202 199640
rect 169168 199588 169174 199600
rect 168282 199560 168288 199572
rect 168024 199532 168288 199560
rect 167788 199520 167794 199532
rect 168282 199520 168288 199532
rect 168340 199520 168346 199572
rect 168374 199520 168380 199572
rect 168432 199532 168466 199572
rect 168432 199520 168438 199532
rect 168466 199492 168472 199504
rect 167472 199464 168472 199492
rect 168466 199452 168472 199464
rect 168524 199452 168530 199504
rect 169110 199452 169116 199504
rect 169168 199492 169174 199504
rect 169266 199492 169294 199792
rect 169450 199696 169478 199792
rect 169404 199668 169478 199696
rect 169404 199640 169432 199668
rect 169542 199640 169570 199792
rect 169386 199588 169392 199640
rect 169444 199588 169450 199640
rect 169478 199588 169484 199640
rect 169536 199600 169570 199640
rect 169536 199588 169542 199600
rect 169570 199520 169576 199572
rect 169628 199560 169634 199572
rect 169680 199560 169708 199804
rect 170168 199792 170174 199804
rect 170226 199792 170232 199844
rect 170278 199708 170306 199940
rect 170214 199656 170220 199708
rect 170272 199668 170306 199708
rect 170370 199940 170582 199968
rect 171244 199940 171640 199968
rect 172486 200144 213920 200172
rect 170272 199656 170278 199668
rect 170370 199628 170398 199940
rect 170996 199900 171002 199912
rect 170554 199872 171002 199900
rect 170444 199792 170450 199844
rect 170502 199792 170508 199844
rect 169628 199532 169708 199560
rect 169956 199600 170398 199628
rect 169628 199520 169634 199532
rect 169956 199504 169984 199600
rect 170462 199572 170490 199792
rect 170398 199520 170404 199572
rect 170456 199532 170490 199572
rect 170456 199520 170462 199532
rect 170554 199504 170582 199872
rect 170996 199860 171002 199872
rect 171054 199860 171060 199912
rect 171088 199860 171094 199912
rect 171146 199900 171152 199912
rect 171146 199860 171180 199900
rect 170812 199792 170818 199844
rect 170870 199792 170876 199844
rect 170720 199764 170726 199776
rect 170646 199736 170726 199764
rect 170646 199560 170674 199736
rect 170720 199724 170726 199736
rect 170778 199724 170784 199776
rect 170830 199696 170858 199792
rect 171042 199696 171048 199708
rect 170830 199668 171048 199696
rect 171042 199656 171048 199668
rect 171100 199656 171106 199708
rect 171152 199640 171180 199860
rect 171244 199640 171272 199940
rect 171456 199860 171462 199912
rect 171514 199860 171520 199912
rect 171548 199860 171554 199912
rect 171606 199860 171612 199912
rect 172008 199900 172014 199912
rect 171888 199872 172014 199900
rect 171134 199588 171140 199640
rect 171192 199588 171198 199640
rect 171226 199588 171232 199640
rect 171284 199588 171290 199640
rect 170766 199560 170772 199572
rect 170646 199532 170772 199560
rect 170766 199520 170772 199532
rect 170824 199520 170830 199572
rect 169168 199464 169294 199492
rect 169168 199452 169174 199464
rect 169938 199452 169944 199504
rect 169996 199452 170002 199504
rect 170490 199452 170496 199504
rect 170548 199464 170582 199504
rect 171474 199504 171502 199860
rect 171566 199560 171594 199860
rect 171732 199792 171738 199844
rect 171790 199792 171796 199844
rect 171750 199640 171778 199792
rect 171888 199640 171916 199872
rect 172008 199860 172014 199872
rect 172066 199860 172072 199912
rect 172376 199900 172382 199912
rect 172118 199872 172382 199900
rect 172118 199640 172146 199872
rect 172376 199860 172382 199872
rect 172434 199860 172440 199912
rect 172486 199832 172514 200144
rect 213914 200132 213920 200144
rect 213972 200132 213978 200184
rect 173222 200076 186314 200104
rect 172836 199900 172842 199912
rect 172256 199804 172514 199832
rect 172624 199872 172842 199900
rect 172256 199640 172284 199804
rect 172376 199764 172382 199776
rect 172348 199724 172382 199764
rect 172434 199724 172440 199776
rect 171686 199588 171692 199640
rect 171744 199600 171778 199640
rect 171744 199588 171750 199600
rect 171870 199588 171876 199640
rect 171928 199588 171934 199640
rect 172118 199600 172152 199640
rect 172146 199588 172152 199600
rect 172204 199588 172210 199640
rect 172238 199588 172244 199640
rect 172296 199588 172302 199640
rect 172348 199572 172376 199724
rect 172054 199560 172060 199572
rect 171566 199532 172060 199560
rect 172054 199520 172060 199532
rect 172112 199520 172118 199572
rect 172330 199520 172336 199572
rect 172388 199520 172394 199572
rect 171474 199464 171508 199504
rect 170548 199452 170554 199464
rect 171502 199452 171508 199464
rect 171560 199452 171566 199504
rect 172422 199452 172428 199504
rect 172480 199492 172486 199504
rect 172624 199492 172652 199872
rect 172836 199860 172842 199872
rect 172894 199860 172900 199912
rect 172946 199872 173158 199900
rect 172946 199832 172974 199872
rect 172716 199804 172974 199832
rect 172716 199504 172744 199804
rect 173020 199792 173026 199844
rect 173078 199792 173084 199844
rect 173038 199628 173066 199792
rect 173130 199696 173158 199872
rect 173222 199776 173250 200076
rect 178034 200036 178040 200048
rect 173682 200008 178040 200036
rect 173682 199900 173710 200008
rect 178034 199996 178040 200008
rect 178092 199996 178098 200048
rect 181990 199968 181996 199980
rect 173774 199940 174078 199968
rect 173774 199912 173802 199940
rect 173636 199872 173710 199900
rect 173204 199724 173210 199776
rect 173262 199724 173268 199776
rect 173636 199696 173664 199872
rect 173756 199860 173762 199912
rect 173814 199860 173820 199912
rect 173848 199860 173854 199912
rect 173906 199860 173912 199912
rect 173940 199860 173946 199912
rect 173998 199860 174004 199912
rect 173866 199832 173894 199860
rect 173130 199668 173664 199696
rect 173728 199804 173894 199832
rect 172992 199600 173066 199628
rect 172992 199504 173020 199600
rect 173728 199560 173756 199804
rect 173958 199776 173986 199860
rect 173802 199724 173808 199776
rect 173860 199724 173866 199776
rect 173894 199724 173900 199776
rect 173952 199736 173986 199776
rect 173952 199724 173958 199736
rect 173820 199696 173848 199724
rect 174050 199696 174078 199940
rect 174280 199940 174814 199968
rect 174124 199860 174130 199912
rect 174182 199860 174188 199912
rect 173820 199668 174078 199696
rect 174142 199628 174170 199860
rect 174280 199640 174308 199940
rect 174786 199912 174814 199940
rect 175522 199940 181996 199968
rect 175522 199912 175550 199940
rect 181990 199928 181996 199940
rect 182048 199928 182054 199980
rect 174492 199860 174498 199912
rect 174550 199860 174556 199912
rect 174768 199860 174774 199912
rect 174826 199860 174832 199912
rect 174860 199860 174866 199912
rect 174918 199860 174924 199912
rect 174952 199860 174958 199912
rect 175010 199860 175016 199912
rect 175320 199900 175326 199912
rect 175246 199872 175326 199900
rect 174510 199776 174538 199860
rect 174676 199832 174682 199844
rect 174446 199724 174452 199776
rect 174504 199736 174538 199776
rect 174602 199804 174682 199832
rect 174504 199724 174510 199736
rect 174602 199708 174630 199804
rect 174676 199792 174682 199804
rect 174734 199792 174740 199844
rect 174878 199832 174906 199860
rect 174832 199804 174906 199832
rect 174538 199656 174544 199708
rect 174596 199668 174630 199708
rect 174596 199656 174602 199668
rect 173912 199600 174170 199628
rect 173802 199560 173808 199572
rect 173728 199532 173808 199560
rect 173802 199520 173808 199532
rect 173860 199520 173866 199572
rect 172480 199464 172652 199492
rect 172480 199452 172486 199464
rect 172698 199452 172704 199504
rect 172756 199452 172762 199504
rect 172974 199452 172980 199504
rect 173032 199452 173038 199504
rect 173912 199492 173940 199600
rect 174262 199588 174268 199640
rect 174320 199588 174326 199640
rect 173986 199520 173992 199572
rect 174044 199560 174050 199572
rect 174538 199560 174544 199572
rect 174044 199532 174544 199560
rect 174044 199520 174050 199532
rect 174538 199520 174544 199532
rect 174596 199520 174602 199572
rect 174832 199504 174860 199804
rect 174970 199708 174998 199860
rect 174906 199656 174912 199708
rect 174964 199668 174998 199708
rect 174964 199656 174970 199668
rect 175246 199504 175274 199872
rect 175320 199860 175326 199872
rect 175378 199860 175384 199912
rect 175504 199860 175510 199912
rect 175562 199860 175568 199912
rect 175964 199900 175970 199912
rect 175660 199872 175970 199900
rect 175412 199792 175418 199844
rect 175470 199792 175476 199844
rect 175430 199640 175458 199792
rect 175366 199588 175372 199640
rect 175424 199600 175458 199640
rect 175424 199588 175430 199600
rect 175660 199504 175688 199872
rect 175964 199860 175970 199872
rect 176022 199860 176028 199912
rect 176056 199860 176062 199912
rect 176114 199860 176120 199912
rect 176792 199860 176798 199912
rect 176850 199860 176856 199912
rect 176884 199860 176890 199912
rect 176942 199900 176948 199912
rect 178862 199900 178868 199912
rect 176942 199872 178868 199900
rect 176942 199860 176948 199872
rect 178862 199860 178868 199872
rect 178920 199860 178926 199912
rect 176074 199776 176102 199860
rect 176010 199724 176016 199776
rect 176068 199736 176102 199776
rect 176810 199776 176838 199860
rect 177666 199792 177672 199844
rect 177724 199832 177730 199844
rect 180150 199832 180156 199844
rect 177724 199804 180156 199832
rect 177724 199792 177730 199804
rect 180150 199792 180156 199804
rect 180208 199792 180214 199844
rect 176810 199736 176844 199776
rect 176068 199724 176074 199736
rect 176838 199724 176844 199736
rect 176896 199724 176902 199776
rect 180334 199764 180340 199776
rect 177684 199736 180340 199764
rect 177684 199696 177712 199736
rect 180334 199724 180340 199736
rect 180392 199724 180398 199776
rect 186286 199764 186314 200076
rect 187878 199764 187884 199776
rect 186286 199736 187884 199764
rect 187878 199724 187884 199736
rect 187936 199724 187942 199776
rect 214006 199696 214012 199708
rect 175936 199668 177712 199696
rect 177776 199668 214012 199696
rect 175936 199640 175964 199668
rect 175918 199588 175924 199640
rect 175976 199588 175982 199640
rect 176746 199588 176752 199640
rect 176804 199628 176810 199640
rect 177666 199628 177672 199640
rect 176804 199600 177672 199628
rect 176804 199588 176810 199600
rect 177666 199588 177672 199600
rect 177724 199588 177730 199640
rect 177776 199560 177804 199668
rect 214006 199656 214012 199668
rect 214064 199656 214070 199708
rect 177942 199588 177948 199640
rect 178000 199628 178006 199640
rect 215846 199628 215852 199640
rect 178000 199600 215852 199628
rect 178000 199588 178006 199600
rect 215846 199588 215852 199600
rect 215904 199588 215910 199640
rect 175798 199532 177804 199560
rect 174170 199492 174176 199504
rect 173912 199464 174176 199492
rect 174170 199452 174176 199464
rect 174228 199452 174234 199504
rect 174262 199452 174268 199504
rect 174320 199492 174326 199504
rect 174722 199492 174728 199504
rect 174320 199464 174728 199492
rect 174320 199452 174326 199464
rect 174722 199452 174728 199464
rect 174780 199452 174786 199504
rect 174814 199452 174820 199504
rect 174872 199452 174878 199504
rect 175182 199452 175188 199504
rect 175240 199464 175274 199504
rect 175240 199452 175246 199464
rect 175642 199452 175648 199504
rect 175700 199452 175706 199504
rect 163648 199396 163728 199424
rect 163648 199384 163654 199396
rect 163958 199384 163964 199436
rect 164016 199424 164022 199436
rect 169202 199424 169208 199436
rect 164016 199396 169208 199424
rect 164016 199384 164022 199396
rect 169202 199384 169208 199396
rect 169260 199384 169266 199436
rect 169754 199384 169760 199436
rect 169812 199424 169818 199436
rect 175798 199424 175826 199532
rect 175918 199452 175924 199504
rect 175976 199492 175982 199504
rect 180150 199492 180156 199504
rect 175976 199464 180156 199492
rect 175976 199452 175982 199464
rect 180150 199452 180156 199464
rect 180208 199452 180214 199504
rect 182910 199452 182916 199504
rect 182968 199492 182974 199504
rect 190454 199492 190460 199504
rect 182968 199464 190460 199492
rect 182968 199452 182974 199464
rect 190454 199452 190460 199464
rect 190512 199452 190518 199504
rect 169812 199396 175826 199424
rect 169812 199384 169818 199396
rect 181070 199384 181076 199436
rect 181128 199424 181134 199436
rect 190546 199424 190552 199436
rect 181128 199396 190552 199424
rect 181128 199384 181134 199396
rect 190546 199384 190552 199396
rect 190604 199384 190610 199436
rect 215570 199356 215576 199368
rect 159376 199260 163544 199288
rect 163608 199328 215576 199356
rect 157242 199180 157248 199232
rect 157300 199220 157306 199232
rect 161658 199220 161664 199232
rect 157300 199192 161664 199220
rect 157300 199180 157306 199192
rect 161658 199180 161664 199192
rect 161716 199180 161722 199232
rect 163608 199152 163636 199328
rect 215570 199316 215576 199328
rect 215628 199316 215634 199368
rect 163682 199248 163688 199300
rect 163740 199288 163746 199300
rect 193214 199288 193220 199300
rect 163740 199260 193220 199288
rect 163740 199248 163746 199260
rect 193214 199248 193220 199260
rect 193272 199248 193278 199300
rect 189994 199220 190000 199232
rect 154546 199124 163636 199152
rect 163700 199192 190000 199220
rect 108574 199044 108580 199096
rect 108632 199084 108638 199096
rect 131574 199084 131580 199096
rect 108632 199056 131580 199084
rect 108632 199044 108638 199056
rect 131574 199044 131580 199056
rect 131632 199044 131638 199096
rect 133506 199084 133512 199096
rect 132696 199056 133512 199084
rect 115842 198976 115848 199028
rect 115900 199016 115906 199028
rect 131758 199016 131764 199028
rect 115900 198988 131764 199016
rect 115900 198976 115906 198988
rect 131758 198976 131764 198988
rect 131816 198976 131822 199028
rect 132034 198976 132040 199028
rect 132092 199016 132098 199028
rect 132696 199016 132724 199056
rect 133506 199044 133512 199056
rect 133564 199044 133570 199096
rect 135070 199044 135076 199096
rect 135128 199084 135134 199096
rect 135714 199084 135720 199096
rect 135128 199056 135720 199084
rect 135128 199044 135134 199056
rect 135714 199044 135720 199056
rect 135772 199044 135778 199096
rect 135898 199044 135904 199096
rect 135956 199084 135962 199096
rect 144822 199084 144828 199096
rect 135956 199056 144828 199084
rect 135956 199044 135962 199056
rect 144822 199044 144828 199056
rect 144880 199044 144886 199096
rect 154574 199044 154580 199096
rect 154632 199084 154638 199096
rect 156414 199084 156420 199096
rect 154632 199056 156420 199084
rect 154632 199044 154638 199056
rect 156414 199044 156420 199056
rect 156472 199044 156478 199096
rect 156690 199044 156696 199096
rect 156748 199084 156754 199096
rect 156748 199056 160508 199084
rect 156748 199044 156754 199056
rect 132092 198988 132264 199016
rect 132092 198976 132098 198988
rect 130010 198908 130016 198960
rect 130068 198948 130074 198960
rect 132126 198948 132132 198960
rect 130068 198920 132132 198948
rect 130068 198908 130074 198920
rect 132126 198908 132132 198920
rect 132184 198908 132190 198960
rect 132236 198948 132264 198988
rect 132512 198988 132724 199016
rect 132512 198948 132540 198988
rect 138290 198976 138296 199028
rect 138348 199016 138354 199028
rect 147674 199016 147680 199028
rect 138348 198988 147680 199016
rect 138348 198976 138354 198988
rect 147674 198976 147680 198988
rect 147732 198976 147738 199028
rect 150710 198976 150716 199028
rect 150768 199016 150774 199028
rect 157794 199016 157800 199028
rect 150768 198988 157800 199016
rect 150768 198976 150774 198988
rect 157794 198976 157800 198988
rect 157852 198976 157858 199028
rect 160480 199016 160508 199056
rect 161658 199044 161664 199096
rect 161716 199084 161722 199096
rect 163700 199084 163728 199192
rect 189994 199180 190000 199192
rect 190052 199180 190058 199232
rect 163958 199112 163964 199164
rect 164016 199152 164022 199164
rect 189258 199152 189264 199164
rect 164016 199124 189264 199152
rect 164016 199112 164022 199124
rect 189258 199112 189264 199124
rect 189316 199112 189322 199164
rect 190546 199084 190552 199096
rect 161716 199056 163728 199084
rect 164390 199056 190552 199084
rect 161716 199044 161722 199056
rect 160480 198988 164234 199016
rect 132236 198920 132540 198948
rect 132862 198908 132868 198960
rect 132920 198948 132926 198960
rect 135898 198948 135904 198960
rect 132920 198920 135904 198948
rect 132920 198908 132926 198920
rect 135898 198908 135904 198920
rect 135956 198908 135962 198960
rect 137002 198908 137008 198960
rect 137060 198948 137066 198960
rect 139394 198948 139400 198960
rect 137060 198920 139400 198948
rect 137060 198908 137066 198920
rect 139394 198908 139400 198920
rect 139452 198908 139458 198960
rect 141418 198908 141424 198960
rect 141476 198948 141482 198960
rect 141476 198920 142568 198948
rect 141476 198908 141482 198920
rect 121270 198840 121276 198892
rect 121328 198880 121334 198892
rect 142154 198880 142160 198892
rect 121328 198852 142160 198880
rect 121328 198840 121334 198852
rect 142154 198840 142160 198852
rect 142212 198840 142218 198892
rect 142540 198880 142568 198920
rect 142614 198908 142620 198960
rect 142672 198948 142678 198960
rect 142982 198948 142988 198960
rect 142672 198920 142988 198948
rect 142672 198908 142678 198920
rect 142982 198908 142988 198920
rect 143040 198908 143046 198960
rect 143902 198908 143908 198960
rect 143960 198948 143966 198960
rect 146294 198948 146300 198960
rect 143960 198920 146300 198948
rect 143960 198908 143966 198920
rect 146294 198908 146300 198920
rect 146352 198908 146358 198960
rect 152274 198908 152280 198960
rect 152332 198948 152338 198960
rect 152332 198920 160094 198948
rect 152332 198908 152338 198920
rect 143166 198880 143172 198892
rect 142540 198852 143172 198880
rect 143166 198840 143172 198852
rect 143224 198840 143230 198892
rect 160066 198880 160094 198920
rect 160186 198908 160192 198960
rect 160244 198948 160250 198960
rect 163222 198948 163228 198960
rect 160244 198920 163228 198948
rect 160244 198908 160250 198920
rect 163222 198908 163228 198920
rect 163280 198908 163286 198960
rect 164206 198948 164234 198988
rect 164206 198920 164326 198948
rect 164298 198880 164326 198920
rect 164390 198880 164418 199056
rect 190546 199044 190552 199056
rect 190604 199044 190610 199096
rect 165338 198976 165344 199028
rect 165396 199016 165402 199028
rect 168466 199016 168472 199028
rect 165396 198988 168472 199016
rect 165396 198976 165402 198988
rect 168466 198976 168472 198988
rect 168524 198976 168530 199028
rect 168650 198976 168656 199028
rect 168708 199016 168714 199028
rect 200298 199016 200304 199028
rect 168708 198988 200304 199016
rect 168708 198976 168714 198988
rect 200298 198976 200304 198988
rect 200356 198976 200362 199028
rect 168282 198908 168288 198960
rect 168340 198948 168346 198960
rect 171226 198948 171232 198960
rect 168340 198920 171232 198948
rect 168340 198908 168346 198920
rect 171226 198908 171232 198920
rect 171284 198908 171290 198960
rect 172054 198908 172060 198960
rect 172112 198948 172118 198960
rect 172698 198948 172704 198960
rect 172112 198920 172704 198948
rect 172112 198908 172118 198920
rect 172698 198908 172704 198920
rect 172756 198908 172762 198960
rect 174262 198908 174268 198960
rect 174320 198948 174326 198960
rect 178862 198948 178868 198960
rect 174320 198920 178868 198948
rect 174320 198908 174326 198920
rect 178862 198908 178868 198920
rect 178920 198908 178926 198960
rect 186590 198948 186596 198960
rect 186286 198920 186596 198948
rect 186286 198880 186314 198920
rect 186590 198908 186596 198920
rect 186648 198908 186654 198960
rect 160066 198852 164234 198880
rect 164298 198852 164418 198880
rect 166828 198852 186314 198880
rect 126330 198772 126336 198824
rect 126388 198812 126394 198824
rect 147858 198812 147864 198824
rect 126388 198784 147864 198812
rect 126388 198772 126394 198784
rect 147858 198772 147864 198784
rect 147916 198772 147922 198824
rect 154758 198772 154764 198824
rect 154816 198812 154822 198824
rect 163958 198812 163964 198824
rect 154816 198784 163964 198812
rect 154816 198772 154822 198784
rect 163958 198772 163964 198784
rect 164016 198772 164022 198824
rect 164206 198812 164234 198852
rect 166828 198812 166856 198852
rect 164206 198784 166856 198812
rect 168466 198772 168472 198824
rect 168524 198812 168530 198824
rect 182818 198812 182824 198824
rect 168524 198784 182824 198812
rect 168524 198772 168530 198784
rect 182818 198772 182824 198784
rect 182876 198772 182882 198824
rect 126422 198704 126428 198756
rect 126480 198744 126486 198756
rect 149054 198744 149060 198756
rect 126480 198716 149060 198744
rect 126480 198704 126486 198716
rect 149054 198704 149060 198716
rect 149112 198704 149118 198756
rect 157334 198704 157340 198756
rect 157392 198744 157398 198756
rect 180058 198744 180064 198756
rect 157392 198716 180064 198744
rect 157392 198704 157398 198716
rect 180058 198704 180064 198716
rect 180116 198704 180122 198756
rect 184290 198704 184296 198756
rect 184348 198744 184354 198756
rect 189166 198744 189172 198756
rect 184348 198716 189172 198744
rect 184348 198704 184354 198716
rect 189166 198704 189172 198716
rect 189224 198704 189230 198756
rect 129274 198636 129280 198688
rect 129332 198676 129338 198688
rect 144086 198676 144092 198688
rect 129332 198648 144092 198676
rect 129332 198636 129338 198648
rect 144086 198636 144092 198648
rect 144144 198636 144150 198688
rect 154850 198636 154856 198688
rect 154908 198676 154914 198688
rect 162486 198676 162492 198688
rect 154908 198648 162492 198676
rect 154908 198636 154914 198648
rect 162486 198636 162492 198648
rect 162544 198636 162550 198688
rect 164510 198636 164516 198688
rect 164568 198676 164574 198688
rect 170674 198676 170680 198688
rect 164568 198648 170680 198676
rect 164568 198636 164574 198648
rect 170674 198636 170680 198648
rect 170732 198636 170738 198688
rect 170858 198636 170864 198688
rect 170916 198676 170922 198688
rect 177850 198676 177856 198688
rect 170916 198648 177856 198676
rect 170916 198636 170922 198648
rect 177850 198636 177856 198648
rect 177908 198636 177914 198688
rect 128998 198568 129004 198620
rect 129056 198608 129062 198620
rect 149330 198608 149336 198620
rect 129056 198580 149336 198608
rect 129056 198568 129062 198580
rect 149330 198568 149336 198580
rect 149388 198568 149394 198620
rect 157702 198568 157708 198620
rect 157760 198608 157766 198620
rect 157760 198580 165568 198608
rect 157760 198568 157766 198580
rect 165540 198552 165568 198580
rect 167086 198568 167092 198620
rect 167144 198608 167150 198620
rect 170214 198608 170220 198620
rect 167144 198580 170220 198608
rect 167144 198568 167150 198580
rect 170214 198568 170220 198580
rect 170272 198568 170278 198620
rect 172606 198568 172612 198620
rect 172664 198608 172670 198620
rect 211338 198608 211344 198620
rect 172664 198580 211344 198608
rect 172664 198568 172670 198580
rect 211338 198568 211344 198580
rect 211396 198568 211402 198620
rect 126514 198500 126520 198552
rect 126572 198540 126578 198552
rect 147766 198540 147772 198552
rect 126572 198512 147772 198540
rect 126572 198500 126578 198512
rect 147766 198500 147772 198512
rect 147824 198500 147830 198552
rect 165522 198500 165528 198552
rect 165580 198500 165586 198552
rect 172974 198500 172980 198552
rect 173032 198540 173038 198552
rect 211522 198540 211528 198552
rect 173032 198512 211528 198540
rect 173032 198500 173038 198512
rect 211522 198500 211528 198512
rect 211580 198500 211586 198552
rect 122374 198432 122380 198484
rect 122432 198472 122438 198484
rect 147122 198472 147128 198484
rect 122432 198444 147128 198472
rect 122432 198432 122438 198444
rect 147122 198432 147128 198444
rect 147180 198432 147186 198484
rect 159542 198432 159548 198484
rect 159600 198472 159606 198484
rect 166258 198472 166264 198484
rect 159600 198444 166264 198472
rect 159600 198432 159606 198444
rect 166258 198432 166264 198444
rect 166316 198432 166322 198484
rect 168834 198432 168840 198484
rect 168892 198472 168898 198484
rect 170858 198472 170864 198484
rect 168892 198444 170864 198472
rect 168892 198432 168898 198444
rect 170858 198432 170864 198444
rect 170916 198432 170922 198484
rect 170950 198432 170956 198484
rect 171008 198472 171014 198484
rect 208854 198472 208860 198484
rect 171008 198444 208860 198472
rect 171008 198432 171014 198444
rect 208854 198432 208860 198444
rect 208912 198432 208918 198484
rect 125042 198364 125048 198416
rect 125100 198404 125106 198416
rect 149422 198404 149428 198416
rect 125100 198376 149428 198404
rect 125100 198364 125106 198376
rect 149422 198364 149428 198376
rect 149480 198364 149486 198416
rect 159726 198364 159732 198416
rect 159784 198404 159790 198416
rect 172054 198404 172060 198416
rect 159784 198376 172060 198404
rect 159784 198364 159790 198376
rect 172054 198364 172060 198376
rect 172112 198364 172118 198416
rect 173802 198364 173808 198416
rect 173860 198404 173866 198416
rect 212718 198404 212724 198416
rect 173860 198376 212724 198404
rect 173860 198364 173866 198376
rect 212718 198364 212724 198376
rect 212776 198364 212782 198416
rect 122282 198296 122288 198348
rect 122340 198336 122346 198348
rect 146846 198336 146852 198348
rect 122340 198308 146852 198336
rect 122340 198296 122346 198308
rect 146846 198296 146852 198308
rect 146904 198296 146910 198348
rect 165706 198336 165712 198348
rect 157306 198308 165712 198336
rect 105722 198228 105728 198280
rect 105780 198268 105786 198280
rect 127526 198268 127532 198280
rect 105780 198240 127532 198268
rect 105780 198228 105786 198240
rect 127526 198228 127532 198240
rect 127584 198228 127590 198280
rect 107010 198160 107016 198212
rect 107068 198200 107074 198212
rect 135990 198200 135996 198212
rect 107068 198172 135996 198200
rect 107068 198160 107074 198172
rect 135990 198160 135996 198172
rect 136048 198160 136054 198212
rect 141050 198160 141056 198212
rect 141108 198200 141114 198212
rect 141510 198200 141516 198212
rect 141108 198172 141516 198200
rect 141108 198160 141114 198172
rect 141510 198160 141516 198172
rect 141568 198160 141574 198212
rect 151722 198160 151728 198212
rect 151780 198200 151786 198212
rect 157306 198200 157334 198308
rect 165706 198296 165712 198308
rect 165764 198296 165770 198348
rect 167086 198296 167092 198348
rect 167144 198336 167150 198348
rect 168098 198336 168104 198348
rect 167144 198308 168104 198336
rect 167144 198296 167150 198308
rect 168098 198296 168104 198308
rect 168156 198296 168162 198348
rect 171134 198296 171140 198348
rect 171192 198336 171198 198348
rect 172606 198336 172612 198348
rect 171192 198308 172612 198336
rect 171192 198296 171198 198308
rect 172606 198296 172612 198308
rect 172664 198296 172670 198348
rect 173618 198296 173624 198348
rect 173676 198336 173682 198348
rect 212902 198336 212908 198348
rect 173676 198308 212908 198336
rect 173676 198296 173682 198308
rect 212902 198296 212908 198308
rect 212960 198296 212966 198348
rect 163038 198228 163044 198280
rect 163096 198268 163102 198280
rect 168834 198268 168840 198280
rect 163096 198240 168840 198268
rect 163096 198228 163102 198240
rect 168834 198228 168840 198240
rect 168892 198228 168898 198280
rect 170490 198228 170496 198280
rect 170548 198268 170554 198280
rect 170950 198268 170956 198280
rect 170548 198240 170956 198268
rect 170548 198228 170554 198240
rect 170950 198228 170956 198240
rect 171008 198228 171014 198280
rect 172514 198228 172520 198280
rect 172572 198268 172578 198280
rect 212626 198268 212632 198280
rect 172572 198240 212632 198268
rect 172572 198228 172578 198240
rect 212626 198228 212632 198240
rect 212684 198228 212690 198280
rect 151780 198172 157334 198200
rect 151780 198160 151786 198172
rect 159818 198160 159824 198212
rect 159876 198200 159882 198212
rect 171134 198200 171140 198212
rect 159876 198172 171140 198200
rect 159876 198160 159882 198172
rect 171134 198160 171140 198172
rect 171192 198160 171198 198212
rect 174906 198160 174912 198212
rect 174964 198200 174970 198212
rect 215478 198200 215484 198212
rect 174964 198172 215484 198200
rect 174964 198160 174970 198172
rect 215478 198160 215484 198172
rect 215536 198160 215542 198212
rect 108942 198092 108948 198144
rect 109000 198132 109006 198144
rect 143350 198132 143356 198144
rect 109000 198104 143356 198132
rect 109000 198092 109006 198104
rect 143350 198092 143356 198104
rect 143408 198092 143414 198144
rect 148410 198092 148416 198144
rect 148468 198132 148474 198144
rect 156230 198132 156236 198144
rect 148468 198104 156236 198132
rect 148468 198092 148474 198104
rect 156230 198092 156236 198104
rect 156288 198092 156294 198144
rect 163406 198092 163412 198144
rect 163464 198132 163470 198144
rect 168098 198132 168104 198144
rect 163464 198104 168104 198132
rect 163464 198092 163470 198104
rect 168098 198092 168104 198104
rect 168156 198092 168162 198144
rect 170030 198092 170036 198144
rect 170088 198132 170094 198144
rect 211798 198132 211804 198144
rect 170088 198104 211804 198132
rect 170088 198092 170094 198104
rect 211798 198092 211804 198104
rect 211856 198092 211862 198144
rect 103146 198024 103152 198076
rect 103204 198064 103210 198076
rect 134058 198064 134064 198076
rect 103204 198036 134064 198064
rect 103204 198024 103210 198036
rect 134058 198024 134064 198036
rect 134116 198024 134122 198076
rect 149330 198024 149336 198076
rect 149388 198064 149394 198076
rect 149882 198064 149888 198076
rect 149388 198036 149888 198064
rect 149388 198024 149394 198036
rect 149882 198024 149888 198036
rect 149940 198024 149946 198076
rect 155770 198024 155776 198076
rect 155828 198064 155834 198076
rect 155828 198036 164924 198064
rect 155828 198024 155834 198036
rect 140774 197956 140780 198008
rect 140832 197996 140838 198008
rect 145282 197996 145288 198008
rect 140832 197968 145288 197996
rect 140832 197956 140838 197968
rect 145282 197956 145288 197968
rect 145340 197956 145346 198008
rect 146202 197956 146208 198008
rect 146260 197996 146266 198008
rect 159450 197996 159456 198008
rect 146260 197968 159456 197996
rect 146260 197956 146266 197968
rect 159450 197956 159456 197968
rect 159508 197956 159514 198008
rect 164896 197996 164924 198036
rect 171502 198024 171508 198076
rect 171560 198064 171566 198076
rect 171870 198064 171876 198076
rect 171560 198036 171876 198064
rect 171560 198024 171566 198036
rect 171870 198024 171876 198036
rect 171928 198024 171934 198076
rect 176120 198036 176608 198064
rect 170490 197996 170496 198008
rect 164896 197968 170496 197996
rect 170490 197956 170496 197968
rect 170548 197956 170554 198008
rect 176120 197996 176148 198036
rect 171796 197968 176148 197996
rect 176580 197996 176608 198036
rect 176654 198024 176660 198076
rect 176712 198064 176718 198076
rect 181162 198064 181168 198076
rect 176712 198036 181168 198064
rect 176712 198024 176718 198036
rect 181162 198024 181168 198036
rect 181220 198024 181226 198076
rect 181438 198024 181444 198076
rect 181496 198064 181502 198076
rect 214374 198064 214380 198076
rect 181496 198036 214380 198064
rect 181496 198024 181502 198036
rect 214374 198024 214380 198036
rect 214432 198024 214438 198076
rect 211430 197996 211436 198008
rect 176580 197968 211436 197996
rect 124858 197888 124864 197940
rect 124916 197928 124922 197940
rect 124916 197900 142752 197928
rect 124916 197888 124922 197900
rect 108390 197820 108396 197872
rect 108448 197860 108454 197872
rect 142522 197860 142528 197872
rect 108448 197832 142528 197860
rect 108448 197820 108454 197832
rect 142522 197820 142528 197832
rect 142580 197820 142586 197872
rect 142724 197860 142752 197900
rect 149606 197888 149612 197940
rect 149664 197928 149670 197940
rect 149882 197928 149888 197940
rect 149664 197900 149888 197928
rect 149664 197888 149670 197900
rect 149882 197888 149888 197900
rect 149940 197888 149946 197940
rect 161566 197888 161572 197940
rect 161624 197928 161630 197940
rect 171796 197928 171824 197968
rect 211430 197956 211436 197968
rect 211488 197956 211494 198008
rect 161624 197900 171824 197928
rect 161624 197888 161630 197900
rect 174170 197888 174176 197940
rect 174228 197928 174234 197940
rect 187050 197928 187056 197940
rect 174228 197900 187056 197928
rect 174228 197888 174234 197900
rect 187050 197888 187056 197900
rect 187108 197888 187114 197940
rect 144638 197860 144644 197872
rect 142724 197832 144644 197860
rect 144638 197820 144644 197832
rect 144696 197820 144702 197872
rect 149238 197820 149244 197872
rect 149296 197860 149302 197872
rect 171042 197860 171048 197872
rect 149296 197832 171048 197860
rect 149296 197820 149302 197832
rect 171042 197820 171048 197832
rect 171100 197820 171106 197872
rect 181438 197860 181444 197872
rect 179386 197832 181444 197860
rect 124950 197752 124956 197804
rect 125008 197792 125014 197804
rect 144454 197792 144460 197804
rect 125008 197764 144460 197792
rect 125008 197752 125014 197764
rect 144454 197752 144460 197764
rect 144512 197752 144518 197804
rect 149974 197752 149980 197804
rect 150032 197792 150038 197804
rect 151078 197792 151084 197804
rect 150032 197764 151084 197792
rect 150032 197752 150038 197764
rect 151078 197752 151084 197764
rect 151136 197752 151142 197804
rect 160278 197752 160284 197804
rect 160336 197792 160342 197804
rect 169754 197792 169760 197804
rect 160336 197764 169760 197792
rect 160336 197752 160342 197764
rect 169754 197752 169760 197764
rect 169812 197752 169818 197804
rect 171134 197752 171140 197804
rect 171192 197792 171198 197804
rect 172146 197792 172152 197804
rect 171192 197764 172152 197792
rect 171192 197752 171198 197764
rect 172146 197752 172152 197764
rect 172204 197752 172210 197804
rect 160738 197684 160744 197736
rect 160796 197724 160802 197736
rect 173802 197724 173808 197736
rect 160796 197696 173808 197724
rect 160796 197684 160802 197696
rect 173802 197684 173808 197696
rect 173860 197684 173866 197736
rect 176378 197684 176384 197736
rect 176436 197724 176442 197736
rect 177666 197724 177672 197736
rect 176436 197696 177672 197724
rect 176436 197684 176442 197696
rect 177666 197684 177672 197696
rect 177724 197684 177730 197736
rect 129182 197616 129188 197668
rect 129240 197656 129246 197668
rect 143626 197656 143632 197668
rect 129240 197628 143632 197656
rect 129240 197616 129246 197628
rect 143626 197616 143632 197628
rect 143684 197616 143690 197668
rect 157426 197616 157432 197668
rect 157484 197656 157490 197668
rect 171870 197656 171876 197668
rect 157484 197628 171876 197656
rect 157484 197616 157490 197628
rect 171870 197616 171876 197628
rect 171928 197616 171934 197668
rect 179386 197656 179414 197832
rect 181438 197820 181444 197832
rect 181496 197820 181502 197872
rect 173866 197628 179414 197656
rect 149790 197548 149796 197600
rect 149848 197588 149854 197600
rect 150066 197588 150072 197600
rect 149848 197560 150072 197588
rect 149848 197548 149854 197560
rect 150066 197548 150072 197560
rect 150124 197548 150130 197600
rect 156046 197548 156052 197600
rect 156104 197588 156110 197600
rect 156104 197560 166994 197588
rect 156104 197548 156110 197560
rect 149790 197412 149796 197464
rect 149848 197452 149854 197464
rect 153930 197452 153936 197464
rect 149848 197424 153936 197452
rect 149848 197412 149854 197424
rect 153930 197412 153936 197424
rect 153988 197412 153994 197464
rect 133506 197344 133512 197396
rect 133564 197384 133570 197396
rect 141326 197384 141332 197396
rect 133564 197356 141332 197384
rect 133564 197344 133570 197356
rect 141326 197344 141332 197356
rect 141384 197344 141390 197396
rect 156046 197344 156052 197396
rect 156104 197384 156110 197396
rect 156598 197384 156604 197396
rect 156104 197356 156604 197384
rect 156104 197344 156110 197356
rect 156598 197344 156604 197356
rect 156656 197344 156662 197396
rect 166966 197384 166994 197560
rect 167178 197548 167184 197600
rect 167236 197588 167242 197600
rect 173866 197588 173894 197628
rect 188338 197588 188344 197600
rect 167236 197560 173894 197588
rect 176626 197560 188344 197588
rect 167236 197548 167242 197560
rect 169754 197480 169760 197532
rect 169812 197520 169818 197532
rect 175182 197520 175188 197532
rect 169812 197492 175188 197520
rect 169812 197480 169818 197492
rect 175182 197480 175188 197492
rect 175240 197480 175246 197532
rect 167822 197412 167828 197464
rect 167880 197452 167886 197464
rect 168374 197452 168380 197464
rect 167880 197424 168380 197452
rect 167880 197412 167886 197424
rect 168374 197412 168380 197424
rect 168432 197412 168438 197464
rect 173894 197412 173900 197464
rect 173952 197452 173958 197464
rect 174078 197452 174084 197464
rect 173952 197424 174084 197452
rect 173952 197412 173958 197424
rect 174078 197412 174084 197424
rect 174136 197412 174142 197464
rect 175366 197412 175372 197464
rect 175424 197452 175430 197464
rect 176102 197452 176108 197464
rect 175424 197424 176108 197452
rect 175424 197412 175430 197424
rect 176102 197412 176108 197424
rect 176160 197412 176166 197464
rect 176626 197384 176654 197560
rect 188338 197548 188344 197560
rect 188396 197548 188402 197600
rect 166966 197356 176654 197384
rect 177114 197344 177120 197396
rect 177172 197384 177178 197396
rect 182450 197384 182456 197396
rect 177172 197356 182456 197384
rect 177172 197344 177178 197356
rect 182450 197344 182456 197356
rect 182508 197344 182514 197396
rect 105630 197276 105636 197328
rect 105688 197316 105694 197328
rect 130286 197316 130292 197328
rect 105688 197288 130292 197316
rect 105688 197276 105694 197288
rect 130286 197276 130292 197288
rect 130344 197276 130350 197328
rect 131850 197276 131856 197328
rect 131908 197316 131914 197328
rect 139486 197316 139492 197328
rect 131908 197288 139492 197316
rect 131908 197276 131914 197288
rect 139486 197276 139492 197288
rect 139544 197276 139550 197328
rect 139578 197276 139584 197328
rect 139636 197316 139642 197328
rect 139946 197316 139952 197328
rect 139636 197288 139952 197316
rect 139636 197276 139642 197288
rect 139946 197276 139952 197288
rect 140004 197276 140010 197328
rect 141234 197276 141240 197328
rect 141292 197316 141298 197328
rect 141878 197316 141884 197328
rect 141292 197288 141884 197316
rect 141292 197276 141298 197288
rect 141878 197276 141884 197288
rect 141936 197276 141942 197328
rect 166350 197276 166356 197328
rect 166408 197316 166414 197328
rect 179414 197316 179420 197328
rect 166408 197288 179420 197316
rect 166408 197276 166414 197288
rect 179414 197276 179420 197288
rect 179472 197276 179478 197328
rect 121086 197208 121092 197260
rect 121144 197248 121150 197260
rect 145834 197248 145840 197260
rect 121144 197220 145840 197248
rect 121144 197208 121150 197220
rect 145834 197208 145840 197220
rect 145892 197208 145898 197260
rect 157242 197208 157248 197260
rect 157300 197248 157306 197260
rect 158990 197248 158996 197260
rect 157300 197220 158996 197248
rect 157300 197208 157306 197220
rect 158990 197208 158996 197220
rect 159048 197208 159054 197260
rect 160830 197208 160836 197260
rect 160888 197248 160894 197260
rect 180426 197248 180432 197260
rect 160888 197220 180432 197248
rect 160888 197208 160894 197220
rect 180426 197208 180432 197220
rect 180484 197208 180490 197260
rect 108298 197140 108304 197192
rect 108356 197180 108362 197192
rect 137370 197180 137376 197192
rect 108356 197152 137376 197180
rect 108356 197140 108362 197152
rect 137370 197140 137376 197152
rect 137428 197140 137434 197192
rect 137462 197140 137468 197192
rect 137520 197180 137526 197192
rect 138106 197180 138112 197192
rect 137520 197152 138112 197180
rect 137520 197140 137526 197152
rect 138106 197140 138112 197152
rect 138164 197140 138170 197192
rect 139762 197140 139768 197192
rect 139820 197180 139826 197192
rect 140038 197180 140044 197192
rect 139820 197152 140044 197180
rect 139820 197140 139826 197152
rect 140038 197140 140044 197152
rect 140096 197140 140102 197192
rect 141878 197140 141884 197192
rect 141936 197180 141942 197192
rect 142338 197180 142344 197192
rect 141936 197152 142344 197180
rect 141936 197140 141942 197152
rect 142338 197140 142344 197152
rect 142396 197140 142402 197192
rect 160002 197140 160008 197192
rect 160060 197180 160066 197192
rect 160646 197180 160652 197192
rect 160060 197152 160652 197180
rect 160060 197140 160066 197152
rect 160646 197140 160652 197152
rect 160704 197140 160710 197192
rect 162762 197140 162768 197192
rect 162820 197180 162826 197192
rect 167914 197180 167920 197192
rect 162820 197152 167920 197180
rect 162820 197140 162826 197152
rect 167914 197140 167920 197152
rect 167972 197140 167978 197192
rect 168098 197140 168104 197192
rect 168156 197180 168162 197192
rect 197354 197180 197360 197192
rect 168156 197152 197360 197180
rect 168156 197140 168162 197152
rect 197354 197140 197360 197152
rect 197412 197140 197418 197192
rect 119062 197072 119068 197124
rect 119120 197112 119126 197124
rect 151814 197112 151820 197124
rect 119120 197084 151820 197112
rect 119120 197072 119126 197084
rect 151814 197072 151820 197084
rect 151872 197072 151878 197124
rect 164694 197072 164700 197124
rect 164752 197112 164758 197124
rect 199654 197112 199660 197124
rect 164752 197084 199660 197112
rect 164752 197072 164758 197084
rect 199654 197072 199660 197084
rect 199712 197072 199718 197124
rect 112990 197004 112996 197056
rect 113048 197044 113054 197056
rect 142062 197044 142068 197056
rect 113048 197016 142068 197044
rect 113048 197004 113054 197016
rect 142062 197004 142068 197016
rect 142120 197004 142126 197056
rect 171226 197004 171232 197056
rect 171284 197044 171290 197056
rect 201678 197044 201684 197056
rect 171284 197016 201684 197044
rect 171284 197004 171290 197016
rect 201678 197004 201684 197016
rect 201736 197004 201742 197056
rect 111518 196936 111524 196988
rect 111576 196976 111582 196988
rect 143258 196976 143264 196988
rect 111576 196948 143264 196976
rect 111576 196936 111582 196948
rect 143258 196936 143264 196948
rect 143316 196936 143322 196988
rect 154666 196936 154672 196988
rect 154724 196976 154730 196988
rect 155402 196976 155408 196988
rect 154724 196948 155408 196976
rect 154724 196936 154730 196948
rect 155402 196936 155408 196948
rect 155460 196936 155466 196988
rect 159082 196936 159088 196988
rect 159140 196976 159146 196988
rect 159910 196976 159916 196988
rect 159140 196948 159916 196976
rect 159140 196936 159146 196948
rect 159910 196936 159916 196948
rect 159968 196936 159974 196988
rect 164418 196936 164424 196988
rect 164476 196976 164482 196988
rect 197538 196976 197544 196988
rect 164476 196948 197544 196976
rect 164476 196936 164482 196948
rect 197538 196936 197544 196948
rect 197596 196936 197602 196988
rect 112714 196868 112720 196920
rect 112772 196908 112778 196920
rect 132862 196908 132868 196920
rect 112772 196880 132868 196908
rect 112772 196868 112778 196880
rect 132862 196868 132868 196880
rect 132920 196868 132926 196920
rect 137278 196868 137284 196920
rect 137336 196908 137342 196920
rect 138382 196908 138388 196920
rect 137336 196880 138388 196908
rect 137336 196868 137342 196880
rect 138382 196868 138388 196880
rect 138440 196868 138446 196920
rect 139670 196868 139676 196920
rect 139728 196908 139734 196920
rect 140498 196908 140504 196920
rect 139728 196880 140504 196908
rect 139728 196868 139734 196880
rect 140498 196868 140504 196880
rect 140556 196868 140562 196920
rect 143442 196868 143448 196920
rect 143500 196908 143506 196920
rect 143810 196908 143816 196920
rect 143500 196880 143816 196908
rect 143500 196868 143506 196880
rect 143810 196868 143816 196880
rect 143868 196868 143874 196920
rect 155310 196868 155316 196920
rect 155368 196908 155374 196920
rect 189166 196908 189172 196920
rect 155368 196880 189172 196908
rect 155368 196868 155374 196880
rect 189166 196868 189172 196880
rect 189224 196868 189230 196920
rect 114278 196800 114284 196852
rect 114336 196840 114342 196852
rect 146110 196840 146116 196852
rect 114336 196812 146116 196840
rect 114336 196800 114342 196812
rect 146110 196800 146116 196812
rect 146168 196800 146174 196852
rect 160370 196800 160376 196852
rect 160428 196840 160434 196852
rect 160554 196840 160560 196852
rect 160428 196812 160560 196840
rect 160428 196800 160434 196812
rect 160554 196800 160560 196812
rect 160612 196800 160618 196852
rect 161934 196800 161940 196852
rect 161992 196840 161998 196852
rect 196342 196840 196348 196852
rect 161992 196812 196348 196840
rect 161992 196800 161998 196812
rect 196342 196800 196348 196812
rect 196400 196800 196406 196852
rect 111150 196732 111156 196784
rect 111208 196772 111214 196784
rect 133138 196772 133144 196784
rect 111208 196744 133144 196772
rect 111208 196732 111214 196744
rect 133138 196732 133144 196744
rect 133196 196732 133202 196784
rect 139854 196732 139860 196784
rect 139912 196772 139918 196784
rect 140314 196772 140320 196784
rect 139912 196744 140320 196772
rect 139912 196732 139918 196744
rect 140314 196732 140320 196744
rect 140372 196732 140378 196784
rect 164326 196732 164332 196784
rect 164384 196772 164390 196784
rect 165338 196772 165344 196784
rect 164384 196744 165344 196772
rect 164384 196732 164390 196744
rect 165338 196732 165344 196744
rect 165396 196732 165402 196784
rect 172790 196732 172796 196784
rect 172848 196772 172854 196784
rect 173342 196772 173348 196784
rect 172848 196744 173348 196772
rect 172848 196732 172854 196744
rect 173342 196732 173348 196744
rect 173400 196732 173406 196784
rect 175550 196732 175556 196784
rect 175608 196772 175614 196784
rect 176470 196772 176476 196784
rect 175608 196744 176476 196772
rect 175608 196732 175614 196744
rect 176470 196732 176476 196744
rect 176528 196732 176534 196784
rect 177114 196732 177120 196784
rect 177172 196772 177178 196784
rect 177390 196772 177396 196784
rect 177172 196744 177396 196772
rect 177172 196732 177178 196744
rect 177390 196732 177396 196744
rect 177448 196732 177454 196784
rect 181162 196732 181168 196784
rect 181220 196772 181226 196784
rect 215294 196772 215300 196784
rect 181220 196744 215300 196772
rect 181220 196732 181226 196744
rect 215294 196732 215300 196744
rect 215352 196732 215358 196784
rect 105538 196664 105544 196716
rect 105596 196704 105602 196716
rect 136634 196704 136640 196716
rect 105596 196676 136640 196704
rect 105596 196664 105602 196676
rect 136634 196664 136640 196676
rect 136692 196664 136698 196716
rect 138566 196664 138572 196716
rect 138624 196704 138630 196716
rect 138842 196704 138848 196716
rect 138624 196676 138848 196704
rect 138624 196664 138630 196676
rect 138842 196664 138848 196676
rect 138900 196664 138906 196716
rect 139946 196664 139952 196716
rect 140004 196704 140010 196716
rect 140406 196704 140412 196716
rect 140004 196676 140412 196704
rect 140004 196664 140010 196676
rect 140406 196664 140412 196676
rect 140464 196664 140470 196716
rect 141418 196664 141424 196716
rect 141476 196704 141482 196716
rect 143718 196704 143724 196716
rect 141476 196676 143724 196704
rect 141476 196664 141482 196676
rect 143718 196664 143724 196676
rect 143776 196664 143782 196716
rect 148686 196664 148692 196716
rect 148744 196704 148750 196716
rect 155494 196704 155500 196716
rect 148744 196676 155500 196704
rect 148744 196664 148750 196676
rect 155494 196664 155500 196676
rect 155552 196664 155558 196716
rect 157518 196664 157524 196716
rect 157576 196704 157582 196716
rect 157702 196704 157708 196716
rect 157576 196676 157708 196704
rect 157576 196664 157582 196676
rect 157702 196664 157708 196676
rect 157760 196664 157766 196716
rect 160278 196664 160284 196716
rect 160336 196704 160342 196716
rect 160922 196704 160928 196716
rect 160336 196676 160928 196704
rect 160336 196664 160342 196676
rect 160922 196664 160928 196676
rect 160980 196664 160986 196716
rect 161382 196664 161388 196716
rect 161440 196704 161446 196716
rect 162762 196704 162768 196716
rect 161440 196676 162768 196704
rect 161440 196664 161446 196676
rect 162762 196664 162768 196676
rect 162820 196664 162826 196716
rect 164510 196664 164516 196716
rect 164568 196704 164574 196716
rect 165614 196704 165620 196716
rect 164568 196676 165620 196704
rect 164568 196664 164574 196676
rect 165614 196664 165620 196676
rect 165672 196664 165678 196716
rect 165706 196664 165712 196716
rect 165764 196704 165770 196716
rect 166718 196704 166724 196716
rect 165764 196676 166724 196704
rect 165764 196664 165770 196676
rect 166718 196664 166724 196676
rect 166776 196664 166782 196716
rect 166994 196664 167000 196716
rect 167052 196704 167058 196716
rect 168190 196704 168196 196716
rect 167052 196676 168196 196704
rect 167052 196664 167058 196676
rect 168190 196664 168196 196676
rect 168248 196664 168254 196716
rect 168466 196664 168472 196716
rect 168524 196704 168530 196716
rect 169294 196704 169300 196716
rect 168524 196676 169300 196704
rect 168524 196664 168530 196676
rect 169294 196664 169300 196676
rect 169352 196664 169358 196716
rect 169570 196664 169576 196716
rect 169628 196704 169634 196716
rect 169846 196704 169852 196716
rect 169628 196676 169852 196704
rect 169628 196664 169634 196676
rect 169846 196664 169852 196676
rect 169904 196664 169910 196716
rect 172882 196664 172888 196716
rect 172940 196704 172946 196716
rect 173526 196704 173532 196716
rect 172940 196676 173532 196704
rect 172940 196664 172946 196676
rect 173526 196664 173532 196676
rect 173584 196664 173590 196716
rect 177022 196664 177028 196716
rect 177080 196704 177086 196716
rect 177574 196704 177580 196716
rect 177080 196676 177580 196704
rect 177080 196664 177086 196676
rect 177574 196664 177580 196676
rect 177632 196664 177638 196716
rect 181990 196664 181996 196716
rect 182048 196704 182054 196716
rect 215662 196704 215668 196716
rect 182048 196676 215668 196704
rect 182048 196664 182054 196676
rect 215662 196664 215668 196676
rect 215720 196664 215726 196716
rect 97902 196596 97908 196648
rect 97960 196636 97966 196648
rect 97960 196608 122834 196636
rect 97960 196596 97966 196608
rect 122806 196568 122834 196608
rect 140866 196596 140872 196648
rect 140924 196636 140930 196648
rect 141786 196636 141792 196648
rect 140924 196608 141792 196636
rect 140924 196596 140930 196608
rect 141786 196596 141792 196608
rect 141844 196596 141850 196648
rect 142982 196596 142988 196648
rect 143040 196636 143046 196648
rect 143166 196636 143172 196648
rect 143040 196608 143172 196636
rect 143040 196596 143046 196608
rect 143166 196596 143172 196608
rect 143224 196596 143230 196648
rect 147214 196596 147220 196648
rect 147272 196636 147278 196648
rect 151354 196636 151360 196648
rect 147272 196608 151360 196636
rect 147272 196596 147278 196608
rect 151354 196596 151360 196608
rect 151412 196596 151418 196648
rect 151814 196596 151820 196648
rect 151872 196636 151878 196648
rect 152366 196636 152372 196648
rect 151872 196608 152372 196636
rect 151872 196596 151878 196608
rect 152366 196596 152372 196608
rect 152424 196596 152430 196648
rect 152642 196596 152648 196648
rect 152700 196636 152706 196648
rect 152918 196636 152924 196648
rect 152700 196608 152924 196636
rect 152700 196596 152706 196608
rect 152918 196596 152924 196608
rect 152976 196596 152982 196648
rect 154758 196596 154764 196648
rect 154816 196636 154822 196648
rect 155678 196636 155684 196648
rect 154816 196608 155684 196636
rect 154816 196596 154822 196608
rect 155678 196596 155684 196608
rect 155736 196596 155742 196648
rect 165982 196596 165988 196648
rect 166040 196636 166046 196648
rect 166902 196636 166908 196648
rect 166040 196608 166908 196636
rect 166040 196596 166046 196608
rect 166902 196596 166908 196608
rect 166960 196596 166966 196648
rect 167638 196596 167644 196648
rect 167696 196636 167702 196648
rect 170030 196636 170036 196648
rect 167696 196608 170036 196636
rect 167696 196596 167702 196608
rect 170030 196596 170036 196608
rect 170088 196596 170094 196648
rect 170122 196596 170128 196648
rect 170180 196636 170186 196648
rect 216674 196636 216680 196648
rect 170180 196608 216680 196636
rect 170180 196596 170186 196608
rect 216674 196596 216680 196608
rect 216732 196596 216738 196648
rect 133506 196568 133512 196580
rect 122806 196540 133512 196568
rect 133506 196528 133512 196540
rect 133564 196528 133570 196580
rect 149330 196528 149336 196580
rect 149388 196568 149394 196580
rect 150250 196568 150256 196580
rect 149388 196540 150256 196568
rect 149388 196528 149394 196540
rect 150250 196528 150256 196540
rect 150308 196528 150314 196580
rect 154942 196528 154948 196580
rect 155000 196568 155006 196580
rect 156598 196568 156604 196580
rect 155000 196540 156604 196568
rect 155000 196528 155006 196540
rect 156598 196528 156604 196540
rect 156656 196528 156662 196580
rect 176654 196528 176660 196580
rect 176712 196568 176718 196580
rect 177206 196568 177212 196580
rect 176712 196540 177212 196568
rect 176712 196528 176718 196540
rect 177206 196528 177212 196540
rect 177264 196528 177270 196580
rect 177298 196528 177304 196580
rect 177356 196568 177362 196580
rect 178218 196568 178224 196580
rect 177356 196540 178224 196568
rect 177356 196528 177362 196540
rect 178218 196528 178224 196540
rect 178276 196528 178282 196580
rect 126698 196460 126704 196512
rect 126756 196500 126762 196512
rect 146570 196500 146576 196512
rect 126756 196472 146576 196500
rect 126756 196460 126762 196472
rect 146570 196460 146576 196472
rect 146628 196460 146634 196512
rect 164878 196460 164884 196512
rect 164936 196500 164942 196512
rect 165430 196500 165436 196512
rect 164936 196472 165436 196500
rect 164936 196460 164942 196472
rect 165430 196460 165436 196472
rect 165488 196460 165494 196512
rect 169846 196460 169852 196512
rect 169904 196500 169910 196512
rect 170214 196500 170220 196512
rect 169904 196472 170220 196500
rect 169904 196460 169910 196472
rect 170214 196460 170220 196472
rect 170272 196460 170278 196512
rect 175826 196460 175832 196512
rect 175884 196500 175890 196512
rect 182266 196500 182272 196512
rect 175884 196472 182272 196500
rect 175884 196460 175890 196472
rect 182266 196460 182272 196472
rect 182324 196460 182330 196512
rect 129918 196392 129924 196444
rect 129976 196432 129982 196444
rect 140590 196432 140596 196444
rect 129976 196404 140596 196432
rect 129976 196392 129982 196404
rect 140590 196392 140596 196404
rect 140648 196392 140654 196444
rect 162946 196392 162952 196444
rect 163004 196432 163010 196444
rect 163222 196432 163228 196444
rect 163004 196404 163228 196432
rect 163004 196392 163010 196404
rect 163222 196392 163228 196404
rect 163280 196392 163286 196444
rect 169018 196392 169024 196444
rect 169076 196392 169082 196444
rect 126606 196324 126612 196376
rect 126664 196364 126670 196376
rect 148318 196364 148324 196376
rect 126664 196336 148324 196364
rect 126664 196324 126670 196336
rect 148318 196324 148324 196336
rect 148376 196324 148382 196376
rect 161934 196324 161940 196376
rect 161992 196364 161998 196376
rect 162670 196364 162676 196376
rect 161992 196336 162676 196364
rect 161992 196324 161998 196336
rect 162670 196324 162676 196336
rect 162728 196324 162734 196376
rect 132862 196256 132868 196308
rect 132920 196296 132926 196308
rect 144546 196296 144552 196308
rect 132920 196268 144552 196296
rect 132920 196256 132926 196268
rect 144546 196256 144552 196268
rect 144604 196256 144610 196308
rect 144914 196256 144920 196308
rect 144972 196296 144978 196308
rect 145834 196296 145840 196308
rect 144972 196268 145840 196296
rect 144972 196256 144978 196268
rect 145834 196256 145840 196268
rect 145892 196256 145898 196308
rect 151906 196256 151912 196308
rect 151964 196296 151970 196308
rect 153010 196296 153016 196308
rect 151964 196268 153016 196296
rect 151964 196256 151970 196268
rect 153010 196256 153016 196268
rect 153068 196256 153074 196308
rect 157978 196256 157984 196308
rect 158036 196296 158042 196308
rect 159542 196296 159548 196308
rect 158036 196268 159548 196296
rect 158036 196256 158042 196268
rect 159542 196256 159548 196268
rect 159600 196256 159606 196308
rect 131022 196188 131028 196240
rect 131080 196228 131086 196240
rect 134702 196228 134708 196240
rect 131080 196200 134708 196228
rect 131080 196188 131086 196200
rect 134702 196188 134708 196200
rect 134760 196188 134766 196240
rect 143902 196188 143908 196240
rect 143960 196228 143966 196240
rect 144086 196228 144092 196240
rect 143960 196200 144092 196228
rect 143960 196188 143966 196200
rect 144086 196188 144092 196200
rect 144144 196188 144150 196240
rect 157794 196188 157800 196240
rect 157852 196228 157858 196240
rect 158438 196228 158444 196240
rect 157852 196200 158444 196228
rect 157852 196188 157858 196200
rect 158438 196188 158444 196200
rect 158496 196188 158502 196240
rect 133138 196120 133144 196172
rect 133196 196160 133202 196172
rect 143994 196160 144000 196172
rect 133196 196132 144000 196160
rect 133196 196120 133202 196132
rect 143994 196120 144000 196132
rect 144052 196120 144058 196172
rect 144914 196120 144920 196172
rect 144972 196160 144978 196172
rect 146478 196160 146484 196172
rect 144972 196132 146484 196160
rect 144972 196120 144978 196132
rect 146478 196120 146484 196132
rect 146536 196120 146542 196172
rect 161750 196120 161756 196172
rect 161808 196120 161814 196172
rect 168558 196120 168564 196172
rect 168616 196160 168622 196172
rect 169036 196160 169064 196392
rect 169386 196324 169392 196376
rect 169444 196364 169450 196376
rect 183002 196364 183008 196376
rect 169444 196336 183008 196364
rect 169444 196324 169450 196336
rect 183002 196324 183008 196336
rect 183060 196324 183066 196376
rect 176930 196256 176936 196308
rect 176988 196296 176994 196308
rect 177482 196296 177488 196308
rect 176988 196268 177488 196296
rect 176988 196256 176994 196268
rect 177482 196256 177488 196268
rect 177540 196256 177546 196308
rect 171042 196188 171048 196240
rect 171100 196228 171106 196240
rect 178954 196228 178960 196240
rect 171100 196200 178960 196228
rect 171100 196188 171106 196200
rect 178954 196188 178960 196200
rect 179012 196188 179018 196240
rect 168616 196132 169064 196160
rect 168616 196120 168622 196132
rect 176838 196120 176844 196172
rect 176896 196160 176902 196172
rect 177758 196160 177764 196172
rect 176896 196132 177764 196160
rect 176896 196120 176902 196132
rect 177758 196120 177764 196132
rect 177816 196120 177822 196172
rect 141602 196052 141608 196104
rect 141660 196092 141666 196104
rect 143902 196092 143908 196104
rect 141660 196064 143908 196092
rect 141660 196052 141666 196064
rect 143902 196052 143908 196064
rect 143960 196052 143966 196104
rect 138474 195984 138480 196036
rect 138532 196024 138538 196036
rect 138658 196024 138664 196036
rect 138532 195996 138664 196024
rect 138532 195984 138538 195996
rect 138658 195984 138664 195996
rect 138716 195984 138722 196036
rect 145466 195984 145472 196036
rect 145524 196024 145530 196036
rect 146018 196024 146024 196036
rect 145524 195996 146024 196024
rect 145524 195984 145530 195996
rect 146018 195984 146024 195996
rect 146076 195984 146082 196036
rect 120718 195916 120724 195968
rect 120776 195956 120782 195968
rect 145190 195956 145196 195968
rect 120776 195928 145196 195956
rect 120776 195916 120782 195928
rect 145190 195916 145196 195928
rect 145248 195916 145254 195968
rect 145374 195916 145380 195968
rect 145432 195956 145438 195968
rect 146570 195956 146576 195968
rect 145432 195928 146576 195956
rect 145432 195916 145438 195928
rect 146570 195916 146576 195928
rect 146628 195916 146634 195968
rect 153470 195916 153476 195968
rect 153528 195956 153534 195968
rect 153654 195956 153660 195968
rect 153528 195928 153660 195956
rect 153528 195916 153534 195928
rect 153654 195916 153660 195928
rect 153712 195916 153718 195968
rect 156230 195916 156236 195968
rect 156288 195956 156294 195968
rect 157978 195956 157984 195968
rect 156288 195928 157984 195956
rect 156288 195916 156294 195928
rect 157978 195916 157984 195928
rect 158036 195916 158042 195968
rect 161658 195916 161664 195968
rect 161716 195956 161722 195968
rect 161768 195956 161796 196120
rect 161716 195928 161796 195956
rect 161716 195916 161722 195928
rect 169386 195916 169392 195968
rect 169444 195956 169450 195968
rect 183094 195956 183100 195968
rect 169444 195928 183100 195956
rect 169444 195916 169450 195928
rect 183094 195916 183100 195928
rect 183152 195916 183158 195968
rect 123478 195848 123484 195900
rect 123536 195888 123542 195900
rect 149146 195888 149152 195900
rect 123536 195860 149152 195888
rect 123536 195848 123542 195860
rect 149146 195848 149152 195860
rect 149204 195848 149210 195900
rect 157426 195848 157432 195900
rect 157484 195888 157490 195900
rect 158070 195888 158076 195900
rect 157484 195860 158076 195888
rect 157484 195848 157490 195860
rect 158070 195848 158076 195860
rect 158128 195848 158134 195900
rect 158990 195848 158996 195900
rect 159048 195888 159054 195900
rect 159266 195888 159272 195900
rect 159048 195860 159272 195888
rect 159048 195848 159054 195860
rect 159266 195848 159272 195860
rect 159324 195848 159330 195900
rect 161290 195848 161296 195900
rect 161348 195888 161354 195900
rect 176194 195888 176200 195900
rect 161348 195860 176200 195888
rect 161348 195848 161354 195860
rect 176194 195848 176200 195860
rect 176252 195848 176258 195900
rect 119890 195780 119896 195832
rect 119948 195820 119954 195832
rect 148962 195820 148968 195832
rect 119948 195792 148968 195820
rect 119948 195780 119954 195792
rect 148962 195780 148968 195792
rect 149020 195780 149026 195832
rect 153470 195780 153476 195832
rect 153528 195820 153534 195832
rect 154298 195820 154304 195832
rect 153528 195792 154304 195820
rect 153528 195780 153534 195792
rect 154298 195780 154304 195792
rect 154356 195780 154362 195832
rect 156230 195780 156236 195832
rect 156288 195820 156294 195832
rect 156506 195820 156512 195832
rect 156288 195792 156512 195820
rect 156288 195780 156294 195792
rect 156506 195780 156512 195792
rect 156564 195780 156570 195832
rect 175182 195780 175188 195832
rect 175240 195820 175246 195832
rect 194594 195820 194600 195832
rect 175240 195792 194600 195820
rect 175240 195780 175246 195792
rect 194594 195780 194600 195792
rect 194652 195780 194658 195832
rect 118510 195712 118516 195764
rect 118568 195752 118574 195764
rect 148134 195752 148140 195764
rect 118568 195724 148140 195752
rect 118568 195712 118574 195724
rect 148134 195712 148140 195724
rect 148192 195712 148198 195764
rect 150986 195712 150992 195764
rect 151044 195752 151050 195764
rect 151630 195752 151636 195764
rect 151044 195724 151636 195752
rect 151044 195712 151050 195724
rect 151630 195712 151636 195724
rect 151688 195712 151694 195764
rect 173802 195712 173808 195764
rect 173860 195752 173866 195764
rect 194686 195752 194692 195764
rect 173860 195724 194692 195752
rect 173860 195712 173866 195724
rect 194686 195712 194692 195724
rect 194744 195712 194750 195764
rect 117130 195644 117136 195696
rect 117188 195684 117194 195696
rect 147858 195684 147864 195696
rect 117188 195656 147864 195684
rect 117188 195644 117194 195656
rect 147858 195644 147864 195656
rect 147916 195644 147922 195696
rect 172054 195644 172060 195696
rect 172112 195684 172118 195696
rect 193398 195684 193404 195696
rect 172112 195656 173664 195684
rect 172112 195644 172118 195656
rect 111334 195576 111340 195628
rect 111392 195616 111398 195628
rect 128446 195616 128452 195628
rect 111392 195588 128452 195616
rect 111392 195576 111398 195588
rect 128446 195576 128452 195588
rect 128504 195576 128510 195628
rect 162486 195576 162492 195628
rect 162544 195616 162550 195628
rect 173526 195616 173532 195628
rect 162544 195588 173532 195616
rect 162544 195576 162550 195588
rect 173526 195576 173532 195588
rect 173584 195576 173590 195628
rect 173636 195616 173664 195656
rect 177316 195656 193404 195684
rect 177316 195616 177344 195656
rect 193398 195644 193404 195656
rect 193456 195644 193462 195696
rect 173636 195588 177344 195616
rect 182450 195576 182456 195628
rect 182508 195616 182514 195628
rect 203610 195616 203616 195628
rect 182508 195588 203616 195616
rect 182508 195576 182514 195588
rect 203610 195576 203616 195588
rect 203668 195576 203674 195628
rect 115658 195508 115664 195560
rect 115716 195548 115722 195560
rect 147306 195548 147312 195560
rect 115716 195520 147312 195548
rect 115716 195508 115722 195520
rect 147306 195508 147312 195520
rect 147364 195508 147370 195560
rect 158806 195508 158812 195560
rect 158864 195548 158870 195560
rect 173710 195548 173716 195560
rect 158864 195520 173716 195548
rect 158864 195508 158870 195520
rect 173710 195508 173716 195520
rect 173768 195508 173774 195560
rect 179966 195508 179972 195560
rect 180024 195548 180030 195560
rect 203702 195548 203708 195560
rect 180024 195520 203708 195548
rect 180024 195508 180030 195520
rect 203702 195508 203708 195520
rect 203760 195508 203766 195560
rect 104434 195440 104440 195492
rect 104492 195480 104498 195492
rect 137646 195480 137652 195492
rect 104492 195452 137652 195480
rect 104492 195440 104498 195452
rect 137646 195440 137652 195452
rect 137704 195440 137710 195492
rect 138290 195440 138296 195492
rect 138348 195480 138354 195492
rect 139026 195480 139032 195492
rect 138348 195452 139032 195480
rect 138348 195440 138354 195452
rect 139026 195440 139032 195452
rect 139084 195440 139090 195492
rect 154574 195440 154580 195492
rect 154632 195480 154638 195492
rect 155034 195480 155040 195492
rect 154632 195452 155040 195480
rect 154632 195440 154638 195452
rect 155034 195440 155040 195452
rect 155092 195440 155098 195492
rect 157058 195440 157064 195492
rect 157116 195480 157122 195492
rect 190454 195480 190460 195492
rect 157116 195452 190460 195480
rect 157116 195440 157122 195452
rect 190454 195440 190460 195452
rect 190512 195440 190518 195492
rect 104526 195372 104532 195424
rect 104584 195412 104590 195424
rect 123386 195412 123392 195424
rect 104584 195384 123392 195412
rect 104584 195372 104590 195384
rect 123386 195372 123392 195384
rect 123444 195372 123450 195424
rect 123570 195372 123576 195424
rect 123628 195412 123634 195424
rect 142798 195412 142804 195424
rect 123628 195384 142804 195412
rect 123628 195372 123634 195384
rect 142798 195372 142804 195384
rect 142856 195372 142862 195424
rect 149974 195412 149980 195424
rect 143460 195384 149980 195412
rect 109954 195304 109960 195356
rect 110012 195344 110018 195356
rect 110012 195316 125594 195344
rect 110012 195304 110018 195316
rect 108850 195236 108856 195288
rect 108908 195276 108914 195288
rect 125566 195276 125594 195316
rect 143350 195276 143356 195288
rect 108908 195248 115934 195276
rect 125566 195248 143356 195276
rect 108908 195236 108914 195248
rect 115906 195208 115934 195248
rect 143350 195236 143356 195248
rect 143408 195236 143414 195288
rect 123570 195208 123576 195220
rect 115906 195180 123576 195208
rect 123570 195168 123576 195180
rect 123628 195168 123634 195220
rect 128170 195168 128176 195220
rect 128228 195208 128234 195220
rect 128228 195180 142292 195208
rect 128228 195168 128234 195180
rect 132126 195100 132132 195152
rect 132184 195140 132190 195152
rect 142264 195140 142292 195180
rect 143460 195140 143488 195384
rect 149974 195372 149980 195384
rect 150032 195372 150038 195424
rect 154482 195372 154488 195424
rect 154540 195412 154546 195424
rect 187786 195412 187792 195424
rect 154540 195384 187792 195412
rect 154540 195372 154546 195384
rect 187786 195372 187792 195384
rect 187844 195372 187850 195424
rect 158714 195304 158720 195356
rect 158772 195344 158778 195356
rect 192018 195344 192024 195356
rect 158772 195316 192024 195344
rect 158772 195304 158778 195316
rect 192018 195304 192024 195316
rect 192076 195304 192082 195356
rect 159358 195236 159364 195288
rect 159416 195276 159422 195288
rect 218146 195276 218152 195288
rect 159416 195248 218152 195276
rect 159416 195236 159422 195248
rect 218146 195236 218152 195248
rect 218204 195236 218210 195288
rect 163130 195168 163136 195220
rect 163188 195208 163194 195220
rect 164050 195208 164056 195220
rect 163188 195180 164056 195208
rect 163188 195168 163194 195180
rect 164050 195168 164056 195180
rect 164108 195168 164114 195220
rect 168926 195168 168932 195220
rect 168984 195208 168990 195220
rect 183186 195208 183192 195220
rect 168984 195180 183192 195208
rect 168984 195168 168990 195180
rect 183186 195168 183192 195180
rect 183244 195168 183250 195220
rect 132184 195112 142154 195140
rect 142264 195112 143488 195140
rect 132184 195100 132190 195112
rect 123386 195032 123392 195084
rect 123444 195072 123450 195084
rect 137922 195072 137928 195084
rect 123444 195044 137928 195072
rect 123444 195032 123450 195044
rect 137922 195032 137928 195044
rect 137980 195032 137986 195084
rect 128446 194964 128452 195016
rect 128504 195004 128510 195016
rect 142126 195004 142154 195112
rect 163038 195100 163044 195152
rect 163096 195140 163102 195152
rect 163774 195140 163780 195152
rect 163096 195112 163780 195140
rect 163096 195100 163102 195112
rect 163774 195100 163780 195112
rect 163832 195100 163838 195152
rect 165982 195100 165988 195152
rect 166040 195140 166046 195152
rect 166442 195140 166448 195152
rect 166040 195112 166448 195140
rect 166040 195100 166046 195112
rect 166442 195100 166448 195112
rect 166500 195100 166506 195152
rect 173986 195100 173992 195152
rect 174044 195140 174050 195152
rect 174722 195140 174728 195152
rect 174044 195112 174728 195140
rect 174044 195100 174050 195112
rect 174722 195100 174728 195112
rect 174780 195100 174786 195152
rect 176562 195100 176568 195152
rect 176620 195140 176626 195152
rect 177206 195140 177212 195152
rect 176620 195112 177212 195140
rect 176620 195100 176626 195112
rect 177206 195100 177212 195112
rect 177264 195100 177270 195152
rect 155126 195032 155132 195084
rect 155184 195072 155190 195084
rect 155678 195072 155684 195084
rect 155184 195044 155684 195072
rect 155184 195032 155190 195044
rect 155678 195032 155684 195044
rect 155736 195032 155742 195084
rect 175642 195032 175648 195084
rect 175700 195072 175706 195084
rect 176378 195072 176384 195084
rect 175700 195044 176384 195072
rect 175700 195032 175706 195044
rect 176378 195032 176384 195044
rect 176436 195032 176442 195084
rect 148594 195004 148600 195016
rect 128504 194976 133874 195004
rect 142126 194976 148600 195004
rect 128504 194964 128510 194976
rect 133846 194936 133874 194976
rect 148594 194964 148600 194976
rect 148652 194964 148658 195016
rect 142890 194936 142896 194948
rect 133846 194908 142896 194936
rect 142890 194896 142896 194908
rect 142948 194896 142954 194948
rect 155954 194896 155960 194948
rect 156012 194936 156018 194948
rect 156782 194936 156788 194948
rect 156012 194908 156788 194936
rect 156012 194896 156018 194908
rect 156782 194896 156788 194908
rect 156840 194896 156846 194948
rect 165246 194896 165252 194948
rect 165304 194936 165310 194948
rect 165304 194908 176240 194936
rect 165304 194896 165310 194908
rect 167178 194828 167184 194880
rect 167236 194868 167242 194880
rect 167822 194868 167828 194880
rect 167236 194840 167828 194868
rect 167236 194828 167242 194840
rect 167822 194828 167828 194840
rect 167880 194828 167886 194880
rect 173710 194828 173716 194880
rect 173768 194868 173774 194880
rect 176102 194868 176108 194880
rect 173768 194840 176108 194868
rect 173768 194828 173774 194840
rect 176102 194828 176108 194840
rect 176160 194828 176166 194880
rect 176212 194868 176240 194908
rect 177574 194868 177580 194880
rect 176212 194840 177580 194868
rect 177574 194828 177580 194840
rect 177632 194828 177638 194880
rect 132034 194760 132040 194812
rect 132092 194800 132098 194812
rect 139210 194800 139216 194812
rect 132092 194772 139216 194800
rect 132092 194760 132098 194772
rect 139210 194760 139216 194772
rect 139268 194760 139274 194812
rect 176194 194760 176200 194812
rect 176252 194800 176258 194812
rect 180334 194800 180340 194812
rect 176252 194772 180340 194800
rect 176252 194760 176258 194772
rect 180334 194760 180340 194772
rect 180392 194760 180398 194812
rect 183830 194692 183836 194744
rect 183888 194732 183894 194744
rect 186498 194732 186504 194744
rect 183888 194704 186504 194732
rect 183888 194692 183894 194704
rect 186498 194692 186504 194704
rect 186556 194692 186562 194744
rect 174078 194556 174084 194608
rect 174136 194596 174142 194608
rect 174998 194596 175004 194608
rect 174136 194568 175004 194596
rect 174136 194556 174142 194568
rect 174998 194556 175004 194568
rect 175056 194556 175062 194608
rect 130562 194488 130568 194540
rect 130620 194528 130626 194540
rect 144914 194528 144920 194540
rect 130620 194500 144920 194528
rect 130620 194488 130626 194500
rect 144914 194488 144920 194500
rect 144972 194488 144978 194540
rect 130378 194420 130384 194472
rect 130436 194460 130442 194472
rect 146754 194460 146760 194472
rect 130436 194432 146760 194460
rect 130436 194420 130442 194432
rect 146754 194420 146760 194432
rect 146812 194420 146818 194472
rect 130930 194352 130936 194404
rect 130988 194392 130994 194404
rect 147582 194392 147588 194404
rect 130988 194364 147588 194392
rect 130988 194352 130994 194364
rect 147582 194352 147588 194364
rect 147640 194352 147646 194404
rect 156138 194352 156144 194404
rect 156196 194392 156202 194404
rect 181438 194392 181444 194404
rect 156196 194364 181444 194392
rect 156196 194352 156202 194364
rect 181438 194352 181444 194364
rect 181496 194352 181502 194404
rect 127802 194284 127808 194336
rect 127860 194324 127866 194336
rect 144638 194324 144644 194336
rect 127860 194296 144644 194324
rect 127860 194284 127866 194296
rect 144638 194284 144644 194296
rect 144696 194284 144702 194336
rect 153378 194284 153384 194336
rect 153436 194324 153442 194336
rect 181530 194324 181536 194336
rect 153436 194296 181536 194324
rect 153436 194284 153442 194296
rect 181530 194284 181536 194296
rect 181588 194284 181594 194336
rect 127986 194216 127992 194268
rect 128044 194256 128050 194268
rect 148042 194256 148048 194268
rect 128044 194228 148048 194256
rect 128044 194216 128050 194228
rect 148042 194216 148048 194228
rect 148100 194216 148106 194268
rect 176286 194216 176292 194268
rect 176344 194256 176350 194268
rect 209958 194256 209964 194268
rect 176344 194228 209964 194256
rect 176344 194216 176350 194228
rect 209958 194216 209964 194228
rect 210016 194216 210022 194268
rect 122190 194148 122196 194200
rect 122248 194188 122254 194200
rect 143534 194188 143540 194200
rect 122248 194160 143540 194188
rect 122248 194148 122254 194160
rect 143534 194148 143540 194160
rect 143592 194148 143598 194200
rect 173802 194148 173808 194200
rect 173860 194188 173866 194200
rect 207290 194188 207296 194200
rect 173860 194160 207296 194188
rect 173860 194148 173866 194160
rect 207290 194148 207296 194160
rect 207348 194148 207354 194200
rect 108482 194080 108488 194132
rect 108540 194120 108546 194132
rect 140774 194120 140780 194132
rect 108540 194092 140780 194120
rect 108540 194080 108546 194092
rect 140774 194080 140780 194092
rect 140832 194080 140838 194132
rect 170858 194080 170864 194132
rect 170916 194120 170922 194132
rect 203058 194120 203064 194132
rect 170916 194092 203064 194120
rect 170916 194080 170922 194092
rect 203058 194080 203064 194092
rect 203116 194080 203122 194132
rect 108666 194012 108672 194064
rect 108724 194052 108730 194064
rect 139118 194052 139124 194064
rect 108724 194024 139124 194052
rect 108724 194012 108730 194024
rect 139118 194012 139124 194024
rect 139176 194012 139182 194064
rect 174354 194012 174360 194064
rect 174412 194052 174418 194064
rect 208762 194052 208768 194064
rect 174412 194024 208768 194052
rect 174412 194012 174418 194024
rect 208762 194012 208768 194024
rect 208820 194012 208826 194064
rect 113910 193944 113916 193996
rect 113968 193984 113974 193996
rect 145558 193984 145564 193996
rect 113968 193956 145564 193984
rect 113968 193944 113974 193956
rect 145558 193944 145564 193956
rect 145616 193944 145622 193996
rect 153286 193944 153292 193996
rect 153344 193984 153350 193996
rect 154022 193984 154028 193996
rect 153344 193956 154028 193984
rect 153344 193944 153350 193956
rect 154022 193944 154028 193956
rect 154080 193944 154086 193996
rect 173434 193944 173440 193996
rect 173492 193984 173498 193996
rect 207566 193984 207572 193996
rect 173492 193956 207572 193984
rect 173492 193944 173498 193956
rect 207566 193944 207572 193956
rect 207624 193944 207630 193996
rect 111426 193876 111432 193928
rect 111484 193916 111490 193928
rect 145650 193916 145656 193928
rect 111484 193888 145656 193916
rect 111484 193876 111490 193888
rect 145650 193876 145656 193888
rect 145708 193876 145714 193928
rect 173618 193876 173624 193928
rect 173676 193916 173682 193928
rect 207658 193916 207664 193928
rect 173676 193888 207664 193916
rect 173676 193876 173682 193888
rect 207658 193876 207664 193888
rect 207716 193876 207722 193928
rect 111242 193808 111248 193860
rect 111300 193848 111306 193860
rect 145006 193848 145012 193860
rect 111300 193820 145012 193848
rect 111300 193808 111306 193820
rect 145006 193808 145012 193820
rect 145064 193808 145070 193860
rect 166810 193808 166816 193860
rect 166868 193848 166874 193860
rect 213086 193848 213092 193860
rect 166868 193820 213092 193848
rect 166868 193808 166874 193820
rect 213086 193808 213092 193820
rect 213144 193808 213150 193860
rect 130746 193740 130752 193792
rect 130804 193780 130810 193792
rect 147490 193780 147496 193792
rect 130804 193752 147496 193780
rect 130804 193740 130810 193752
rect 147490 193740 147496 193752
rect 147548 193740 147554 193792
rect 130562 193672 130568 193724
rect 130620 193712 130626 193724
rect 144086 193712 144092 193724
rect 130620 193684 144092 193712
rect 130620 193672 130626 193684
rect 144086 193672 144092 193684
rect 144144 193672 144150 193724
rect 174262 193672 174268 193724
rect 174320 193712 174326 193724
rect 174814 193712 174820 193724
rect 174320 193684 174820 193712
rect 174320 193672 174326 193684
rect 174814 193672 174820 193684
rect 174872 193672 174878 193724
rect 130838 193604 130844 193656
rect 130896 193644 130902 193656
rect 145098 193644 145104 193656
rect 130896 193616 145104 193644
rect 130896 193604 130902 193616
rect 145098 193604 145104 193616
rect 145156 193604 145162 193656
rect 141694 193536 141700 193588
rect 141752 193576 141758 193588
rect 143626 193576 143632 193588
rect 141752 193548 143632 193576
rect 141752 193536 141758 193548
rect 143626 193536 143632 193548
rect 143684 193536 143690 193588
rect 149698 193536 149704 193588
rect 149756 193576 149762 193588
rect 150434 193576 150440 193588
rect 149756 193548 150440 193576
rect 149756 193536 149762 193548
rect 150434 193536 150440 193548
rect 150492 193536 150498 193588
rect 150618 193128 150624 193180
rect 150676 193168 150682 193180
rect 151538 193168 151544 193180
rect 150676 193140 151544 193168
rect 150676 193128 150682 193140
rect 151538 193128 151544 193140
rect 151596 193128 151602 193180
rect 189810 193128 189816 193180
rect 189868 193168 189874 193180
rect 580166 193168 580172 193180
rect 189868 193140 580172 193168
rect 189868 193128 189874 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 107102 193060 107108 193112
rect 107160 193100 107166 193112
rect 130010 193100 130016 193112
rect 107160 193072 130016 193100
rect 107160 193060 107166 193072
rect 130010 193060 130016 193072
rect 130068 193060 130074 193112
rect 162118 193060 162124 193112
rect 162176 193100 162182 193112
rect 162670 193100 162676 193112
rect 162176 193072 162676 193100
rect 162176 193060 162182 193072
rect 162670 193060 162676 193072
rect 162728 193060 162734 193112
rect 174446 193060 174452 193112
rect 174504 193100 174510 193112
rect 175090 193100 175096 193112
rect 174504 193072 175096 193100
rect 174504 193060 174510 193072
rect 175090 193060 175096 193072
rect 175148 193060 175154 193112
rect 179414 193060 179420 193112
rect 179472 193100 179478 193112
rect 198918 193100 198924 193112
rect 179472 193072 198924 193100
rect 179472 193060 179478 193072
rect 198918 193060 198924 193072
rect 198976 193060 198982 193112
rect 105814 192992 105820 193044
rect 105872 193032 105878 193044
rect 129918 193032 129924 193044
rect 105872 193004 129924 193032
rect 105872 192992 105878 193004
rect 129918 192992 129924 193004
rect 129976 192992 129982 193044
rect 138474 192992 138480 193044
rect 138532 193032 138538 193044
rect 139302 193032 139308 193044
rect 138532 193004 139308 193032
rect 138532 192992 138538 193004
rect 139302 192992 139308 193004
rect 139360 192992 139366 193044
rect 171594 192992 171600 193044
rect 171652 193032 171658 193044
rect 204714 193032 204720 193044
rect 171652 193004 204720 193032
rect 171652 192992 171658 193004
rect 204714 192992 204720 193004
rect 204772 192992 204778 193044
rect 122466 192924 122472 192976
rect 122524 192964 122530 192976
rect 147214 192964 147220 192976
rect 122524 192936 147220 192964
rect 122524 192924 122530 192936
rect 147214 192924 147220 192936
rect 147272 192924 147278 192976
rect 157518 192924 157524 192976
rect 157576 192964 157582 192976
rect 158346 192964 158352 192976
rect 157576 192936 158352 192964
rect 157576 192924 157582 192936
rect 158346 192924 158352 192936
rect 158404 192924 158410 192976
rect 178034 192924 178040 192976
rect 178092 192964 178098 192976
rect 205910 192964 205916 192976
rect 178092 192936 205916 192964
rect 178092 192924 178098 192936
rect 205910 192924 205916 192936
rect 205968 192924 205974 192976
rect 100478 192856 100484 192908
rect 100536 192896 100542 192908
rect 128538 192896 128544 192908
rect 100536 192868 128544 192896
rect 100536 192856 100542 192868
rect 128538 192856 128544 192868
rect 128596 192856 128602 192908
rect 170766 192856 170772 192908
rect 170824 192896 170830 192908
rect 204530 192896 204536 192908
rect 170824 192868 204536 192896
rect 170824 192856 170830 192868
rect 204530 192856 204536 192868
rect 204588 192856 204594 192908
rect 110322 192788 110328 192840
rect 110380 192828 110386 192840
rect 144362 192828 144368 192840
rect 110380 192800 144368 192828
rect 110380 192788 110386 192800
rect 144362 192788 144368 192800
rect 144420 192788 144426 192840
rect 173158 192788 173164 192840
rect 173216 192828 173222 192840
rect 206002 192828 206008 192840
rect 173216 192800 206008 192828
rect 173216 192788 173222 192800
rect 206002 192788 206008 192800
rect 206060 192788 206066 192840
rect 110138 192720 110144 192772
rect 110196 192760 110202 192772
rect 144178 192760 144184 192772
rect 110196 192732 144184 192760
rect 110196 192720 110202 192732
rect 144178 192720 144184 192732
rect 144236 192720 144242 192772
rect 150526 192720 150532 192772
rect 150584 192760 150590 192772
rect 185670 192760 185676 192772
rect 150584 192732 185676 192760
rect 150584 192720 150590 192732
rect 185670 192720 185676 192732
rect 185728 192720 185734 192772
rect 123938 192652 123944 192704
rect 123996 192692 124002 192704
rect 161842 192692 161848 192704
rect 123996 192664 161848 192692
rect 123996 192652 124002 192664
rect 161842 192652 161848 192664
rect 161900 192652 161906 192704
rect 170214 192652 170220 192704
rect 170272 192692 170278 192704
rect 204898 192692 204904 192704
rect 170272 192664 204904 192692
rect 170272 192652 170278 192664
rect 204898 192652 204904 192664
rect 204956 192652 204962 192704
rect 108758 192584 108764 192636
rect 108816 192624 108822 192636
rect 143074 192624 143080 192636
rect 108816 192596 143080 192624
rect 108816 192584 108822 192596
rect 143074 192584 143080 192596
rect 143132 192584 143138 192636
rect 156874 192584 156880 192636
rect 156932 192624 156938 192636
rect 210326 192624 210332 192636
rect 156932 192596 210332 192624
rect 156932 192584 156938 192596
rect 210326 192584 210332 192596
rect 210384 192584 210390 192636
rect 104342 192516 104348 192568
rect 104400 192556 104406 192568
rect 138014 192556 138020 192568
rect 104400 192528 138020 192556
rect 104400 192516 104406 192528
rect 138014 192516 138020 192528
rect 138072 192516 138078 192568
rect 155862 192516 155868 192568
rect 155920 192556 155926 192568
rect 209774 192556 209780 192568
rect 155920 192528 209780 192556
rect 155920 192516 155926 192528
rect 209774 192516 209780 192528
rect 209832 192516 209838 192568
rect 110046 192448 110052 192500
rect 110104 192488 110110 192500
rect 143534 192488 143540 192500
rect 110104 192460 143540 192488
rect 110104 192448 110110 192460
rect 143534 192448 143540 192460
rect 143592 192448 143598 192500
rect 155218 192448 155224 192500
rect 155276 192488 155282 192500
rect 211154 192488 211160 192500
rect 155276 192460 211160 192488
rect 155276 192448 155282 192460
rect 211154 192448 211160 192460
rect 211212 192448 211218 192500
rect 161842 192380 161848 192432
rect 161900 192420 161906 192432
rect 162394 192420 162400 192432
rect 161900 192392 162400 192420
rect 161900 192380 161906 192392
rect 162394 192380 162400 192392
rect 162452 192380 162458 192432
rect 168374 192108 168380 192160
rect 168432 192148 168438 192160
rect 169662 192148 169668 192160
rect 168432 192120 169668 192148
rect 168432 192108 168438 192120
rect 169662 192108 169668 192120
rect 169720 192108 169726 192160
rect 158622 192040 158628 192092
rect 158680 192080 158686 192092
rect 160646 192080 160652 192092
rect 158680 192052 160652 192080
rect 158680 192040 158686 192052
rect 160646 192040 160652 192052
rect 160704 192040 160710 192092
rect 171318 192040 171324 192092
rect 171376 192080 171382 192092
rect 205726 192080 205732 192092
rect 171376 192052 205732 192080
rect 171376 192040 171382 192052
rect 205726 192040 205732 192052
rect 205784 192040 205790 192092
rect 170674 191972 170680 192024
rect 170732 192012 170738 192024
rect 204346 192012 204352 192024
rect 170732 191984 204352 192012
rect 170732 191972 170738 191984
rect 204346 191972 204352 191984
rect 204404 191972 204410 192024
rect 171962 191904 171968 191956
rect 172020 191944 172026 191956
rect 206094 191944 206100 191956
rect 172020 191916 206100 191944
rect 172020 191904 172026 191916
rect 206094 191904 206100 191916
rect 206152 191904 206158 191956
rect 170950 191836 170956 191888
rect 171008 191876 171014 191888
rect 204806 191876 204812 191888
rect 171008 191848 204812 191876
rect 171008 191836 171014 191848
rect 204806 191836 204812 191848
rect 204864 191836 204870 191888
rect 171318 191768 171324 191820
rect 171376 191808 171382 191820
rect 172238 191808 172244 191820
rect 171376 191780 172244 191808
rect 171376 191768 171382 191780
rect 172238 191768 172244 191780
rect 172296 191768 172302 191820
rect 132586 191700 132592 191752
rect 132644 191740 132650 191752
rect 133414 191740 133420 191752
rect 132644 191712 133420 191740
rect 132644 191700 132650 191712
rect 133414 191700 133420 191712
rect 133472 191700 133478 191752
rect 130286 191632 130292 191684
rect 130344 191672 130350 191684
rect 132494 191672 132500 191684
rect 130344 191644 132500 191672
rect 130344 191632 130350 191644
rect 132494 191632 132500 191644
rect 132552 191632 132558 191684
rect 131022 191564 131028 191616
rect 131080 191604 131086 191616
rect 135254 191604 135260 191616
rect 131080 191576 135260 191604
rect 131080 191564 131086 191576
rect 135254 191564 135260 191576
rect 135312 191564 135318 191616
rect 166258 191564 166264 191616
rect 166316 191604 166322 191616
rect 185854 191604 185860 191616
rect 166316 191576 185860 191604
rect 166316 191564 166322 191576
rect 185854 191564 185860 191576
rect 185912 191564 185918 191616
rect 132218 191496 132224 191548
rect 132276 191536 132282 191548
rect 139578 191536 139584 191548
rect 132276 191508 139584 191536
rect 132276 191496 132282 191508
rect 139578 191496 139584 191508
rect 139636 191496 139642 191548
rect 164142 191496 164148 191548
rect 164200 191536 164206 191548
rect 184198 191536 184204 191548
rect 164200 191508 184204 191536
rect 164200 191496 164206 191508
rect 184198 191496 184204 191508
rect 184256 191496 184262 191548
rect 122558 191428 122564 191480
rect 122616 191468 122622 191480
rect 141234 191468 141240 191480
rect 122616 191440 141240 191468
rect 122616 191428 122622 191440
rect 141234 191428 141240 191440
rect 141292 191428 141298 191480
rect 162670 191428 162676 191480
rect 162728 191468 162734 191480
rect 185762 191468 185768 191480
rect 162728 191440 185768 191468
rect 162728 191428 162734 191440
rect 185762 191428 185768 191440
rect 185820 191428 185826 191480
rect 123846 191360 123852 191412
rect 123904 191400 123910 191412
rect 154574 191400 154580 191412
rect 123904 191372 154580 191400
rect 123904 191360 123910 191372
rect 154574 191360 154580 191372
rect 154632 191360 154638 191412
rect 163590 191360 163596 191412
rect 163648 191400 163654 191412
rect 164142 191400 164148 191412
rect 163648 191372 164148 191400
rect 163648 191360 163654 191372
rect 164142 191360 164148 191372
rect 164200 191360 164206 191412
rect 167638 191360 167644 191412
rect 167696 191400 167702 191412
rect 201494 191400 201500 191412
rect 167696 191372 201500 191400
rect 167696 191360 167702 191372
rect 201494 191360 201500 191372
rect 201552 191360 201558 191412
rect 103330 191292 103336 191344
rect 103388 191332 103394 191344
rect 131022 191332 131028 191344
rect 103388 191304 131028 191332
rect 103388 191292 103394 191304
rect 131022 191292 131028 191304
rect 131080 191292 131086 191344
rect 167454 191292 167460 191344
rect 167512 191332 167518 191344
rect 201770 191332 201776 191344
rect 167512 191304 201776 191332
rect 167512 191292 167518 191304
rect 201770 191292 201776 191304
rect 201828 191292 201834 191344
rect 99190 191224 99196 191276
rect 99248 191264 99254 191276
rect 130286 191264 130292 191276
rect 99248 191236 130292 191264
rect 99248 191224 99254 191236
rect 130286 191224 130292 191236
rect 130344 191224 130350 191276
rect 133966 191264 133972 191276
rect 131316 191236 133972 191264
rect 100386 191156 100392 191208
rect 100444 191196 100450 191208
rect 131316 191196 131344 191236
rect 133966 191224 133972 191236
rect 134024 191224 134030 191276
rect 168650 191224 168656 191276
rect 168708 191264 168714 191276
rect 202966 191264 202972 191276
rect 168708 191236 202972 191264
rect 168708 191224 168714 191236
rect 202966 191224 202972 191236
rect 203024 191224 203030 191276
rect 100444 191168 131344 191196
rect 100444 191156 100450 191168
rect 134058 191156 134064 191208
rect 134116 191196 134122 191208
rect 134518 191196 134524 191208
rect 134116 191168 134524 191196
rect 134116 191156 134122 191168
rect 134518 191156 134524 191168
rect 134576 191156 134582 191208
rect 135714 191156 135720 191208
rect 135772 191196 135778 191208
rect 136266 191196 136272 191208
rect 135772 191168 136272 191196
rect 135772 191156 135778 191168
rect 136266 191156 136272 191168
rect 136324 191156 136330 191208
rect 137094 191156 137100 191208
rect 137152 191196 137158 191208
rect 137554 191196 137560 191208
rect 137152 191168 137560 191196
rect 137152 191156 137158 191168
rect 137554 191156 137560 191168
rect 137612 191156 137618 191208
rect 161198 191156 161204 191208
rect 161256 191196 161262 191208
rect 216766 191196 216772 191208
rect 161256 191168 216772 191196
rect 161256 191156 161262 191168
rect 216766 191156 216772 191168
rect 216824 191156 216830 191208
rect 103054 191088 103060 191140
rect 103112 191128 103118 191140
rect 143442 191128 143448 191140
rect 103112 191100 143448 191128
rect 103112 191088 103118 191100
rect 143442 191088 143448 191100
rect 143500 191088 143506 191140
rect 152182 191088 152188 191140
rect 152240 191128 152246 191140
rect 218330 191128 218336 191140
rect 152240 191100 218336 191128
rect 152240 191088 152246 191100
rect 218330 191088 218336 191100
rect 218388 191088 218394 191140
rect 134150 191020 134156 191072
rect 134208 191060 134214 191072
rect 135162 191060 135168 191072
rect 134208 191032 135168 191060
rect 134208 191020 134214 191032
rect 135162 191020 135168 191032
rect 135220 191020 135226 191072
rect 135530 191020 135536 191072
rect 135588 191060 135594 191072
rect 136450 191060 136456 191072
rect 135588 191032 136456 191060
rect 135588 191020 135594 191032
rect 136450 191020 136456 191032
rect 136508 191020 136514 191072
rect 149882 190952 149888 191004
rect 149940 190992 149946 191004
rect 150158 190992 150164 191004
rect 149940 190964 150164 190992
rect 149940 190952 149946 190964
rect 150158 190952 150164 190964
rect 150216 190952 150222 191004
rect 121822 190408 121828 190460
rect 121880 190448 121886 190460
rect 149974 190448 149980 190460
rect 121880 190420 149980 190448
rect 121880 190408 121886 190420
rect 149974 190408 149980 190420
rect 150032 190408 150038 190460
rect 177206 190408 177212 190460
rect 177264 190448 177270 190460
rect 210418 190448 210424 190460
rect 177264 190420 210424 190448
rect 177264 190408 177270 190420
rect 210418 190408 210424 190420
rect 210476 190408 210482 190460
rect 107378 190340 107384 190392
rect 107436 190380 107442 190392
rect 138658 190380 138664 190392
rect 107436 190352 138664 190380
rect 107436 190340 107442 190352
rect 138658 190340 138664 190352
rect 138716 190340 138722 190392
rect 177298 190340 177304 190392
rect 177356 190380 177362 190392
rect 211706 190380 211712 190392
rect 177356 190352 211712 190380
rect 177356 190340 177362 190352
rect 211706 190340 211712 190352
rect 211764 190340 211770 190392
rect 106182 190272 106188 190324
rect 106240 190312 106246 190324
rect 130286 190312 130292 190324
rect 106240 190284 130292 190312
rect 106240 190272 106246 190284
rect 130286 190272 130292 190284
rect 130344 190272 130350 190324
rect 130654 190272 130660 190324
rect 130712 190312 130718 190324
rect 130930 190312 130936 190324
rect 130712 190284 130936 190312
rect 130712 190272 130718 190284
rect 130930 190272 130936 190284
rect 130988 190272 130994 190324
rect 175550 190272 175556 190324
rect 175608 190312 175614 190324
rect 210050 190312 210056 190324
rect 175608 190284 210056 190312
rect 175608 190272 175614 190284
rect 210050 190272 210056 190284
rect 210108 190272 210114 190324
rect 104250 190204 104256 190256
rect 104308 190244 104314 190256
rect 136358 190244 136364 190256
rect 104308 190216 136364 190244
rect 104308 190204 104314 190216
rect 136358 190204 136364 190216
rect 136416 190204 136422 190256
rect 172882 190204 172888 190256
rect 172940 190244 172946 190256
rect 207474 190244 207480 190256
rect 172940 190216 207480 190244
rect 172940 190204 172946 190216
rect 207474 190204 207480 190216
rect 207532 190204 207538 190256
rect 100570 190136 100576 190188
rect 100628 190176 100634 190188
rect 132310 190176 132316 190188
rect 100628 190148 132316 190176
rect 100628 190136 100634 190148
rect 132310 190136 132316 190148
rect 132368 190136 132374 190188
rect 160554 190136 160560 190188
rect 160612 190176 160618 190188
rect 195146 190176 195152 190188
rect 160612 190148 195152 190176
rect 160612 190136 160618 190148
rect 195146 190136 195152 190148
rect 195204 190136 195210 190188
rect 103422 190068 103428 190120
rect 103480 190108 103486 190120
rect 135622 190108 135628 190120
rect 103480 190080 135628 190108
rect 103480 190068 103486 190080
rect 135622 190068 135628 190080
rect 135680 190068 135686 190120
rect 174262 190068 174268 190120
rect 174320 190108 174326 190120
rect 208946 190108 208952 190120
rect 174320 190080 208952 190108
rect 174320 190068 174326 190080
rect 208946 190068 208952 190080
rect 209004 190068 209010 190120
rect 111610 190000 111616 190052
rect 111668 190040 111674 190052
rect 144730 190040 144736 190052
rect 111668 190012 144736 190040
rect 111668 190000 111674 190012
rect 144730 190000 144736 190012
rect 144788 190000 144794 190052
rect 164694 190000 164700 190052
rect 164752 190040 164758 190052
rect 205818 190040 205824 190052
rect 164752 190012 205824 190040
rect 164752 190000 164758 190012
rect 205818 190000 205824 190012
rect 205876 190000 205882 190052
rect 104618 189932 104624 189984
rect 104676 189972 104682 189984
rect 104676 189944 130240 189972
rect 104676 189932 104682 189944
rect 102870 189864 102876 189916
rect 102928 189904 102934 189916
rect 130102 189904 130108 189916
rect 102928 189876 130108 189904
rect 102928 189864 102934 189876
rect 130102 189864 130108 189876
rect 130160 189864 130166 189916
rect 130212 189904 130240 189944
rect 130286 189932 130292 189984
rect 130344 189972 130350 189984
rect 137738 189972 137744 189984
rect 130344 189944 137744 189972
rect 130344 189932 130350 189944
rect 137738 189932 137744 189944
rect 137796 189932 137802 189984
rect 163498 189932 163504 189984
rect 163556 189972 163562 189984
rect 214282 189972 214288 189984
rect 163556 189944 214288 189972
rect 163556 189932 163562 189944
rect 214282 189932 214288 189944
rect 214340 189932 214346 189984
rect 137278 189904 137284 189916
rect 130212 189876 137284 189904
rect 137278 189864 137284 189876
rect 137336 189864 137342 189916
rect 159174 189864 159180 189916
rect 159232 189904 159238 189916
rect 216950 189904 216956 189916
rect 159232 189876 216956 189904
rect 159232 189864 159238 189876
rect 216950 189864 216956 189876
rect 217008 189864 217014 189916
rect 102962 189796 102968 189848
rect 103020 189836 103026 189848
rect 136910 189836 136916 189848
rect 103020 189808 136916 189836
rect 103020 189796 103026 189808
rect 136910 189796 136916 189808
rect 136968 189796 136974 189848
rect 155402 189796 155408 189848
rect 155460 189836 155466 189848
rect 218238 189836 218244 189848
rect 155460 189808 218244 189836
rect 155460 189796 155466 189808
rect 218238 189796 218244 189808
rect 218296 189796 218302 189848
rect 101582 189728 101588 189780
rect 101640 189768 101646 189780
rect 136082 189768 136088 189780
rect 101640 189740 136088 189768
rect 101640 189728 101646 189740
rect 136082 189728 136088 189740
rect 136140 189728 136146 189780
rect 154390 189728 154396 189780
rect 154448 189768 154454 189780
rect 218422 189768 218428 189780
rect 154448 189740 218428 189768
rect 154448 189728 154454 189740
rect 218422 189728 218428 189740
rect 218480 189728 218486 189780
rect 130102 189660 130108 189712
rect 130160 189700 130166 189712
rect 137462 189700 137468 189712
rect 130160 189672 137468 189700
rect 130160 189660 130166 189672
rect 137462 189660 137468 189672
rect 137520 189660 137526 189712
rect 174446 189660 174452 189712
rect 174504 189700 174510 189712
rect 207382 189700 207388 189712
rect 174504 189672 207388 189700
rect 174504 189660 174510 189672
rect 207382 189660 207388 189672
rect 207440 189660 207446 189712
rect 156322 189592 156328 189644
rect 156380 189632 156386 189644
rect 187418 189632 187424 189644
rect 156380 189604 187424 189632
rect 156380 189592 156386 189604
rect 187418 189592 187424 189604
rect 187476 189592 187482 189644
rect 160462 189524 160468 189576
rect 160520 189564 160526 189576
rect 185578 189564 185584 189576
rect 160520 189536 185584 189564
rect 160520 189524 160526 189536
rect 185578 189524 185584 189536
rect 185636 189524 185642 189576
rect 3418 188980 3424 189032
rect 3476 189020 3482 189032
rect 117774 189020 117780 189032
rect 3476 188992 117780 189020
rect 3476 188980 3482 188992
rect 117774 188980 117780 188992
rect 117832 188980 117838 189032
rect 166074 187552 166080 187604
rect 166132 187592 166138 187604
rect 200390 187592 200396 187604
rect 166132 187564 200396 187592
rect 166132 187552 166138 187564
rect 200390 187552 200396 187564
rect 200448 187552 200454 187604
rect 161842 187484 161848 187536
rect 161900 187524 161906 187536
rect 209038 187524 209044 187536
rect 161900 187496 209044 187524
rect 161900 187484 161906 187496
rect 209038 187484 209044 187496
rect 209096 187484 209102 187536
rect 160002 187416 160008 187468
rect 160060 187456 160066 187468
rect 207014 187456 207020 187468
rect 160060 187428 207020 187456
rect 160060 187416 160066 187428
rect 207014 187416 207020 187428
rect 207072 187416 207078 187468
rect 159082 187348 159088 187400
rect 159140 187388 159146 187400
rect 207106 187388 207112 187400
rect 159140 187360 207112 187388
rect 159140 187348 159146 187360
rect 207106 187348 207112 187360
rect 207164 187348 207170 187400
rect 161934 187280 161940 187332
rect 161992 187320 161998 187332
rect 210142 187320 210148 187332
rect 161992 187292 210148 187320
rect 161992 187280 161998 187292
rect 210142 187280 210148 187292
rect 210200 187280 210206 187332
rect 101490 187212 101496 187264
rect 101548 187252 101554 187264
rect 134978 187252 134984 187264
rect 101548 187224 134984 187252
rect 101548 187212 101554 187224
rect 134978 187212 134984 187224
rect 135036 187212 135042 187264
rect 154758 187212 154764 187264
rect 154816 187252 154822 187264
rect 214190 187252 214196 187264
rect 154816 187224 214196 187252
rect 154816 187212 154822 187224
rect 214190 187212 214196 187224
rect 214248 187212 214254 187264
rect 99098 187144 99104 187196
rect 99156 187184 99162 187196
rect 133598 187184 133604 187196
rect 99156 187156 133604 187184
rect 99156 187144 99162 187156
rect 133598 187144 133604 187156
rect 133656 187144 133662 187196
rect 152826 187144 152832 187196
rect 152884 187184 152890 187196
rect 214098 187184 214104 187196
rect 152884 187156 214104 187184
rect 152884 187144 152890 187156
rect 214098 187144 214104 187156
rect 214156 187144 214162 187196
rect 99282 187076 99288 187128
rect 99340 187116 99346 187128
rect 132770 187116 132776 187128
rect 99340 187088 132776 187116
rect 99340 187076 99346 187088
rect 132770 187076 132776 187088
rect 132828 187076 132834 187128
rect 149330 187076 149336 187128
rect 149388 187116 149394 187128
rect 211614 187116 211620 187128
rect 149388 187088 211620 187116
rect 149388 187076 149394 187088
rect 211614 187076 211620 187088
rect 211672 187076 211678 187128
rect 99006 187008 99012 187060
rect 99064 187048 99070 187060
rect 133230 187048 133236 187060
rect 99064 187020 133236 187048
rect 99064 187008 99070 187020
rect 133230 187008 133236 187020
rect 133288 187008 133294 187060
rect 151078 187008 151084 187060
rect 151136 187048 151142 187060
rect 215754 187048 215760 187060
rect 151136 187020 215760 187048
rect 151136 187008 151142 187020
rect 215754 187008 215760 187020
rect 215812 187008 215818 187060
rect 100202 186940 100208 186992
rect 100260 186980 100266 186992
rect 134334 186980 134340 186992
rect 100260 186952 134340 186980
rect 100260 186940 100266 186952
rect 134334 186940 134340 186952
rect 134392 186940 134398 186992
rect 150802 186940 150808 186992
rect 150860 186980 150866 186992
rect 218514 186980 218520 186992
rect 150860 186952 218520 186980
rect 150860 186940 150866 186952
rect 218514 186940 218520 186952
rect 218572 186940 218578 186992
rect 188522 178032 188528 178084
rect 188580 178072 188586 178084
rect 580166 178072 580172 178084
rect 188580 178044 580172 178072
rect 188580 178032 188586 178044
rect 580166 178032 580172 178044
rect 580224 178032 580230 178084
rect 189810 165588 189816 165640
rect 189868 165628 189874 165640
rect 580166 165628 580172 165640
rect 189868 165600 580172 165628
rect 189868 165588 189874 165600
rect 580166 165588 580172 165600
rect 580224 165588 580230 165640
rect 168742 158380 168748 158432
rect 168800 158420 168806 158432
rect 189718 158420 189724 158432
rect 168800 158392 189724 158420
rect 168800 158380 168806 158392
rect 189718 158380 189724 158392
rect 189776 158380 189782 158432
rect 172882 158312 172888 158364
rect 172940 158352 172946 158364
rect 201954 158352 201960 158364
rect 172940 158324 201960 158352
rect 172940 158312 172946 158324
rect 201954 158312 201960 158324
rect 202012 158312 202018 158364
rect 170030 158244 170036 158296
rect 170088 158284 170094 158296
rect 203242 158284 203248 158296
rect 170088 158256 203248 158284
rect 170088 158244 170094 158256
rect 203242 158244 203248 158256
rect 203300 158244 203306 158296
rect 166074 158176 166080 158228
rect 166132 158216 166138 158228
rect 203150 158216 203156 158228
rect 166132 158188 203156 158216
rect 166132 158176 166138 158188
rect 203150 158176 203156 158188
rect 203208 158176 203214 158228
rect 159726 158108 159732 158160
rect 159784 158148 159790 158160
rect 214466 158148 214472 158160
rect 159784 158120 214472 158148
rect 159784 158108 159790 158120
rect 214466 158108 214472 158120
rect 214524 158108 214530 158160
rect 152090 158040 152096 158092
rect 152148 158080 152154 158092
rect 213178 158080 213184 158092
rect 152148 158052 213184 158080
rect 152148 158040 152154 158052
rect 213178 158040 213184 158052
rect 213236 158040 213242 158092
rect 152182 157972 152188 158024
rect 152240 158012 152246 158024
rect 217134 158012 217140 158024
rect 152240 157984 217140 158012
rect 152240 157972 152246 157984
rect 217134 157972 217140 157984
rect 217192 157972 217198 158024
rect 171502 155864 171508 155916
rect 171560 155904 171566 155916
rect 201862 155904 201868 155916
rect 171560 155876 201868 155904
rect 171560 155864 171566 155876
rect 201862 155864 201868 155876
rect 201920 155864 201926 155916
rect 170214 155796 170220 155848
rect 170272 155836 170278 155848
rect 191006 155836 191012 155848
rect 170272 155808 191012 155836
rect 170272 155796 170278 155808
rect 191006 155796 191012 155808
rect 191064 155796 191070 155848
rect 167270 155728 167276 155780
rect 167328 155768 167334 155780
rect 201862 155768 201868 155780
rect 167328 155740 201868 155768
rect 167328 155728 167334 155740
rect 201862 155728 201868 155740
rect 201920 155728 201926 155780
rect 167546 155660 167552 155712
rect 167604 155700 167610 155712
rect 202230 155700 202236 155712
rect 167604 155672 202236 155700
rect 167604 155660 167610 155672
rect 202230 155660 202236 155672
rect 202288 155660 202294 155712
rect 165982 155592 165988 155644
rect 166040 155632 166046 155644
rect 200758 155632 200764 155644
rect 166040 155604 200764 155632
rect 166040 155592 166046 155604
rect 200758 155592 200764 155604
rect 200816 155592 200822 155644
rect 165890 155524 165896 155576
rect 165948 155564 165954 155576
rect 200666 155564 200672 155576
rect 165948 155536 200672 155564
rect 165948 155524 165954 155536
rect 200666 155524 200672 155536
rect 200724 155524 200730 155576
rect 167362 155456 167368 155508
rect 167420 155496 167426 155508
rect 202138 155496 202144 155508
rect 167420 155468 202144 155496
rect 167420 155456 167426 155468
rect 202138 155456 202144 155468
rect 202196 155456 202202 155508
rect 177022 155388 177028 155440
rect 177080 155428 177086 155440
rect 211890 155428 211896 155440
rect 177080 155400 211896 155428
rect 177080 155388 177086 155400
rect 211890 155388 211896 155400
rect 211948 155388 211954 155440
rect 168558 155320 168564 155372
rect 168616 155360 168622 155372
rect 203426 155360 203432 155372
rect 168616 155332 203432 155360
rect 168616 155320 168622 155332
rect 203426 155320 203432 155332
rect 203484 155320 203490 155372
rect 168650 155252 168656 155304
rect 168708 155292 168714 155304
rect 203518 155292 203524 155304
rect 168708 155264 203524 155292
rect 168708 155252 168714 155264
rect 203518 155252 203524 155264
rect 203576 155252 203582 155304
rect 168282 155184 168288 155236
rect 168340 155224 168346 155236
rect 202322 155224 202328 155236
rect 168340 155196 202328 155224
rect 168340 155184 168346 155196
rect 202322 155184 202328 155196
rect 202380 155184 202386 155236
rect 174262 155116 174268 155168
rect 174320 155156 174326 155168
rect 193858 155156 193864 155168
rect 174320 155128 193864 155156
rect 174320 155116 174326 155128
rect 193858 155116 193864 155128
rect 193916 155116 193922 155168
rect 183554 154504 183560 154556
rect 183612 154544 183618 154556
rect 184290 154544 184296 154556
rect 183612 154516 184296 154544
rect 183612 154504 183618 154516
rect 184290 154504 184296 154516
rect 184348 154504 184354 154556
rect 112438 154368 112444 154420
rect 112496 154408 112502 154420
rect 132678 154408 132684 154420
rect 112496 154380 132684 154408
rect 112496 154368 112502 154380
rect 132678 154368 132684 154380
rect 132736 154368 132742 154420
rect 116578 154300 116584 154352
rect 116636 154340 116642 154352
rect 143534 154340 143540 154352
rect 116636 154312 143540 154340
rect 116636 154300 116642 154312
rect 143534 154300 143540 154312
rect 143592 154300 143598 154352
rect 113726 154232 113732 154284
rect 113784 154272 113790 154284
rect 141234 154272 141240 154284
rect 113784 154244 141240 154272
rect 113784 154232 113790 154244
rect 141234 154232 141240 154244
rect 141292 154232 141298 154284
rect 115106 154164 115112 154216
rect 115164 154204 115170 154216
rect 146386 154204 146392 154216
rect 115164 154176 146392 154204
rect 115164 154164 115170 154176
rect 146386 154164 146392 154176
rect 146444 154164 146450 154216
rect 101214 154096 101220 154148
rect 101272 154136 101278 154148
rect 134150 154136 134156 154148
rect 101272 154108 134156 154136
rect 101272 154096 101278 154108
rect 134150 154096 134156 154108
rect 134208 154096 134214 154148
rect 98914 154028 98920 154080
rect 98972 154068 98978 154080
rect 133322 154068 133328 154080
rect 98972 154040 133328 154068
rect 98972 154028 98978 154040
rect 133322 154028 133328 154040
rect 133380 154028 133386 154080
rect 100018 153960 100024 154012
rect 100076 154000 100082 154012
rect 134334 154000 134340 154012
rect 100076 153972 134340 154000
rect 100076 153960 100082 153972
rect 134334 153960 134340 153972
rect 134392 153960 134398 154012
rect 100110 153892 100116 153944
rect 100168 153932 100174 153944
rect 134426 153932 134432 153944
rect 100168 153904 134432 153932
rect 100168 153892 100174 153904
rect 134426 153892 134432 153904
rect 134484 153892 134490 153944
rect 99926 153824 99932 153876
rect 99984 153864 99990 153876
rect 134058 153864 134064 153876
rect 99984 153836 134064 153864
rect 99984 153824 99990 153836
rect 134058 153824 134064 153836
rect 134116 153824 134122 153876
rect 97258 153212 97264 153264
rect 97316 153252 97322 153264
rect 183554 153252 183560 153264
rect 97316 153224 183560 153252
rect 97316 153212 97322 153224
rect 183554 153212 183560 153224
rect 183612 153212 183618 153264
rect 160370 153144 160376 153196
rect 160428 153184 160434 153196
rect 184658 153184 184664 153196
rect 160428 153156 184664 153184
rect 160428 153144 160434 153156
rect 184658 153144 184664 153156
rect 184716 153144 184722 153196
rect 161658 153076 161664 153128
rect 161716 153116 161722 153128
rect 185946 153116 185952 153128
rect 161716 153088 185952 153116
rect 161716 153076 161722 153088
rect 185946 153076 185952 153088
rect 186004 153076 186010 153128
rect 161750 153008 161756 153060
rect 161808 153048 161814 153060
rect 186130 153048 186136 153060
rect 161808 153020 186136 153048
rect 161808 153008 161814 153020
rect 186130 153008 186136 153020
rect 186188 153008 186194 153060
rect 158898 152940 158904 152992
rect 158956 152980 158962 152992
rect 184566 152980 184572 152992
rect 158956 152952 184572 152980
rect 158956 152940 158962 152952
rect 184566 152940 184572 152952
rect 184624 152940 184630 152992
rect 158990 152872 158996 152924
rect 159048 152912 159054 152924
rect 185486 152912 185492 152924
rect 159048 152884 185492 152912
rect 159048 152872 159054 152884
rect 185486 152872 185492 152884
rect 185544 152872 185550 152924
rect 157794 152804 157800 152856
rect 157852 152844 157858 152856
rect 184382 152844 184388 152856
rect 157852 152816 184388 152844
rect 157852 152804 157858 152816
rect 184382 152804 184388 152816
rect 184440 152804 184446 152856
rect 157702 152736 157708 152788
rect 157760 152776 157766 152788
rect 184474 152776 184480 152788
rect 157760 152748 184480 152776
rect 157760 152736 157766 152748
rect 184474 152736 184480 152748
rect 184532 152736 184538 152788
rect 178954 152668 178960 152720
rect 179012 152708 179018 152720
rect 210510 152708 210516 152720
rect 179012 152680 210516 152708
rect 179012 152668 179018 152680
rect 210510 152668 210516 152680
rect 210568 152668 210574 152720
rect 176838 152600 176844 152652
rect 176896 152640 176902 152652
rect 210602 152640 210608 152652
rect 176896 152612 210608 152640
rect 176896 152600 176902 152612
rect 210602 152600 210608 152612
rect 210660 152600 210666 152652
rect 166902 152532 166908 152584
rect 166960 152572 166966 152584
rect 200574 152572 200580 152584
rect 166960 152544 200580 152572
rect 166960 152532 166966 152544
rect 200574 152532 200580 152544
rect 200632 152532 200638 152584
rect 176930 152464 176936 152516
rect 176988 152504 176994 152516
rect 211982 152504 211988 152516
rect 176988 152476 211988 152504
rect 176988 152464 176994 152476
rect 211982 152464 211988 152476
rect 212040 152464 212046 152516
rect 165706 152396 165712 152448
rect 165764 152436 165770 152448
rect 186222 152436 186228 152448
rect 165764 152408 186228 152436
rect 165764 152396 165770 152408
rect 186222 152396 186228 152408
rect 186280 152396 186286 152448
rect 165246 152328 165252 152380
rect 165304 152368 165310 152380
rect 184290 152368 184296 152380
rect 165304 152340 184296 152368
rect 165304 152328 165310 152340
rect 184290 152328 184296 152340
rect 184348 152328 184354 152380
rect 188430 151784 188436 151836
rect 188488 151824 188494 151836
rect 579982 151824 579988 151836
rect 188488 151796 579988 151824
rect 188488 151784 188494 151796
rect 579982 151784 579988 151796
rect 580040 151784 580046 151836
rect 115106 151648 115112 151700
rect 115164 151688 115170 151700
rect 141142 151688 141148 151700
rect 115164 151660 141148 151688
rect 115164 151648 115170 151660
rect 141142 151648 141148 151660
rect 141200 151648 141206 151700
rect 113542 151580 113548 151632
rect 113600 151620 113606 151632
rect 142982 151620 142988 151632
rect 113600 151592 142988 151620
rect 113600 151580 113606 151592
rect 142982 151580 142988 151592
rect 143040 151580 143046 151632
rect 168466 151580 168472 151632
rect 168524 151620 168530 151632
rect 186774 151620 186780 151632
rect 168524 151592 186780 151620
rect 168524 151580 168530 151592
rect 186774 151580 186780 151592
rect 186832 151580 186838 151632
rect 111978 151512 111984 151564
rect 112036 151552 112042 151564
rect 142430 151552 142436 151564
rect 112036 151524 142436 151552
rect 112036 151512 112042 151524
rect 142430 151512 142436 151524
rect 142488 151512 142494 151564
rect 157610 151512 157616 151564
rect 157668 151552 157674 151564
rect 188706 151552 188712 151564
rect 157668 151524 188712 151552
rect 157668 151512 157674 151524
rect 188706 151512 188712 151524
rect 188764 151512 188770 151564
rect 106826 151444 106832 151496
rect 106884 151484 106890 151496
rect 138198 151484 138204 151496
rect 106884 151456 138204 151484
rect 106884 151444 106890 151456
rect 138198 151444 138204 151456
rect 138256 151444 138262 151496
rect 156230 151444 156236 151496
rect 156288 151484 156294 151496
rect 187234 151484 187240 151496
rect 156288 151456 187240 151484
rect 156288 151444 156294 151456
rect 187234 151444 187240 151456
rect 187292 151444 187298 151496
rect 109586 151376 109592 151428
rect 109644 151416 109650 151428
rect 140958 151416 140964 151428
rect 109644 151388 140964 151416
rect 109644 151376 109650 151388
rect 140958 151376 140964 151388
rect 141016 151376 141022 151428
rect 162762 151376 162768 151428
rect 162820 151416 162826 151428
rect 198458 151416 198464 151428
rect 162820 151388 198464 151416
rect 162820 151376 162826 151388
rect 198458 151376 198464 151388
rect 198516 151376 198522 151428
rect 104158 151308 104164 151360
rect 104216 151348 104222 151360
rect 137186 151348 137192 151360
rect 104216 151320 137192 151348
rect 104216 151308 104222 151320
rect 137186 151308 137192 151320
rect 137244 151308 137250 151360
rect 163314 151308 163320 151360
rect 163372 151348 163378 151360
rect 204990 151348 204996 151360
rect 163372 151320 204996 151348
rect 163372 151308 163378 151320
rect 204990 151308 204996 151320
rect 205048 151308 205054 151360
rect 99834 151240 99840 151292
rect 99892 151280 99898 151292
rect 132586 151280 132592 151292
rect 99892 151252 132592 151280
rect 99892 151240 99898 151252
rect 132586 151240 132592 151252
rect 132644 151240 132650 151292
rect 163406 151240 163412 151292
rect 163464 151280 163470 151292
rect 207842 151280 207848 151292
rect 163464 151252 207848 151280
rect 163464 151240 163470 151252
rect 207842 151240 207848 151252
rect 207900 151240 207906 151292
rect 106734 151172 106740 151224
rect 106792 151212 106798 151224
rect 139670 151212 139676 151224
rect 106792 151184 139676 151212
rect 106792 151172 106798 151184
rect 139670 151172 139676 151184
rect 139728 151172 139734 151224
rect 154758 151172 154764 151224
rect 154816 151212 154822 151224
rect 204438 151212 204444 151224
rect 154816 151184 204444 151212
rect 154816 151172 154822 151184
rect 204438 151172 204444 151184
rect 204496 151172 204502 151224
rect 102594 151104 102600 151156
rect 102652 151144 102658 151156
rect 135530 151144 135536 151156
rect 102652 151116 135536 151144
rect 102652 151104 102658 151116
rect 135530 151104 135536 151116
rect 135588 151104 135594 151156
rect 150618 151104 150624 151156
rect 150676 151144 150682 151156
rect 209130 151144 209136 151156
rect 150676 151116 209136 151144
rect 150676 151104 150682 151116
rect 209130 151104 209136 151116
rect 209188 151104 209194 151156
rect 104066 151036 104072 151088
rect 104124 151076 104130 151088
rect 138290 151076 138296 151088
rect 104124 151048 138296 151076
rect 104124 151036 104130 151048
rect 138290 151036 138296 151048
rect 138348 151036 138354 151088
rect 154666 151036 154672 151088
rect 154724 151076 154730 151088
rect 217226 151076 217232 151088
rect 154724 151048 217232 151076
rect 154724 151036 154730 151048
rect 217226 151036 217232 151048
rect 217284 151036 217290 151088
rect 124766 150424 124772 150476
rect 124824 150464 124830 150476
rect 125134 150464 125140 150476
rect 124824 150436 125140 150464
rect 124824 150424 124830 150436
rect 125134 150424 125140 150436
rect 125192 150464 125198 150476
rect 580442 150464 580448 150476
rect 125192 150436 580448 150464
rect 125192 150424 125198 150436
rect 580442 150424 580448 150436
rect 580500 150424 580506 150476
rect 176746 150356 176752 150408
rect 176804 150396 176810 150408
rect 207750 150396 207756 150408
rect 176804 150368 207756 150396
rect 176804 150356 176810 150368
rect 207750 150356 207756 150368
rect 207808 150356 207814 150408
rect 182082 150016 182088 150068
rect 182140 150056 182146 150068
rect 197998 150056 198004 150068
rect 182140 150028 198004 150056
rect 182140 150016 182146 150028
rect 197998 150016 198004 150028
rect 198056 150016 198062 150068
rect 172790 149948 172796 150000
rect 172848 149988 172854 150000
rect 203794 149988 203800 150000
rect 172848 149960 203800 149988
rect 172848 149948 172854 149960
rect 203794 149948 203800 149960
rect 203852 149948 203858 150000
rect 175366 149880 175372 149932
rect 175424 149920 175430 149932
rect 206462 149920 206468 149932
rect 175424 149892 206468 149920
rect 175424 149880 175430 149892
rect 206462 149880 206468 149892
rect 206520 149880 206526 149932
rect 112162 149812 112168 149864
rect 112220 149852 112226 149864
rect 141786 149852 141792 149864
rect 112220 149824 141792 149852
rect 112220 149812 112226 149824
rect 141786 149812 141792 149824
rect 141844 149812 141850 149864
rect 174078 149812 174084 149864
rect 174136 149852 174142 149864
rect 206278 149852 206284 149864
rect 174136 149824 206284 149852
rect 174136 149812 174142 149824
rect 206278 149812 206284 149824
rect 206336 149812 206342 149864
rect 102686 149744 102692 149796
rect 102744 149784 102750 149796
rect 135806 149784 135812 149796
rect 102744 149756 135812 149784
rect 102744 149744 102750 149756
rect 135806 149744 135812 149756
rect 135864 149744 135870 149796
rect 173986 149744 173992 149796
rect 174044 149784 174050 149796
rect 206370 149784 206376 149796
rect 174044 149756 206376 149784
rect 174044 149744 174050 149756
rect 206370 149744 206376 149756
rect 206428 149744 206434 149796
rect 101306 149676 101312 149728
rect 101364 149716 101370 149728
rect 135898 149716 135904 149728
rect 101364 149688 135904 149716
rect 101364 149676 101370 149688
rect 135898 149676 135904 149688
rect 135956 149676 135962 149728
rect 172698 149676 172704 149728
rect 172756 149716 172762 149728
rect 205082 149716 205088 149728
rect 172756 149688 205088 149716
rect 172756 149676 172762 149688
rect 205082 149676 205088 149688
rect 205140 149676 205146 149728
rect 3142 149132 3148 149184
rect 3200 149172 3206 149184
rect 180886 149172 180892 149184
rect 3200 149144 180892 149172
rect 3200 149132 3206 149144
rect 180886 149132 180892 149144
rect 180944 149172 180950 149184
rect 182082 149172 182088 149184
rect 180944 149144 182088 149172
rect 180944 149132 180950 149144
rect 182082 149132 182088 149144
rect 182140 149132 182146 149184
rect 119246 149064 119252 149116
rect 119304 149104 119310 149116
rect 119982 149104 119988 149116
rect 119304 149076 119988 149104
rect 119304 149064 119310 149076
rect 119982 149064 119988 149076
rect 120040 149104 120046 149116
rect 580258 149104 580264 149116
rect 120040 149076 580264 149104
rect 120040 149064 120046 149076
rect 580258 149064 580264 149076
rect 580316 149064 580322 149116
rect 122558 148996 122564 149048
rect 122616 149036 122622 149048
rect 149790 149036 149796 149048
rect 122616 149008 149796 149036
rect 122616 148996 122622 149008
rect 149790 148996 149796 149008
rect 149848 148996 149854 149048
rect 160278 148996 160284 149048
rect 160336 149036 160342 149048
rect 186958 149036 186964 149048
rect 160336 149008 186964 149036
rect 160336 148996 160342 149008
rect 186958 148996 186964 149008
rect 187016 148996 187022 149048
rect 203610 148996 203616 149048
rect 203668 149036 203674 149048
rect 203794 149036 203800 149048
rect 203668 149008 203800 149036
rect 203668 148996 203674 149008
rect 203794 148996 203800 149008
rect 203852 148996 203858 149048
rect 113818 148928 113824 148980
rect 113876 148968 113882 148980
rect 125134 148968 125140 148980
rect 113876 148940 125140 148968
rect 113876 148928 113882 148940
rect 125134 148928 125140 148940
rect 125192 148928 125198 148980
rect 158806 148928 158812 148980
rect 158864 148968 158870 148980
rect 188614 148968 188620 148980
rect 158864 148940 188620 148968
rect 158864 148928 158870 148940
rect 188614 148928 188620 148940
rect 188672 148928 188678 148980
rect 115198 148860 115204 148912
rect 115256 148900 115262 148912
rect 128354 148900 128360 148912
rect 115256 148872 128360 148900
rect 115256 148860 115262 148872
rect 128354 148860 128360 148872
rect 128412 148860 128418 148912
rect 157518 148860 157524 148912
rect 157576 148900 157582 148912
rect 188154 148900 188160 148912
rect 157576 148872 188160 148900
rect 157576 148860 157582 148872
rect 188154 148860 188160 148872
rect 188212 148860 188218 148912
rect 116946 148792 116952 148844
rect 117004 148832 117010 148844
rect 142522 148832 142528 148844
rect 117004 148804 142528 148832
rect 117004 148792 117010 148804
rect 142522 148792 142528 148804
rect 142580 148792 142586 148844
rect 161566 148792 161572 148844
rect 161624 148832 161630 148844
rect 194778 148832 194784 148844
rect 161624 148804 194784 148832
rect 161624 148792 161630 148804
rect 194778 148792 194784 148804
rect 194836 148792 194842 148844
rect 122098 148724 122104 148776
rect 122156 148764 122162 148776
rect 149698 148764 149704 148776
rect 122156 148736 149704 148764
rect 122156 148724 122162 148736
rect 149698 148724 149704 148736
rect 149756 148724 149762 148776
rect 163222 148724 163228 148776
rect 163280 148764 163286 148776
rect 198366 148764 198372 148776
rect 163280 148736 198372 148764
rect 163280 148724 163286 148736
rect 198366 148724 198372 148736
rect 198424 148724 198430 148776
rect 112070 148656 112076 148708
rect 112128 148696 112134 148708
rect 142706 148696 142712 148708
rect 112128 148668 142712 148696
rect 112128 148656 112134 148668
rect 142706 148656 142712 148668
rect 142764 148656 142770 148708
rect 163130 148656 163136 148708
rect 163188 148696 163194 148708
rect 198274 148696 198280 148708
rect 163188 148668 198280 148696
rect 163188 148656 163194 148668
rect 198274 148656 198280 148668
rect 198332 148656 198338 148708
rect 114922 148588 114928 148640
rect 114980 148628 114986 148640
rect 145466 148628 145472 148640
rect 114980 148600 145472 148628
rect 114980 148588 114986 148600
rect 145466 148588 145472 148600
rect 145524 148588 145530 148640
rect 164602 148588 164608 148640
rect 164660 148628 164666 148640
rect 199838 148628 199844 148640
rect 164660 148600 199844 148628
rect 164660 148588 164666 148600
rect 199838 148588 199844 148600
rect 199896 148588 199902 148640
rect 115566 148520 115572 148572
rect 115624 148560 115630 148572
rect 145558 148560 145564 148572
rect 115624 148532 145564 148560
rect 115624 148520 115630 148532
rect 145558 148520 145564 148532
rect 145616 148520 145622 148572
rect 157150 148520 157156 148572
rect 157208 148560 157214 148572
rect 191006 148560 191012 148572
rect 157208 148532 191012 148560
rect 157208 148520 157214 148532
rect 191006 148520 191012 148532
rect 191064 148520 191070 148572
rect 116302 148452 116308 148504
rect 116360 148492 116366 148504
rect 146662 148492 146668 148504
rect 116360 148464 146668 148492
rect 116360 148452 116366 148464
rect 146662 148452 146668 148464
rect 146720 148452 146726 148504
rect 164418 148452 164424 148504
rect 164476 148492 164482 148504
rect 199378 148492 199384 148504
rect 164476 148464 199384 148492
rect 164476 148452 164482 148464
rect 199378 148452 199384 148464
rect 199436 148452 199442 148504
rect 112530 148384 112536 148436
rect 112588 148424 112594 148436
rect 145190 148424 145196 148436
rect 112588 148396 145196 148424
rect 112588 148384 112594 148396
rect 145190 148384 145196 148396
rect 145248 148384 145254 148436
rect 158622 148384 158628 148436
rect 158680 148424 158686 148436
rect 196986 148424 196992 148436
rect 158680 148396 196992 148424
rect 158680 148384 158686 148396
rect 196986 148384 196992 148396
rect 197044 148384 197050 148436
rect 98822 148316 98828 148368
rect 98880 148356 98886 148368
rect 132954 148356 132960 148368
rect 98880 148328 132960 148356
rect 98880 148316 98886 148328
rect 132954 148316 132960 148328
rect 133012 148316 133018 148368
rect 155678 148316 155684 148368
rect 155736 148356 155742 148368
rect 217042 148356 217048 148368
rect 155736 148328 217048 148356
rect 155736 148316 155742 148328
rect 217042 148316 217048 148328
rect 217100 148316 217106 148368
rect 164510 148248 164516 148300
rect 164568 148288 164574 148300
rect 191098 148288 191104 148300
rect 164568 148260 191104 148288
rect 164568 148248 164574 148260
rect 191098 148248 191104 148260
rect 191156 148248 191162 148300
rect 177574 148180 177580 148232
rect 177632 148220 177638 148232
rect 199930 148220 199936 148232
rect 177632 148192 199936 148220
rect 177632 148180 177638 148192
rect 199930 148180 199936 148192
rect 199988 148180 199994 148232
rect 180426 148112 180432 148164
rect 180484 148152 180490 148164
rect 193950 148152 193956 148164
rect 180484 148124 193956 148152
rect 180484 148112 180490 148124
rect 193950 148112 193956 148124
rect 194008 148112 194014 148164
rect 128354 147636 128360 147688
rect 128412 147676 128418 147688
rect 128630 147676 128636 147688
rect 128412 147648 128636 147676
rect 128412 147636 128418 147648
rect 128630 147636 128636 147648
rect 128688 147676 128694 147688
rect 136174 147676 136180 147688
rect 128688 147648 136180 147676
rect 128688 147636 128694 147648
rect 136174 147636 136180 147648
rect 136232 147636 136238 147688
rect 169846 147568 169852 147620
rect 169904 147608 169910 147620
rect 196434 147608 196440 147620
rect 169904 147580 196440 147608
rect 169904 147568 169910 147580
rect 196434 147568 196440 147580
rect 196492 147568 196498 147620
rect 172606 147500 172612 147552
rect 172664 147540 172670 147552
rect 198734 147540 198740 147552
rect 172664 147512 198740 147540
rect 172664 147500 172670 147512
rect 198734 147500 198740 147512
rect 198792 147500 198798 147552
rect 117682 147432 117688 147484
rect 117740 147472 117746 147484
rect 132126 147472 132132 147484
rect 117740 147444 132132 147472
rect 117740 147432 117746 147444
rect 132126 147432 132132 147444
rect 132184 147432 132190 147484
rect 171226 147432 171232 147484
rect 171284 147472 171290 147484
rect 180426 147472 180432 147484
rect 171284 147444 180432 147472
rect 171284 147432 171290 147444
rect 180426 147432 180432 147444
rect 180484 147432 180490 147484
rect 113726 147364 113732 147416
rect 113784 147404 113790 147416
rect 130746 147404 130752 147416
rect 113784 147376 130752 147404
rect 113784 147364 113790 147376
rect 130746 147364 130752 147376
rect 130804 147364 130810 147416
rect 179598 147364 179604 147416
rect 179656 147404 179662 147416
rect 197722 147404 197728 147416
rect 179656 147376 197728 147404
rect 179656 147364 179662 147376
rect 197722 147364 197728 147376
rect 197780 147364 197786 147416
rect 111886 147296 111892 147348
rect 111944 147336 111950 147348
rect 130838 147336 130844 147348
rect 111944 147308 130844 147336
rect 111944 147296 111950 147308
rect 130838 147296 130844 147308
rect 130896 147296 130902 147348
rect 179690 147296 179696 147348
rect 179748 147336 179754 147348
rect 199194 147336 199200 147348
rect 179748 147308 199200 147336
rect 179748 147296 179754 147308
rect 199194 147296 199200 147308
rect 199252 147296 199258 147348
rect 109678 147228 109684 147280
rect 109736 147268 109742 147280
rect 132034 147268 132040 147280
rect 109736 147240 132040 147268
rect 109736 147228 109742 147240
rect 132034 147228 132040 147240
rect 132092 147228 132098 147280
rect 161446 147240 166994 147268
rect 116210 147160 116216 147212
rect 116268 147200 116274 147212
rect 143718 147200 143724 147212
rect 116268 147172 143724 147200
rect 116268 147160 116274 147172
rect 143718 147160 143724 147172
rect 143776 147160 143782 147212
rect 156230 147160 156236 147212
rect 156288 147200 156294 147212
rect 161446 147200 161474 147240
rect 156288 147172 161474 147200
rect 156288 147160 156294 147172
rect 113818 147092 113824 147144
rect 113876 147132 113882 147144
rect 143902 147132 143908 147144
rect 113876 147104 143908 147132
rect 113876 147092 113882 147104
rect 143902 147092 143908 147104
rect 143960 147092 143966 147144
rect 166966 147132 166994 147240
rect 178954 147228 178960 147280
rect 179012 147268 179018 147280
rect 197906 147268 197912 147280
rect 179012 147240 197912 147268
rect 179012 147228 179018 147240
rect 197906 147228 197912 147240
rect 197964 147228 197970 147280
rect 179506 147160 179512 147212
rect 179564 147200 179570 147212
rect 199102 147200 199108 147212
rect 179564 147172 199108 147200
rect 179564 147160 179570 147172
rect 199102 147160 199108 147172
rect 199160 147160 199166 147212
rect 180242 147132 180248 147144
rect 166966 147104 180248 147132
rect 180242 147092 180248 147104
rect 180300 147092 180306 147144
rect 198090 147132 198096 147144
rect 180352 147104 198096 147132
rect 110782 147024 110788 147076
rect 110840 147064 110846 147076
rect 143626 147064 143632 147076
rect 110840 147036 143632 147064
rect 110840 147024 110846 147036
rect 143626 147024 143632 147036
rect 143684 147024 143690 147076
rect 171410 147024 171416 147076
rect 171468 147064 171474 147076
rect 180352 147064 180380 147104
rect 198090 147092 198096 147104
rect 198148 147092 198154 147144
rect 171468 147036 180380 147064
rect 171468 147024 171474 147036
rect 180426 147024 180432 147076
rect 180484 147064 180490 147076
rect 198182 147064 198188 147076
rect 180484 147036 198188 147064
rect 180484 147024 180490 147036
rect 198182 147024 198188 147036
rect 198240 147024 198246 147076
rect 109770 146956 109776 147008
rect 109828 146996 109834 147008
rect 143810 146996 143816 147008
rect 109828 146968 143816 146996
rect 109828 146956 109834 146968
rect 143810 146956 143816 146968
rect 143868 146956 143874 147008
rect 157242 146956 157248 147008
rect 157300 146996 157306 147008
rect 193858 146996 193864 147008
rect 157300 146968 193864 146996
rect 157300 146956 157306 146968
rect 193858 146956 193864 146968
rect 193916 146956 193922 147008
rect 109494 146888 109500 146940
rect 109552 146928 109558 146940
rect 145282 146928 145288 146940
rect 109552 146900 145288 146928
rect 109552 146888 109558 146900
rect 145282 146888 145288 146900
rect 145340 146888 145346 146940
rect 146202 146888 146208 146940
rect 146260 146928 146266 146940
rect 184750 146928 184756 146940
rect 146260 146900 184756 146928
rect 146260 146888 146266 146900
rect 184750 146888 184756 146900
rect 184808 146888 184814 146940
rect 185854 146888 185860 146940
rect 185912 146928 185918 146940
rect 186038 146928 186044 146940
rect 185912 146900 186044 146928
rect 185912 146888 185918 146900
rect 186038 146888 186044 146900
rect 186096 146888 186102 146940
rect 185670 146752 185676 146804
rect 185728 146792 185734 146804
rect 186038 146792 186044 146804
rect 185728 146764 186044 146792
rect 185728 146752 185734 146764
rect 186038 146752 186044 146764
rect 186096 146752 186102 146804
rect 176102 146208 176108 146260
rect 176160 146248 176166 146260
rect 194134 146248 194140 146260
rect 176160 146220 194140 146248
rect 176160 146208 176166 146220
rect 194134 146208 194140 146220
rect 194192 146208 194198 146260
rect 120350 146140 120356 146192
rect 120408 146180 120414 146192
rect 131758 146180 131764 146192
rect 120408 146152 131764 146180
rect 120408 146140 120414 146152
rect 131758 146140 131764 146152
rect 131816 146140 131822 146192
rect 178402 146140 178408 146192
rect 178460 146180 178466 146192
rect 196710 146180 196716 146192
rect 178460 146152 196716 146180
rect 178460 146140 178466 146152
rect 196710 146140 196716 146152
rect 196768 146140 196774 146192
rect 117958 146072 117964 146124
rect 118016 146112 118022 146124
rect 129734 146112 129740 146124
rect 118016 146084 129740 146112
rect 118016 146072 118022 146084
rect 129734 146072 129740 146084
rect 129792 146072 129798 146124
rect 177206 146072 177212 146124
rect 177264 146112 177270 146124
rect 199286 146112 199292 146124
rect 177264 146084 199292 146112
rect 177264 146072 177270 146084
rect 199286 146072 199292 146084
rect 199344 146072 199350 146124
rect 115382 146004 115388 146056
rect 115440 146044 115446 146056
rect 131298 146044 131304 146056
rect 115440 146016 131304 146044
rect 115440 146004 115446 146016
rect 131298 146004 131304 146016
rect 131356 146004 131362 146056
rect 157518 146004 157524 146056
rect 157576 146044 157582 146056
rect 188430 146044 188436 146056
rect 157576 146016 188436 146044
rect 157576 146004 157582 146016
rect 188430 146004 188436 146016
rect 188488 146004 188494 146056
rect 114002 145936 114008 145988
rect 114060 145976 114066 145988
rect 130286 145976 130292 145988
rect 114060 145948 130292 145976
rect 114060 145936 114066 145948
rect 130286 145936 130292 145948
rect 130344 145936 130350 145988
rect 159910 145936 159916 145988
rect 159968 145976 159974 145988
rect 192846 145976 192852 145988
rect 159968 145948 192852 145976
rect 159968 145936 159974 145948
rect 192846 145936 192852 145948
rect 192904 145936 192910 145988
rect 111058 145868 111064 145920
rect 111116 145908 111122 145920
rect 126974 145908 126980 145920
rect 111116 145880 126980 145908
rect 111116 145868 111122 145880
rect 126974 145868 126980 145880
rect 127032 145868 127038 145920
rect 161290 145868 161296 145920
rect 161348 145908 161354 145920
rect 194226 145908 194232 145920
rect 161348 145880 194232 145908
rect 161348 145868 161354 145880
rect 194226 145868 194232 145880
rect 194284 145868 194290 145920
rect 120626 145800 120632 145852
rect 120684 145840 120690 145852
rect 143626 145840 143632 145852
rect 120684 145812 143632 145840
rect 120684 145800 120690 145812
rect 143626 145800 143632 145812
rect 143684 145800 143690 145852
rect 155954 145800 155960 145852
rect 156012 145840 156018 145852
rect 189442 145840 189448 145852
rect 156012 145812 189448 145840
rect 156012 145800 156018 145812
rect 189442 145800 189448 145812
rect 189500 145800 189506 145852
rect 117958 145732 117964 145784
rect 118016 145772 118022 145784
rect 146570 145772 146576 145784
rect 118016 145744 146576 145772
rect 118016 145732 118022 145744
rect 146570 145732 146576 145744
rect 146628 145732 146634 145784
rect 160186 145732 160192 145784
rect 160244 145772 160250 145784
rect 195514 145772 195520 145784
rect 160244 145744 195520 145772
rect 160244 145732 160250 145744
rect 195514 145732 195520 145744
rect 195572 145732 195578 145784
rect 115198 145664 115204 145716
rect 115256 145704 115262 145716
rect 148226 145704 148232 145716
rect 115256 145676 148232 145704
rect 115256 145664 115262 145676
rect 148226 145664 148232 145676
rect 148284 145664 148290 145716
rect 162302 145664 162308 145716
rect 162360 145704 162366 145716
rect 196526 145704 196532 145716
rect 162360 145676 196532 145704
rect 162360 145664 162366 145676
rect 196526 145664 196532 145676
rect 196584 145664 196590 145716
rect 112806 145596 112812 145648
rect 112864 145636 112870 145648
rect 145006 145636 145012 145648
rect 112864 145608 145012 145636
rect 112864 145596 112870 145608
rect 145006 145596 145012 145608
rect 145064 145596 145070 145648
rect 156046 145596 156052 145648
rect 156104 145636 156110 145648
rect 191190 145636 191196 145648
rect 156104 145608 191196 145636
rect 156104 145596 156110 145608
rect 191190 145596 191196 145608
rect 191248 145596 191254 145648
rect 3510 145528 3516 145580
rect 3568 145568 3574 145580
rect 3568 145540 161474 145568
rect 3568 145528 3574 145540
rect 161446 145364 161474 145540
rect 183462 145528 183468 145580
rect 183520 145568 183526 145580
rect 197814 145568 197820 145580
rect 183520 145540 197820 145568
rect 183520 145528 183526 145540
rect 197814 145528 197820 145540
rect 197872 145528 197878 145580
rect 178310 145460 178316 145512
rect 178368 145500 178374 145512
rect 195974 145500 195980 145512
rect 178368 145472 195980 145500
rect 178368 145460 178374 145472
rect 195974 145460 195980 145472
rect 196032 145460 196038 145512
rect 178218 145392 178224 145444
rect 178276 145432 178282 145444
rect 193766 145432 193772 145444
rect 178276 145404 193772 145432
rect 178276 145392 178282 145404
rect 193766 145392 193772 145404
rect 193824 145392 193830 145444
rect 179782 145364 179788 145376
rect 161446 145336 179788 145364
rect 179782 145324 179788 145336
rect 179840 145364 179846 145376
rect 192662 145364 192668 145376
rect 179840 145336 192668 145364
rect 179840 145324 179846 145336
rect 192662 145324 192668 145336
rect 192720 145324 192726 145376
rect 118786 144916 118792 144968
rect 118844 144956 118850 144968
rect 182266 144956 182272 144968
rect 118844 144928 182272 144956
rect 118844 144916 118850 144928
rect 182266 144916 182272 144928
rect 182324 144956 182330 144968
rect 183462 144956 183468 144968
rect 182324 144928 183468 144956
rect 182324 144916 182330 144928
rect 183462 144916 183468 144928
rect 183520 144916 183526 144968
rect 116670 144848 116676 144900
rect 116728 144888 116734 144900
rect 133874 144888 133880 144900
rect 116728 144860 133880 144888
rect 116728 144848 116734 144860
rect 133874 144848 133880 144860
rect 133932 144848 133938 144900
rect 184106 144848 184112 144900
rect 184164 144888 184170 144900
rect 196802 144888 196808 144900
rect 184164 144860 196808 144888
rect 184164 144848 184170 144860
rect 196802 144848 196808 144860
rect 196860 144848 196866 144900
rect 112438 144780 112444 144832
rect 112496 144820 112502 144832
rect 130562 144820 130568 144832
rect 112496 144792 130568 144820
rect 112496 144780 112502 144792
rect 130562 144780 130568 144792
rect 130620 144780 130626 144832
rect 177114 144780 177120 144832
rect 177172 144820 177178 144832
rect 195054 144820 195060 144832
rect 177172 144792 195060 144820
rect 177172 144780 177178 144792
rect 195054 144780 195060 144792
rect 195112 144780 195118 144832
rect 119522 144712 119528 144764
rect 119580 144752 119586 144764
rect 138106 144752 138112 144764
rect 119580 144724 138112 144752
rect 119580 144712 119586 144724
rect 138106 144712 138112 144724
rect 138164 144712 138170 144764
rect 172330 144712 172336 144764
rect 172388 144752 172394 144764
rect 185670 144752 185676 144764
rect 172388 144724 185676 144752
rect 172388 144712 172394 144724
rect 185670 144712 185676 144724
rect 185728 144712 185734 144764
rect 115474 144644 115480 144696
rect 115532 144684 115538 144696
rect 135438 144684 135444 144696
rect 115532 144656 135444 144684
rect 115532 144644 115538 144656
rect 135438 144644 135444 144656
rect 135496 144644 135502 144696
rect 172422 144644 172428 144696
rect 172480 144684 172486 144696
rect 196618 144684 196624 144696
rect 172480 144656 196624 144684
rect 172480 144644 172486 144656
rect 196618 144644 196624 144656
rect 196676 144644 196682 144696
rect 120258 144576 120264 144628
rect 120316 144616 120322 144628
rect 150066 144616 150072 144628
rect 120316 144588 150072 144616
rect 120316 144576 120322 144588
rect 150066 144576 150072 144588
rect 150124 144576 150130 144628
rect 165522 144576 165528 144628
rect 165580 144616 165586 144628
rect 193582 144616 193588 144628
rect 165580 144588 193588 144616
rect 165580 144576 165586 144588
rect 193582 144576 193588 144588
rect 193640 144576 193646 144628
rect 118878 144508 118884 144560
rect 118936 144548 118942 144560
rect 151814 144548 151820 144560
rect 118936 144520 151820 144548
rect 118936 144508 118942 144520
rect 151814 144508 151820 144520
rect 151872 144508 151878 144560
rect 163958 144508 163964 144560
rect 164016 144548 164022 144560
rect 192478 144548 192484 144560
rect 164016 144520 192484 144548
rect 164016 144508 164022 144520
rect 192478 144508 192484 144520
rect 192536 144508 192542 144560
rect 119614 144440 119620 144492
rect 119672 144480 119678 144492
rect 152458 144480 152464 144492
rect 119672 144452 152464 144480
rect 119672 144440 119678 144452
rect 152458 144440 152464 144452
rect 152516 144440 152522 144492
rect 154482 144440 154488 144492
rect 154540 144480 154546 144492
rect 187970 144480 187976 144492
rect 154540 144452 187976 144480
rect 154540 144440 154546 144452
rect 187970 144440 187976 144452
rect 188028 144440 188034 144492
rect 117866 144372 117872 144424
rect 117924 144412 117930 144424
rect 151906 144412 151912 144424
rect 117924 144384 151912 144412
rect 117924 144372 117930 144384
rect 151906 144372 151912 144384
rect 151964 144372 151970 144424
rect 157794 144372 157800 144424
rect 157852 144412 157858 144424
rect 192386 144412 192392 144424
rect 157852 144384 192392 144412
rect 157852 144372 157858 144384
rect 192386 144372 192392 144384
rect 192444 144372 192450 144424
rect 103974 144304 103980 144356
rect 104032 144344 104038 144356
rect 145742 144344 145748 144356
rect 104032 144316 145748 144344
rect 104032 144304 104038 144316
rect 145742 144304 145748 144316
rect 145800 144304 145806 144356
rect 159542 144304 159548 144356
rect 159600 144344 159606 144356
rect 193674 144344 193680 144356
rect 159600 144316 193680 144344
rect 159600 144304 159606 144316
rect 193674 144304 193680 144316
rect 193732 144304 193738 144356
rect 112622 144236 112628 144288
rect 112680 144276 112686 144288
rect 131206 144276 131212 144288
rect 112680 144248 131212 144276
rect 112680 144236 112686 144248
rect 131206 144236 131212 144248
rect 131264 144276 131270 144288
rect 188522 144276 188528 144288
rect 131264 144248 188528 144276
rect 131264 144236 131270 144248
rect 188522 144236 188528 144248
rect 188580 144236 188586 144288
rect 116854 144168 116860 144220
rect 116912 144208 116918 144220
rect 130194 144208 130200 144220
rect 116912 144180 130200 144208
rect 116912 144168 116918 144180
rect 130194 144168 130200 144180
rect 130252 144208 130258 144220
rect 189810 144208 189816 144220
rect 130252 144180 189816 144208
rect 130252 144168 130258 144180
rect 189810 144168 189816 144180
rect 189868 144168 189874 144220
rect 113634 144100 113640 144152
rect 113692 144140 113698 144152
rect 130470 144140 130476 144152
rect 113692 144112 130476 144140
rect 113692 144100 113698 144112
rect 130470 144100 130476 144112
rect 130528 144100 130534 144152
rect 185670 144100 185676 144152
rect 185728 144140 185734 144152
rect 192938 144140 192944 144152
rect 185728 144112 192944 144140
rect 185728 144100 185734 144112
rect 192938 144100 192944 144112
rect 192996 144100 193002 144152
rect 112346 144032 112352 144084
rect 112404 144072 112410 144084
rect 122650 144072 122656 144084
rect 112404 144044 122656 144072
rect 112404 144032 112410 144044
rect 122650 144032 122656 144044
rect 122708 144032 122714 144084
rect 117590 143964 117596 144016
rect 117648 144004 117654 144016
rect 128170 144004 128176 144016
rect 117648 143976 128176 144004
rect 117648 143964 117654 143976
rect 128170 143964 128176 143976
rect 128228 143964 128234 144016
rect 125226 143556 125232 143608
rect 125284 143596 125290 143608
rect 126238 143596 126244 143608
rect 125284 143568 126244 143596
rect 125284 143556 125290 143568
rect 126238 143556 126244 143568
rect 126296 143596 126302 143608
rect 580534 143596 580540 143608
rect 126296 143568 580540 143596
rect 126296 143556 126302 143568
rect 580534 143556 580540 143568
rect 580592 143556 580598 143608
rect 118234 143488 118240 143540
rect 118292 143528 118298 143540
rect 128446 143528 128452 143540
rect 118292 143500 128452 143528
rect 118292 143488 118298 143500
rect 128446 143488 128452 143500
rect 128504 143488 128510 143540
rect 147674 143488 147680 143540
rect 147732 143528 147738 143540
rect 150802 143528 150808 143540
rect 147732 143500 150808 143528
rect 147732 143488 147738 143500
rect 150802 143488 150808 143500
rect 150860 143488 150866 143540
rect 170030 143488 170036 143540
rect 170088 143528 170094 143540
rect 170306 143528 170312 143540
rect 170088 143500 170312 143528
rect 170088 143488 170094 143500
rect 170306 143488 170312 143500
rect 170364 143488 170370 143540
rect 172882 143488 172888 143540
rect 172940 143528 172946 143540
rect 173526 143528 173532 143540
rect 172940 143500 173532 143528
rect 172940 143488 172946 143500
rect 173526 143488 173532 143500
rect 173584 143488 173590 143540
rect 174262 143488 174268 143540
rect 174320 143528 174326 143540
rect 179690 143528 179696 143540
rect 174320 143500 179696 143528
rect 174320 143488 174326 143500
rect 179690 143488 179696 143500
rect 179748 143488 179754 143540
rect 185762 143488 185768 143540
rect 185820 143528 185826 143540
rect 189350 143528 189356 143540
rect 185820 143500 189356 143528
rect 185820 143488 185826 143500
rect 189350 143488 189356 143500
rect 189408 143488 189414 143540
rect 131482 143460 131488 143472
rect 118666 143432 131488 143460
rect 118326 143352 118332 143404
rect 118384 143392 118390 143404
rect 118666 143392 118694 143432
rect 131482 143420 131488 143432
rect 131540 143420 131546 143472
rect 176286 143420 176292 143472
rect 176344 143460 176350 143472
rect 179598 143460 179604 143472
rect 176344 143432 179604 143460
rect 176344 143420 176350 143432
rect 179598 143420 179604 143432
rect 179656 143420 179662 143472
rect 181530 143420 181536 143472
rect 181588 143460 181594 143472
rect 187970 143460 187976 143472
rect 181588 143432 187976 143460
rect 181588 143420 181594 143432
rect 187970 143420 187976 143432
rect 188028 143420 188034 143472
rect 188062 143420 188068 143472
rect 188120 143460 188126 143472
rect 191374 143460 191380 143472
rect 188120 143432 191380 143460
rect 188120 143420 188126 143432
rect 191374 143420 191380 143432
rect 191432 143420 191438 143472
rect 130378 143392 130384 143404
rect 118384 143364 118694 143392
rect 120920 143364 130384 143392
rect 118384 143352 118390 143364
rect 115290 143216 115296 143268
rect 115348 143256 115354 143268
rect 120920 143256 120948 143364
rect 130378 143352 130384 143364
rect 130436 143352 130442 143404
rect 131114 143352 131120 143404
rect 131172 143392 131178 143404
rect 137554 143392 137560 143404
rect 131172 143364 137560 143392
rect 131172 143352 131178 143364
rect 137554 143352 137560 143364
rect 137612 143352 137618 143404
rect 175734 143352 175740 143404
rect 175792 143392 175798 143404
rect 178310 143392 178316 143404
rect 175792 143364 178316 143392
rect 175792 143352 175798 143364
rect 178310 143352 178316 143364
rect 178368 143352 178374 143404
rect 178862 143352 178868 143404
rect 178920 143392 178926 143404
rect 190270 143392 190276 143404
rect 178920 143364 190276 143392
rect 178920 143352 178926 143364
rect 190270 143352 190276 143364
rect 190328 143352 190334 143404
rect 120994 143284 121000 143336
rect 121052 143324 121058 143336
rect 134794 143324 134800 143336
rect 121052 143296 134800 143324
rect 121052 143284 121058 143296
rect 134794 143284 134800 143296
rect 134852 143284 134858 143336
rect 170950 143284 170956 143336
rect 171008 143324 171014 143336
rect 179506 143324 179512 143336
rect 171008 143296 179512 143324
rect 171008 143284 171014 143296
rect 179506 143284 179512 143296
rect 179564 143284 179570 143336
rect 181714 143284 181720 143336
rect 181772 143324 181778 143336
rect 193490 143324 193496 143336
rect 181772 143296 193496 143324
rect 181772 143284 181778 143296
rect 193490 143284 193496 143296
rect 193548 143284 193554 143336
rect 115348 143228 120948 143256
rect 115348 143216 115354 143228
rect 129734 143216 129740 143268
rect 129792 143256 129798 143268
rect 137002 143256 137008 143268
rect 129792 143228 137008 143256
rect 129792 143216 129798 143228
rect 137002 143216 137008 143228
rect 137060 143216 137066 143268
rect 169662 143216 169668 143268
rect 169720 143256 169726 143268
rect 179414 143256 179420 143268
rect 169720 143228 179420 143256
rect 169720 143216 169726 143228
rect 179414 143216 179420 143228
rect 179472 143216 179478 143268
rect 184290 143216 184296 143268
rect 184348 143256 184354 143268
rect 196434 143256 196440 143268
rect 184348 143228 196440 143256
rect 184348 143216 184354 143228
rect 196434 143216 196440 143228
rect 196492 143216 196498 143268
rect 116762 143148 116768 143200
rect 116820 143188 116826 143200
rect 133138 143188 133144 143200
rect 116820 143160 133144 143188
rect 116820 143148 116826 143160
rect 133138 143148 133144 143160
rect 133196 143148 133202 143200
rect 173158 143148 173164 143200
rect 173216 143188 173222 143200
rect 190638 143188 190644 143200
rect 173216 143160 190644 143188
rect 173216 143148 173222 143160
rect 190638 143148 190644 143160
rect 190696 143148 190702 143200
rect 120902 143080 120908 143132
rect 120960 143120 120966 143132
rect 139762 143120 139768 143132
rect 120960 143092 139768 143120
rect 120960 143080 120966 143092
rect 139762 143080 139768 143092
rect 139820 143080 139826 143132
rect 168190 143080 168196 143132
rect 168248 143120 168254 143132
rect 181346 143120 181352 143132
rect 168248 143092 181352 143120
rect 168248 143080 168254 143092
rect 181346 143080 181352 143092
rect 181404 143080 181410 143132
rect 181438 143080 181444 143132
rect 181496 143120 181502 143132
rect 188062 143120 188068 143132
rect 181496 143092 188068 143120
rect 181496 143080 181502 143092
rect 188062 143080 188068 143092
rect 188120 143080 188126 143132
rect 119706 143012 119712 143064
rect 119764 143052 119770 143064
rect 141418 143052 141424 143064
rect 119764 143024 141424 143052
rect 119764 143012 119770 143024
rect 141418 143012 141424 143024
rect 141476 143012 141482 143064
rect 166626 143012 166632 143064
rect 166684 143052 166690 143064
rect 190914 143052 190920 143064
rect 166684 143024 190920 143052
rect 166684 143012 166690 143024
rect 190914 143012 190920 143024
rect 190972 143012 190978 143064
rect 119338 142944 119344 142996
rect 119396 142984 119402 142996
rect 144914 142984 144920 142996
rect 119396 142956 144920 142984
rect 119396 142944 119402 142956
rect 144914 142944 144920 142956
rect 144972 142944 144978 142996
rect 154298 142944 154304 142996
rect 154356 142984 154362 142996
rect 188246 142984 188252 142996
rect 154356 142956 188252 142984
rect 154356 142944 154362 142956
rect 188246 142944 188252 142956
rect 188304 142944 188310 142996
rect 119430 142876 119436 142928
rect 119488 142916 119494 142928
rect 148042 142916 148048 142928
rect 119488 142888 148048 142916
rect 119488 142876 119494 142888
rect 148042 142876 148048 142888
rect 148100 142876 148106 142928
rect 168374 142876 168380 142928
rect 168432 142916 168438 142928
rect 209222 142916 209228 142928
rect 168432 142888 209228 142916
rect 168432 142876 168438 142888
rect 209222 142876 209228 142888
rect 209280 142876 209286 142928
rect 116854 142808 116860 142860
rect 116912 142848 116918 142860
rect 149698 142848 149704 142860
rect 116912 142820 149704 142848
rect 116912 142808 116918 142820
rect 149698 142808 149704 142820
rect 149756 142808 149762 142860
rect 155494 142808 155500 142860
rect 155552 142848 155558 142860
rect 207842 142848 207848 142860
rect 155552 142820 207848 142848
rect 155552 142808 155558 142820
rect 207842 142808 207848 142820
rect 207900 142808 207906 142860
rect 186038 142740 186044 142792
rect 186096 142780 186102 142792
rect 192662 142780 192668 142792
rect 186096 142752 192668 142780
rect 186096 142740 186102 142752
rect 192662 142740 192668 142752
rect 192720 142740 192726 142792
rect 181346 142672 181352 142724
rect 181404 142712 181410 142724
rect 189534 142712 189540 142724
rect 181404 142684 189540 142712
rect 181404 142672 181410 142684
rect 189534 142672 189540 142684
rect 189592 142672 189598 142724
rect 188062 142604 188068 142656
rect 188120 142644 188126 142656
rect 188706 142644 188712 142656
rect 188120 142616 188712 142644
rect 188120 142604 188126 142616
rect 188706 142604 188712 142616
rect 188764 142604 188770 142656
rect 127526 142400 127532 142452
rect 127584 142440 127590 142452
rect 127802 142440 127808 142452
rect 127584 142412 127808 142440
rect 127584 142400 127590 142412
rect 127802 142400 127808 142412
rect 127860 142400 127866 142452
rect 123110 142332 123116 142384
rect 123168 142372 123174 142384
rect 123938 142372 123944 142384
rect 123168 142344 123944 142372
rect 123168 142332 123174 142344
rect 123938 142332 123944 142344
rect 123996 142332 124002 142384
rect 126054 142332 126060 142384
rect 126112 142372 126118 142384
rect 126422 142372 126428 142384
rect 126112 142344 126428 142372
rect 126112 142332 126118 142344
rect 126422 142332 126428 142344
rect 126480 142332 126486 142384
rect 40678 142264 40684 142316
rect 40736 142304 40742 142316
rect 184290 142304 184296 142316
rect 40736 142276 184296 142304
rect 40736 142264 40742 142276
rect 184290 142264 184296 142276
rect 184348 142264 184354 142316
rect 120994 142196 121000 142248
rect 121052 142236 121058 142248
rect 146386 142236 146392 142248
rect 121052 142208 146392 142236
rect 121052 142196 121058 142208
rect 146386 142196 146392 142208
rect 146444 142196 146450 142248
rect 184014 142196 184020 142248
rect 184072 142236 184078 142248
rect 192570 142236 192576 142248
rect 184072 142208 192576 142236
rect 184072 142196 184078 142208
rect 192570 142196 192576 142208
rect 192628 142196 192634 142248
rect 129826 142128 129832 142180
rect 129884 142168 129890 142180
rect 134242 142168 134248 142180
rect 129884 142140 134248 142168
rect 129884 142128 129890 142140
rect 134242 142128 134248 142140
rect 134300 142128 134306 142180
rect 150526 142168 150532 142180
rect 148934 142140 150532 142168
rect 117038 142060 117044 142112
rect 117096 142100 117102 142112
rect 117096 142072 125548 142100
rect 117096 142060 117102 142072
rect 118050 141992 118056 142044
rect 118108 142032 118114 142044
rect 123478 142032 123484 142044
rect 118108 142004 123484 142032
rect 118108 141992 118114 142004
rect 123478 141992 123484 142004
rect 123536 141992 123542 142044
rect 125520 142032 125548 142072
rect 125594 142060 125600 142112
rect 125652 142100 125658 142112
rect 148934 142100 148962 142140
rect 150526 142128 150532 142140
rect 150584 142128 150590 142180
rect 155862 142128 155868 142180
rect 155920 142168 155926 142180
rect 157334 142168 157340 142180
rect 155920 142140 157340 142168
rect 155920 142128 155926 142140
rect 157334 142128 157340 142140
rect 157392 142128 157398 142180
rect 159174 142128 159180 142180
rect 159232 142168 159238 142180
rect 159232 142140 161520 142168
rect 159232 142128 159238 142140
rect 125652 142072 148962 142100
rect 161492 142100 161520 142140
rect 192202 142100 192208 142112
rect 161492 142072 192208 142100
rect 125652 142060 125658 142072
rect 192202 142060 192208 142072
rect 192260 142060 192266 142112
rect 126514 142032 126520 142044
rect 125520 142004 126520 142032
rect 126514 141992 126520 142004
rect 126572 141992 126578 142044
rect 184106 141992 184112 142044
rect 184164 142032 184170 142044
rect 184382 142032 184388 142044
rect 184164 142004 184388 142032
rect 184164 141992 184170 142004
rect 184382 141992 184388 142004
rect 184440 141992 184446 142044
rect 184474 141992 184480 142044
rect 184532 142032 184538 142044
rect 184842 142032 184848 142044
rect 184532 142004 184848 142032
rect 184532 141992 184538 142004
rect 184842 141992 184848 142004
rect 184900 141992 184906 142044
rect 186130 141992 186136 142044
rect 186188 142032 186194 142044
rect 196618 142032 196624 142044
rect 186188 142004 196624 142032
rect 186188 141992 186194 142004
rect 196618 141992 196624 142004
rect 196676 141992 196682 142044
rect 114094 141924 114100 141976
rect 114152 141964 114158 141976
rect 125594 141964 125600 141976
rect 114152 141936 125600 141964
rect 114152 141924 114158 141936
rect 125594 141924 125600 141936
rect 125652 141924 125658 141976
rect 186222 141924 186228 141976
rect 186280 141964 186286 141976
rect 186866 141964 186872 141976
rect 186280 141936 186872 141964
rect 186280 141924 186286 141936
rect 186866 141924 186872 141936
rect 186924 141924 186930 141976
rect 187142 141924 187148 141976
rect 187200 141964 187206 141976
rect 196710 141964 196716 141976
rect 187200 141936 196716 141964
rect 187200 141924 187206 141936
rect 196710 141924 196716 141936
rect 196768 141924 196774 141976
rect 114186 141856 114192 141908
rect 114244 141896 114250 141908
rect 127066 141896 127072 141908
rect 114244 141868 127072 141896
rect 114244 141856 114250 141868
rect 127066 141856 127072 141868
rect 127124 141856 127130 141908
rect 180334 141856 180340 141908
rect 180392 141896 180398 141908
rect 194962 141896 194968 141908
rect 180392 141868 194968 141896
rect 180392 141856 180398 141868
rect 194962 141856 194968 141868
rect 195020 141856 195026 141908
rect 112898 141788 112904 141840
rect 112956 141828 112962 141840
rect 129274 141828 129280 141840
rect 112956 141800 129280 141828
rect 112956 141788 112962 141800
rect 129274 141788 129280 141800
rect 129332 141788 129338 141840
rect 176470 141788 176476 141840
rect 176528 141828 176534 141840
rect 192294 141828 192300 141840
rect 176528 141800 192300 141828
rect 176528 141788 176534 141800
rect 192294 141788 192300 141800
rect 192352 141788 192358 141840
rect 118142 141720 118148 141772
rect 118200 141760 118206 141772
rect 140314 141760 140320 141772
rect 118200 141732 140320 141760
rect 118200 141720 118206 141732
rect 140314 141720 140320 141732
rect 140372 141720 140378 141772
rect 170490 141720 170496 141772
rect 170548 141760 170554 141772
rect 185302 141760 185308 141772
rect 170548 141732 185308 141760
rect 170548 141720 170554 141732
rect 185302 141720 185308 141732
rect 185360 141720 185366 141772
rect 185946 141720 185952 141772
rect 186004 141760 186010 141772
rect 187142 141760 187148 141772
rect 186004 141732 187148 141760
rect 186004 141720 186010 141732
rect 187142 141720 187148 141732
rect 187200 141720 187206 141772
rect 123478 141652 123484 141704
rect 123536 141692 123542 141704
rect 136634 141692 136640 141704
rect 123536 141664 136640 141692
rect 123536 141652 123542 141664
rect 136634 141652 136640 141664
rect 136692 141652 136698 141704
rect 180150 141652 180156 141704
rect 180208 141692 180214 141704
rect 199286 141692 199292 141704
rect 180208 141664 199292 141692
rect 180208 141652 180214 141664
rect 199286 141652 199292 141664
rect 199344 141652 199350 141704
rect 113082 141584 113088 141636
rect 113140 141624 113146 141636
rect 139394 141624 139400 141636
rect 113140 141596 139400 141624
rect 113140 141584 113146 141596
rect 139394 141584 139400 141596
rect 139452 141584 139458 141636
rect 164234 141584 164240 141636
rect 164292 141624 164298 141636
rect 187326 141624 187332 141636
rect 164292 141596 187332 141624
rect 164292 141584 164298 141596
rect 187326 141584 187332 141596
rect 187384 141584 187390 141636
rect 119798 141516 119804 141568
rect 119856 141556 119862 141568
rect 153746 141556 153752 141568
rect 119856 141528 153752 141556
rect 119856 141516 119862 141528
rect 153746 141516 153752 141528
rect 153804 141516 153810 141568
rect 167454 141516 167460 141568
rect 167512 141556 167518 141568
rect 192110 141556 192116 141568
rect 167512 141528 192116 141556
rect 167512 141516 167518 141528
rect 192110 141516 192116 141528
rect 192168 141516 192174 141568
rect 119246 141448 119252 141500
rect 119304 141488 119310 141500
rect 158070 141488 158076 141500
rect 119304 141460 158076 141488
rect 119304 141448 119310 141460
rect 158070 141448 158076 141460
rect 158128 141448 158134 141500
rect 166442 141448 166448 141500
rect 166500 141488 166506 141500
rect 217318 141488 217324 141500
rect 166500 141460 217324 141488
rect 166500 141448 166506 141460
rect 217318 141448 217324 141460
rect 217376 141448 217382 141500
rect 119614 141380 119620 141432
rect 119672 141420 119678 141432
rect 149882 141420 149888 141432
rect 119672 141392 149888 141420
rect 119672 141380 119678 141392
rect 149882 141380 149888 141392
rect 149940 141380 149946 141432
rect 151262 141380 151268 141432
rect 151320 141420 151326 141432
rect 214558 141420 214564 141432
rect 151320 141392 214564 141420
rect 151320 141380 151326 141392
rect 214558 141380 214564 141392
rect 214616 141380 214622 141432
rect 116578 141312 116584 141364
rect 116636 141352 116642 141364
rect 116636 141324 118694 141352
rect 116636 141312 116642 141324
rect 118666 141284 118694 141324
rect 119982 141312 119988 141364
rect 120040 141352 120046 141364
rect 123202 141352 123208 141364
rect 120040 141324 123208 141352
rect 120040 141312 120046 141324
rect 123202 141312 123208 141324
rect 123260 141312 123266 141364
rect 184750 141312 184756 141364
rect 184808 141352 184814 141364
rect 195054 141352 195060 141364
rect 184808 141324 195060 141352
rect 184808 141312 184814 141324
rect 195054 141312 195060 141324
rect 195112 141312 195118 141364
rect 127986 141284 127992 141296
rect 118666 141256 127992 141284
rect 127986 141244 127992 141256
rect 128044 141244 128050 141296
rect 184658 141244 184664 141296
rect 184716 141284 184722 141296
rect 194962 141284 194968 141296
rect 184716 141256 194968 141284
rect 184716 141244 184722 141256
rect 194962 141244 194968 141256
rect 195020 141244 195026 141296
rect 185302 141176 185308 141228
rect 185360 141216 185366 141228
rect 189810 141216 189816 141228
rect 185360 141188 189816 141216
rect 185360 141176 185366 141188
rect 189810 141176 189816 141188
rect 189868 141176 189874 141228
rect 117038 140972 117044 141024
rect 117096 141012 117102 141024
rect 124950 141012 124956 141024
rect 117096 140984 124956 141012
rect 117096 140972 117102 140984
rect 124950 140972 124956 140984
rect 125008 140972 125014 141024
rect 116394 140904 116400 140956
rect 116452 140944 116458 140956
rect 123294 140944 123300 140956
rect 116452 140916 123300 140944
rect 116452 140904 116458 140916
rect 123294 140904 123300 140916
rect 123352 140904 123358 140956
rect 123386 140904 123392 140956
rect 123444 140944 123450 140956
rect 142246 140944 142252 140956
rect 123444 140916 142252 140944
rect 123444 140904 123450 140916
rect 142246 140904 142252 140916
rect 142304 140904 142310 140956
rect 97350 140836 97356 140888
rect 97408 140876 97414 140888
rect 181714 140876 181720 140888
rect 97408 140848 181720 140876
rect 97408 140836 97414 140848
rect 181714 140836 181720 140848
rect 181772 140836 181778 140888
rect 13078 140768 13084 140820
rect 13136 140808 13142 140820
rect 182910 140808 182916 140820
rect 13136 140780 182916 140808
rect 13136 140768 13142 140780
rect 182910 140768 182916 140780
rect 182968 140768 182974 140820
rect 120810 140700 120816 140752
rect 120868 140740 120874 140752
rect 126606 140740 126612 140752
rect 120868 140712 126612 140740
rect 120868 140700 120874 140712
rect 126606 140700 126612 140712
rect 126664 140700 126670 140752
rect 131298 140700 131304 140752
rect 131356 140740 131362 140752
rect 132034 140740 132040 140752
rect 131356 140712 132040 140740
rect 131356 140700 131362 140712
rect 132034 140700 132040 140712
rect 132092 140700 132098 140752
rect 145006 140700 145012 140752
rect 145064 140740 145070 140752
rect 145834 140740 145840 140752
rect 145064 140712 145840 140740
rect 145064 140700 145070 140712
rect 145834 140700 145840 140712
rect 145892 140700 145898 140752
rect 183554 140700 183560 140752
rect 183612 140740 183618 140752
rect 184474 140740 184480 140752
rect 183612 140712 184480 140740
rect 183612 140700 183618 140712
rect 184474 140700 184480 140712
rect 184532 140700 184538 140752
rect 120534 140632 120540 140684
rect 120592 140672 120598 140684
rect 126422 140672 126428 140684
rect 120592 140644 126428 140672
rect 120592 140632 120598 140644
rect 126422 140632 126428 140644
rect 126480 140632 126486 140684
rect 184198 140632 184204 140684
rect 184256 140672 184262 140684
rect 192386 140672 192392 140684
rect 184256 140644 192392 140672
rect 184256 140632 184262 140644
rect 192386 140632 192392 140644
rect 192444 140632 192450 140684
rect 118142 140564 118148 140616
rect 118200 140604 118206 140616
rect 121730 140604 121736 140616
rect 118200 140576 121736 140604
rect 118200 140564 118206 140576
rect 121730 140564 121736 140576
rect 121788 140564 121794 140616
rect 121914 140564 121920 140616
rect 121972 140604 121978 140616
rect 125042 140604 125048 140616
rect 121972 140576 125048 140604
rect 121972 140564 121978 140576
rect 125042 140564 125048 140576
rect 125100 140564 125106 140616
rect 184842 140564 184848 140616
rect 184900 140604 184906 140616
rect 192294 140604 192300 140616
rect 184900 140576 192300 140604
rect 184900 140564 184906 140576
rect 192294 140564 192300 140576
rect 192352 140564 192358 140616
rect 118050 140496 118056 140548
rect 118108 140536 118114 140548
rect 118108 140508 118832 140536
rect 118108 140496 118114 140508
rect 115382 140360 115388 140412
rect 115440 140400 115446 140412
rect 118326 140400 118332 140412
rect 115440 140372 118332 140400
rect 115440 140360 115446 140372
rect 118326 140360 118332 140372
rect 118384 140360 118390 140412
rect 118804 140400 118832 140508
rect 119798 140496 119804 140548
rect 119856 140536 119862 140548
rect 126146 140536 126152 140548
rect 119856 140508 126152 140536
rect 119856 140496 119862 140508
rect 126146 140496 126152 140508
rect 126204 140496 126210 140548
rect 185578 140496 185584 140548
rect 185636 140536 185642 140548
rect 195330 140536 195336 140548
rect 185636 140508 195336 140536
rect 185636 140496 185642 140508
rect 195330 140496 195336 140508
rect 195388 140496 195394 140548
rect 119154 140428 119160 140480
rect 119212 140468 119218 140480
rect 126698 140468 126704 140480
rect 119212 140440 126704 140468
rect 119212 140428 119218 140440
rect 126698 140428 126704 140440
rect 126756 140428 126762 140480
rect 180058 140428 180064 140480
rect 180116 140468 180122 140480
rect 190638 140468 190644 140480
rect 180116 140440 190644 140468
rect 180116 140428 180122 140440
rect 190638 140428 190644 140440
rect 190696 140428 190702 140480
rect 126330 140400 126336 140412
rect 118804 140372 126336 140400
rect 126330 140360 126336 140372
rect 126388 140360 126394 140412
rect 178770 140360 178776 140412
rect 178828 140400 178834 140412
rect 190822 140400 190828 140412
rect 178828 140372 190828 140400
rect 178828 140360 178834 140372
rect 190822 140360 190828 140372
rect 190880 140360 190886 140412
rect 125502 140292 125508 140344
rect 125560 140332 125566 140344
rect 138382 140332 138388 140344
rect 125560 140304 138388 140332
rect 125560 140292 125566 140304
rect 138382 140292 138388 140304
rect 138440 140292 138446 140344
rect 178678 140292 178684 140344
rect 178736 140332 178742 140344
rect 190730 140332 190736 140344
rect 178736 140304 190736 140332
rect 178736 140292 178742 140304
rect 190730 140292 190736 140304
rect 190788 140292 190794 140344
rect 115014 140224 115020 140276
rect 115072 140264 115078 140276
rect 128998 140264 129004 140276
rect 115072 140236 118556 140264
rect 115072 140224 115078 140236
rect 112254 140156 112260 140208
rect 112312 140196 112318 140208
rect 117038 140196 117044 140208
rect 112312 140168 117044 140196
rect 112312 140156 112318 140168
rect 117038 140156 117044 140168
rect 117096 140156 117102 140208
rect 118528 140128 118556 140236
rect 119632 140236 129004 140264
rect 119632 140128 119660 140236
rect 128998 140224 129004 140236
rect 129056 140224 129062 140276
rect 164142 140224 164148 140276
rect 164200 140264 164206 140276
rect 187142 140264 187148 140276
rect 164200 140236 187148 140264
rect 164200 140224 164206 140236
rect 187142 140224 187148 140236
rect 187200 140224 187206 140276
rect 124490 140156 124496 140208
rect 124548 140196 124554 140208
rect 139670 140196 139676 140208
rect 124548 140168 139676 140196
rect 124548 140156 124554 140168
rect 139670 140156 139676 140168
rect 139728 140156 139734 140208
rect 162946 140156 162952 140208
rect 163004 140196 163010 140208
rect 197906 140196 197912 140208
rect 163004 140168 197912 140196
rect 163004 140156 163010 140168
rect 197906 140156 197912 140168
rect 197964 140156 197970 140208
rect 118528 140100 119660 140128
rect 119706 140088 119712 140140
rect 119764 140128 119770 140140
rect 150986 140128 150992 140140
rect 119764 140100 150992 140128
rect 119764 140088 119770 140100
rect 150986 140088 150992 140100
rect 151044 140088 151050 140140
rect 157426 140088 157432 140140
rect 157484 140128 157490 140140
rect 192570 140128 192576 140140
rect 157484 140100 192576 140128
rect 157484 140088 157490 140100
rect 192570 140088 192576 140100
rect 192628 140088 192634 140140
rect 121730 140020 121736 140072
rect 121788 140060 121794 140072
rect 126054 140060 126060 140072
rect 121788 140032 126060 140060
rect 121788 140020 121794 140032
rect 126054 140020 126060 140032
rect 126112 140020 126118 140072
rect 148134 140060 148140 140072
rect 132466 140032 148140 140060
rect 118326 139952 118332 140004
rect 118384 139992 118390 140004
rect 127618 139992 127624 140004
rect 118384 139964 127624 139992
rect 118384 139952 118390 139964
rect 127618 139952 127624 139964
rect 127676 139952 127682 140004
rect 116854 139884 116860 139936
rect 116912 139924 116918 139936
rect 132466 139924 132494 140032
rect 148134 140020 148140 140032
rect 148192 140020 148198 140072
rect 156782 140020 156788 140072
rect 156840 140060 156846 140072
rect 197814 140060 197820 140072
rect 156840 140032 197820 140060
rect 156840 140020 156846 140032
rect 197814 140020 197820 140032
rect 197872 140020 197878 140072
rect 116912 139896 132494 139924
rect 116912 139884 116918 139896
rect 172974 139680 172980 139732
rect 173032 139720 173038 139732
rect 197630 139720 197636 139732
rect 173032 139692 197636 139720
rect 173032 139680 173038 139692
rect 197630 139680 197636 139692
rect 197688 139680 197694 139732
rect 161290 139612 161296 139664
rect 161348 139652 161354 139664
rect 194870 139652 194876 139664
rect 161348 139624 194876 139652
rect 161348 139612 161354 139624
rect 194870 139612 194876 139624
rect 194928 139612 194934 139664
rect 123386 139544 123392 139596
rect 123444 139584 123450 139596
rect 183554 139584 183560 139596
rect 123444 139556 183560 139584
rect 123444 139544 123450 139556
rect 183554 139544 183560 139556
rect 183612 139544 183618 139596
rect 118694 139476 118700 139528
rect 118752 139516 118758 139528
rect 180058 139516 180064 139528
rect 118752 139488 180064 139516
rect 118752 139476 118758 139488
rect 180058 139476 180064 139488
rect 180116 139476 180122 139528
rect 183278 139476 183284 139528
rect 183336 139516 183342 139528
rect 189626 139516 189632 139528
rect 183336 139488 189632 139516
rect 183336 139476 183342 139488
rect 189626 139476 189632 139488
rect 189684 139476 189690 139528
rect 125870 139408 125876 139460
rect 125928 139448 125934 139460
rect 327718 139448 327724 139460
rect 125928 139420 327724 139448
rect 125928 139408 125934 139420
rect 327718 139408 327724 139420
rect 327776 139408 327782 139460
rect 188614 139204 188620 139256
rect 188672 139244 188678 139256
rect 189718 139244 189724 139256
rect 188672 139216 189724 139244
rect 188672 139204 188678 139216
rect 189718 139204 189724 139216
rect 189776 139204 189782 139256
rect 189902 138660 189908 138712
rect 189960 138700 189966 138712
rect 195238 138700 195244 138712
rect 189960 138672 195244 138700
rect 189960 138660 189966 138672
rect 195238 138660 195244 138672
rect 195296 138660 195302 138712
rect 3418 137980 3424 138032
rect 3476 138020 3482 138032
rect 120994 138020 121000 138032
rect 3476 137992 121000 138020
rect 3476 137980 3482 137992
rect 120994 137980 121000 137992
rect 121052 137980 121058 138032
rect 3234 137912 3240 137964
rect 3292 137952 3298 137964
rect 118694 137952 118700 137964
rect 3292 137924 118700 137952
rect 3292 137912 3298 137924
rect 118694 137912 118700 137924
rect 118752 137912 118758 137964
rect 120258 137300 120264 137352
rect 120316 137340 120322 137352
rect 120626 137340 120632 137352
rect 120316 137312 120632 137340
rect 120316 137300 120322 137312
rect 120626 137300 120632 137312
rect 120684 137300 120690 137352
rect 117866 136144 117872 136196
rect 117924 136184 117930 136196
rect 119798 136184 119804 136196
rect 117924 136156 119804 136184
rect 117924 136144 117930 136156
rect 119798 136144 119804 136156
rect 119856 136144 119862 136196
rect 3050 111392 3056 111444
rect 3108 111432 3114 111444
rect 8938 111432 8944 111444
rect 3108 111404 8944 111432
rect 3108 111392 3114 111404
rect 8938 111392 8944 111404
rect 8996 111392 9002 111444
rect 467098 100648 467104 100700
rect 467156 100688 467162 100700
rect 580166 100688 580172 100700
rect 467156 100660 580172 100688
rect 467156 100648 467162 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 188982 99356 188988 99408
rect 189040 99396 189046 99408
rect 189810 99396 189816 99408
rect 189040 99368 189816 99396
rect 189040 99356 189046 99368
rect 189810 99356 189816 99368
rect 189868 99356 189874 99408
rect 190362 98200 190368 98252
rect 190420 98240 190426 98252
rect 192662 98240 192668 98252
rect 190420 98212 192668 98240
rect 190420 98200 190426 98212
rect 192662 98200 192668 98212
rect 192720 98200 192726 98252
rect 188890 92488 188896 92540
rect 188948 92528 188954 92540
rect 191834 92528 191840 92540
rect 188948 92500 191840 92528
rect 188948 92488 188954 92500
rect 191834 92488 191840 92500
rect 191892 92488 191898 92540
rect 464338 86912 464344 86964
rect 464396 86952 464402 86964
rect 579982 86952 579988 86964
rect 464396 86924 579988 86952
rect 464396 86912 464402 86924
rect 579982 86912 579988 86924
rect 580040 86912 580046 86964
rect 3510 85484 3516 85536
rect 3568 85524 3574 85536
rect 97350 85524 97356 85536
rect 3568 85496 97356 85524
rect 3568 85484 3574 85496
rect 97350 85484 97356 85496
rect 97408 85484 97414 85536
rect 186958 81472 186964 81524
rect 187016 81512 187022 81524
rect 187418 81512 187424 81524
rect 187016 81484 187424 81512
rect 187016 81472 187022 81484
rect 187418 81472 187424 81484
rect 187476 81472 187482 81524
rect 186682 81404 186688 81456
rect 186740 81444 186746 81456
rect 187510 81444 187516 81456
rect 186740 81416 187516 81444
rect 186740 81404 186746 81416
rect 187510 81404 187516 81416
rect 187568 81404 187574 81456
rect 155926 81280 167776 81308
rect 155926 81172 155954 81280
rect 154546 81144 155954 81172
rect 159514 81212 164234 81240
rect 112346 81064 112352 81116
rect 112404 81104 112410 81116
rect 121822 81104 121828 81116
rect 112404 81076 121828 81104
rect 112404 81064 112410 81076
rect 121822 81064 121828 81076
rect 121880 81064 121886 81116
rect 122282 80996 122288 81048
rect 122340 81036 122346 81048
rect 122340 81008 145834 81036
rect 122340 80996 122346 81008
rect 114922 80928 114928 80980
rect 114980 80968 114986 80980
rect 114980 80940 144638 80968
rect 114980 80928 114986 80940
rect 117958 80860 117964 80912
rect 118016 80900 118022 80912
rect 118016 80872 143534 80900
rect 118016 80860 118022 80872
rect 113910 80792 113916 80844
rect 113968 80832 113974 80844
rect 113968 80804 131114 80832
rect 113968 80792 113974 80804
rect 112254 80724 112260 80776
rect 112312 80764 112318 80776
rect 131086 80764 131114 80804
rect 131316 80804 139394 80832
rect 112312 80736 130516 80764
rect 131086 80736 131252 80764
rect 112312 80724 112318 80736
rect 113634 80656 113640 80708
rect 113692 80696 113698 80708
rect 113692 80668 130332 80696
rect 113692 80656 113698 80668
rect 121822 80588 121828 80640
rect 121880 80628 121886 80640
rect 125594 80628 125600 80640
rect 121880 80600 125600 80628
rect 121880 80588 121886 80600
rect 125594 80588 125600 80600
rect 125652 80588 125658 80640
rect 105262 80520 105268 80572
rect 105320 80560 105326 80572
rect 105630 80560 105636 80572
rect 105320 80532 105636 80560
rect 105320 80520 105326 80532
rect 105630 80520 105636 80532
rect 105688 80520 105694 80572
rect 130304 80560 130332 80668
rect 130488 80640 130516 80736
rect 130580 80668 131114 80696
rect 130470 80588 130476 80640
rect 130528 80588 130534 80640
rect 130580 80560 130608 80668
rect 131086 80640 131114 80668
rect 131086 80600 131120 80640
rect 131114 80588 131120 80600
rect 131172 80588 131178 80640
rect 130304 80532 130608 80560
rect 131224 80560 131252 80736
rect 131316 80640 131344 80804
rect 131298 80588 131304 80640
rect 131356 80588 131362 80640
rect 139366 80628 139394 80804
rect 139366 80600 143350 80628
rect 131224 80532 143166 80560
rect 130470 80384 130476 80436
rect 130528 80424 130534 80436
rect 130528 80396 141418 80424
rect 130528 80384 130534 80396
rect 130378 80316 130384 80368
rect 130436 80356 130442 80368
rect 130436 80328 140084 80356
rect 130436 80316 130442 80328
rect 128998 80044 129004 80096
rect 129056 80084 129062 80096
rect 129056 80056 134058 80084
rect 129056 80044 129062 80056
rect 132540 79908 132546 79960
rect 132598 79908 132604 79960
rect 132724 79948 132730 79960
rect 132696 79908 132730 79948
rect 132782 79908 132788 79960
rect 132816 79908 132822 79960
rect 132874 79908 132880 79960
rect 132908 79908 132914 79960
rect 132966 79908 132972 79960
rect 133000 79908 133006 79960
rect 133058 79908 133064 79960
rect 133368 79948 133374 79960
rect 133340 79908 133374 79948
rect 133426 79908 133432 79960
rect 133460 79908 133466 79960
rect 133518 79908 133524 79960
rect 132558 79824 132586 79908
rect 132494 79772 132500 79824
rect 132552 79784 132586 79824
rect 132552 79772 132558 79784
rect 113726 79636 113732 79688
rect 113784 79676 113790 79688
rect 130378 79676 130384 79688
rect 113784 79648 130384 79676
rect 113784 79636 113790 79648
rect 130378 79636 130384 79648
rect 130436 79636 130442 79688
rect 132696 79620 132724 79908
rect 132834 79880 132862 79908
rect 132788 79852 132862 79880
rect 132788 79756 132816 79852
rect 132926 79812 132954 79908
rect 132880 79784 132954 79812
rect 132880 79756 132908 79784
rect 133018 79756 133046 79908
rect 133092 79840 133098 79892
rect 133150 79880 133156 79892
rect 133150 79840 133184 79880
rect 133156 79756 133184 79840
rect 132770 79704 132776 79756
rect 132828 79704 132834 79756
rect 132862 79704 132868 79756
rect 132920 79704 132926 79756
rect 132954 79704 132960 79756
rect 133012 79716 133046 79756
rect 133012 79704 133018 79716
rect 133138 79704 133144 79756
rect 133196 79704 133202 79756
rect 133340 79688 133368 79908
rect 133478 79880 133506 79908
rect 134030 79892 134058 80056
rect 138308 80056 139302 80084
rect 135272 79988 136082 80016
rect 134380 79908 134386 79960
rect 134438 79908 134444 79960
rect 134564 79908 134570 79960
rect 134622 79908 134628 79960
rect 135024 79948 135030 79960
rect 134950 79920 135030 79948
rect 133478 79852 133644 79880
rect 133322 79636 133328 79688
rect 133380 79636 133386 79688
rect 133616 79676 133644 79852
rect 133736 79840 133742 79892
rect 133794 79840 133800 79892
rect 133828 79840 133834 79892
rect 133886 79840 133892 79892
rect 133920 79840 133926 79892
rect 133978 79840 133984 79892
rect 134012 79840 134018 79892
rect 134070 79840 134076 79892
rect 134398 79880 134426 79908
rect 134260 79852 134426 79880
rect 133616 79648 133690 79676
rect 109862 79568 109868 79620
rect 109920 79608 109926 79620
rect 130286 79608 130292 79620
rect 109920 79580 130292 79608
rect 109920 79568 109926 79580
rect 130286 79568 130292 79580
rect 130344 79568 130350 79620
rect 132678 79568 132684 79620
rect 132736 79568 132742 79620
rect 119246 79500 119252 79552
rect 119304 79540 119310 79552
rect 130562 79540 130568 79552
rect 119304 79512 130568 79540
rect 119304 79500 119310 79512
rect 130562 79500 130568 79512
rect 130620 79540 130626 79552
rect 130620 79512 132724 79540
rect 130620 79500 130626 79512
rect 111150 79432 111156 79484
rect 111208 79472 111214 79484
rect 131022 79472 131028 79484
rect 111208 79444 131028 79472
rect 111208 79432 111214 79444
rect 131022 79432 131028 79444
rect 131080 79432 131086 79484
rect 108206 79364 108212 79416
rect 108264 79404 108270 79416
rect 129918 79404 129924 79416
rect 108264 79376 129924 79404
rect 108264 79364 108270 79376
rect 129918 79364 129924 79376
rect 129976 79364 129982 79416
rect 132696 79404 132724 79512
rect 132862 79432 132868 79484
rect 132920 79472 132926 79484
rect 133662 79472 133690 79648
rect 133754 79608 133782 79840
rect 133846 79756 133874 79840
rect 133938 79812 133966 79840
rect 133938 79784 134104 79812
rect 133846 79716 133880 79756
rect 133874 79704 133880 79716
rect 133932 79704 133938 79756
rect 134076 79688 134104 79784
rect 134260 79688 134288 79852
rect 134472 79840 134478 79892
rect 134530 79840 134536 79892
rect 134490 79812 134518 79840
rect 134352 79784 134518 79812
rect 134352 79688 134380 79784
rect 134582 79756 134610 79908
rect 134518 79704 134524 79756
rect 134576 79716 134610 79756
rect 134576 79704 134582 79716
rect 134058 79636 134064 79688
rect 134116 79636 134122 79688
rect 134242 79636 134248 79688
rect 134300 79636 134306 79688
rect 134334 79636 134340 79688
rect 134392 79636 134398 79688
rect 133754 79580 134012 79608
rect 133984 79552 134012 79580
rect 133966 79500 133972 79552
rect 134024 79500 134030 79552
rect 134702 79500 134708 79552
rect 134760 79540 134766 79552
rect 134950 79540 134978 79920
rect 135024 79908 135030 79920
rect 135082 79908 135088 79960
rect 135116 79908 135122 79960
rect 135174 79908 135180 79960
rect 135134 79756 135162 79908
rect 135070 79704 135076 79756
rect 135128 79716 135162 79756
rect 135128 79704 135134 79716
rect 135272 79620 135300 79988
rect 136054 79960 136082 79988
rect 135392 79908 135398 79960
rect 135450 79908 135456 79960
rect 135576 79908 135582 79960
rect 135634 79908 135640 79960
rect 135760 79908 135766 79960
rect 135818 79908 135824 79960
rect 135852 79908 135858 79960
rect 135910 79908 135916 79960
rect 136036 79908 136042 79960
rect 136094 79908 136100 79960
rect 136404 79908 136410 79960
rect 136462 79908 136468 79960
rect 136588 79908 136594 79960
rect 136646 79908 136652 79960
rect 136772 79948 136778 79960
rect 136744 79908 136778 79948
rect 136830 79908 136836 79960
rect 137140 79908 137146 79960
rect 137198 79908 137204 79960
rect 137232 79908 137238 79960
rect 137290 79908 137296 79960
rect 137416 79908 137422 79960
rect 137474 79908 137480 79960
rect 137508 79908 137514 79960
rect 137566 79908 137572 79960
rect 138060 79948 138066 79960
rect 137894 79920 138066 79948
rect 135254 79568 135260 79620
rect 135312 79568 135318 79620
rect 135410 79552 135438 79908
rect 135594 79676 135622 79908
rect 135778 79824 135806 79908
rect 135714 79772 135720 79824
rect 135772 79784 135806 79824
rect 135772 79772 135778 79784
rect 135870 79756 135898 79908
rect 136312 79772 136318 79824
rect 136370 79772 136376 79824
rect 135806 79704 135812 79756
rect 135864 79716 135898 79756
rect 135864 79704 135870 79716
rect 136330 79676 136358 79772
rect 135594 79648 135668 79676
rect 135640 79552 135668 79648
rect 135824 79648 136358 79676
rect 134760 79512 134978 79540
rect 134760 79500 134766 79512
rect 135346 79500 135352 79552
rect 135404 79512 135438 79552
rect 135404 79500 135410 79512
rect 135622 79500 135628 79552
rect 135680 79500 135686 79552
rect 135824 79540 135852 79648
rect 135898 79568 135904 79620
rect 135956 79608 135962 79620
rect 136422 79608 136450 79908
rect 136606 79688 136634 79908
rect 136744 79688 136772 79908
rect 136956 79880 136962 79892
rect 136836 79852 136962 79880
rect 136542 79636 136548 79688
rect 136600 79648 136634 79688
rect 136600 79636 136606 79648
rect 136726 79636 136732 79688
rect 136784 79636 136790 79688
rect 136836 79620 136864 79852
rect 136956 79840 136962 79852
rect 137014 79840 137020 79892
rect 137158 79812 137186 79908
rect 137020 79784 137186 79812
rect 137020 79676 137048 79784
rect 137094 79704 137100 79756
rect 137152 79744 137158 79756
rect 137250 79744 137278 79908
rect 137434 79824 137462 79908
rect 137370 79772 137376 79824
rect 137428 79784 137462 79824
rect 137428 79772 137434 79784
rect 137526 79756 137554 79908
rect 137600 79840 137606 79892
rect 137658 79840 137664 79892
rect 137152 79716 137278 79744
rect 137152 79704 137158 79716
rect 137462 79704 137468 79756
rect 137520 79716 137554 79756
rect 137520 79704 137526 79716
rect 137186 79676 137192 79688
rect 137020 79648 137192 79676
rect 137186 79636 137192 79648
rect 137244 79636 137250 79688
rect 137618 79620 137646 79840
rect 137894 79756 137922 79920
rect 138060 79908 138066 79920
rect 138118 79908 138124 79960
rect 138152 79908 138158 79960
rect 138210 79908 138216 79960
rect 137968 79840 137974 79892
rect 138026 79880 138032 79892
rect 138026 79852 138106 79880
rect 138026 79840 138032 79852
rect 137894 79716 137928 79756
rect 137922 79704 137928 79716
rect 137980 79704 137986 79756
rect 138078 79688 138106 79852
rect 138014 79636 138020 79688
rect 138072 79648 138106 79688
rect 138072 79636 138078 79648
rect 138170 79620 138198 79908
rect 138308 79688 138336 80056
rect 139274 79960 139302 80056
rect 140056 80016 140084 80328
rect 141390 80084 141418 80396
rect 143138 80152 143166 80532
rect 143322 80220 143350 80600
rect 143506 80288 143534 80872
rect 144610 80628 144638 80940
rect 145806 80696 145834 81008
rect 154546 80900 154574 81144
rect 153350 80872 154574 80900
rect 145806 80668 145880 80696
rect 145852 80628 145880 80668
rect 144610 80600 145788 80628
rect 145852 80600 146938 80628
rect 145760 80560 145788 80600
rect 145760 80532 146110 80560
rect 143506 80260 145604 80288
rect 143322 80192 144960 80220
rect 143138 80124 144546 80152
rect 141390 80056 144454 80084
rect 140056 79988 141878 80016
rect 138612 79948 138618 79960
rect 138492 79920 138618 79948
rect 138290 79636 138296 79688
rect 138348 79636 138354 79688
rect 138492 79676 138520 79920
rect 138612 79908 138618 79920
rect 138670 79908 138676 79960
rect 138704 79908 138710 79960
rect 138762 79908 138768 79960
rect 138796 79908 138802 79960
rect 138854 79908 138860 79960
rect 139256 79908 139262 79960
rect 139314 79908 139320 79960
rect 139348 79908 139354 79960
rect 139406 79908 139412 79960
rect 139532 79908 139538 79960
rect 139590 79908 139596 79960
rect 139624 79908 139630 79960
rect 139682 79908 139688 79960
rect 139808 79908 139814 79960
rect 139866 79908 139872 79960
rect 139900 79908 139906 79960
rect 139958 79908 139964 79960
rect 140084 79908 140090 79960
rect 140142 79908 140148 79960
rect 140176 79908 140182 79960
rect 140234 79908 140240 79960
rect 140360 79908 140366 79960
rect 140418 79908 140424 79960
rect 140544 79908 140550 79960
rect 140602 79948 140608 79960
rect 140602 79920 140820 79948
rect 140602 79908 140608 79920
rect 138722 79880 138750 79908
rect 138584 79852 138750 79880
rect 138584 79824 138612 79852
rect 138814 79824 138842 79908
rect 139072 79880 139078 79892
rect 138566 79772 138572 79824
rect 138624 79772 138630 79824
rect 138750 79772 138756 79824
rect 138808 79784 138842 79824
rect 139044 79840 139078 79880
rect 139130 79840 139136 79892
rect 138808 79772 138814 79784
rect 139044 79756 139072 79840
rect 139026 79704 139032 79756
rect 139084 79704 139090 79756
rect 139118 79704 139124 79756
rect 139176 79744 139182 79756
rect 139366 79744 139394 79908
rect 139550 79812 139578 79908
rect 139642 79880 139670 79908
rect 139642 79852 139716 79880
rect 139550 79784 139624 79812
rect 139596 79756 139624 79784
rect 139176 79716 139394 79744
rect 139176 79704 139182 79716
rect 139578 79704 139584 79756
rect 139636 79704 139642 79756
rect 138566 79676 138572 79688
rect 138492 79648 138572 79676
rect 138566 79636 138572 79648
rect 138624 79636 138630 79688
rect 138658 79636 138664 79688
rect 138716 79676 138722 79688
rect 139688 79676 139716 79852
rect 139826 79756 139854 79908
rect 139762 79704 139768 79756
rect 139820 79716 139854 79756
rect 139820 79704 139826 79716
rect 138716 79648 139716 79676
rect 138716 79636 138722 79648
rect 135956 79580 136450 79608
rect 135956 79568 135962 79580
rect 136818 79568 136824 79620
rect 136876 79568 136882 79620
rect 137618 79580 137652 79620
rect 137646 79568 137652 79580
rect 137704 79568 137710 79620
rect 138170 79580 138204 79620
rect 138198 79568 138204 79580
rect 138256 79568 138262 79620
rect 139918 79608 139946 79908
rect 140102 79812 140130 79908
rect 140056 79784 140130 79812
rect 140056 79688 140084 79784
rect 140194 79756 140222 79908
rect 140130 79704 140136 79756
rect 140188 79716 140222 79756
rect 140188 79704 140194 79716
rect 140378 79688 140406 79908
rect 140038 79636 140044 79688
rect 140096 79636 140102 79688
rect 140378 79648 140412 79688
rect 140406 79636 140412 79648
rect 140464 79636 140470 79688
rect 140792 79620 140820 79920
rect 140884 79920 141326 79948
rect 140884 79620 140912 79920
rect 141298 79892 141326 79920
rect 141004 79880 141010 79892
rect 140976 79840 141010 79880
rect 141062 79840 141068 79892
rect 141280 79840 141286 79892
rect 141338 79840 141344 79892
rect 141464 79840 141470 79892
rect 141522 79840 141528 79892
rect 141740 79840 141746 79892
rect 141798 79840 141804 79892
rect 140314 79608 140320 79620
rect 139918 79580 140320 79608
rect 140314 79568 140320 79580
rect 140372 79568 140378 79620
rect 140774 79568 140780 79620
rect 140832 79568 140838 79620
rect 140866 79568 140872 79620
rect 140924 79568 140930 79620
rect 136358 79540 136364 79552
rect 135824 79512 136364 79540
rect 136358 79500 136364 79512
rect 136416 79500 136422 79552
rect 136910 79500 136916 79552
rect 136968 79540 136974 79552
rect 138106 79540 138112 79552
rect 136968 79512 138112 79540
rect 136968 79500 136974 79512
rect 138106 79500 138112 79512
rect 138164 79500 138170 79552
rect 140222 79500 140228 79552
rect 140280 79500 140286 79552
rect 132920 79444 133690 79472
rect 132920 79432 132926 79444
rect 133874 79432 133880 79484
rect 133932 79472 133938 79484
rect 140240 79472 140268 79500
rect 133932 79444 140268 79472
rect 140976 79472 141004 79840
rect 141482 79744 141510 79840
rect 141068 79716 141510 79744
rect 141068 79552 141096 79716
rect 141326 79568 141332 79620
rect 141384 79568 141390 79620
rect 141418 79568 141424 79620
rect 141476 79608 141482 79620
rect 141758 79608 141786 79840
rect 141476 79580 141786 79608
rect 141476 79568 141482 79580
rect 141050 79500 141056 79552
rect 141108 79500 141114 79552
rect 141344 79484 141372 79568
rect 141234 79472 141240 79484
rect 140976 79444 141240 79472
rect 133932 79432 133938 79444
rect 141234 79432 141240 79444
rect 141292 79432 141298 79484
rect 141326 79432 141332 79484
rect 141384 79432 141390 79484
rect 139670 79404 139676 79416
rect 132696 79376 139676 79404
rect 139670 79364 139676 79376
rect 139728 79364 139734 79416
rect 140222 79364 140228 79416
rect 140280 79404 140286 79416
rect 140498 79404 140504 79416
rect 140280 79376 140504 79404
rect 140280 79364 140286 79376
rect 140498 79364 140504 79376
rect 140556 79364 140562 79416
rect 141850 79404 141878 79988
rect 142016 79908 142022 79960
rect 142074 79908 142080 79960
rect 142476 79908 142482 79960
rect 142534 79908 142540 79960
rect 142844 79948 142850 79960
rect 142632 79920 142850 79948
rect 142034 79484 142062 79908
rect 142200 79840 142206 79892
rect 142258 79840 142264 79892
rect 142384 79840 142390 79892
rect 142442 79840 142448 79892
rect 142218 79688 142246 79840
rect 142402 79756 142430 79840
rect 142338 79704 142344 79756
rect 142396 79716 142430 79756
rect 142396 79704 142402 79716
rect 142154 79636 142160 79688
rect 142212 79648 142246 79688
rect 142212 79636 142218 79648
rect 142246 79568 142252 79620
rect 142304 79608 142310 79620
rect 142494 79608 142522 79908
rect 142632 79620 142660 79920
rect 142844 79908 142850 79920
rect 142902 79908 142908 79960
rect 143304 79948 143310 79960
rect 143276 79908 143310 79948
rect 143362 79908 143368 79960
rect 143276 79620 143304 79908
rect 142304 79580 142522 79608
rect 142304 79568 142310 79580
rect 142614 79568 142620 79620
rect 142672 79568 142678 79620
rect 143258 79568 143264 79620
rect 143316 79568 143322 79620
rect 143598 79608 143626 80056
rect 143690 79988 143902 80016
rect 143690 79676 143718 79988
rect 143874 79960 143902 79988
rect 144426 79960 144454 80056
rect 144518 80016 144546 80124
rect 144932 80084 144960 80192
rect 145576 80152 145604 80260
rect 145576 80124 145650 80152
rect 144932 80056 145282 80084
rect 144518 79988 145006 80016
rect 143856 79908 143862 79960
rect 143914 79908 143920 79960
rect 144040 79908 144046 79960
rect 144098 79908 144104 79960
rect 144316 79908 144322 79960
rect 144374 79908 144380 79960
rect 144408 79908 144414 79960
rect 144466 79908 144472 79960
rect 144500 79908 144506 79960
rect 144558 79908 144564 79960
rect 144592 79908 144598 79960
rect 144650 79908 144656 79960
rect 144684 79908 144690 79960
rect 144742 79908 144748 79960
rect 144868 79948 144874 79960
rect 144840 79908 144874 79948
rect 144926 79908 144932 79960
rect 144058 79824 144086 79908
rect 144132 79840 144138 79892
rect 144190 79840 144196 79892
rect 144040 79772 144046 79824
rect 144098 79772 144104 79824
rect 143902 79676 143908 79688
rect 143690 79648 143908 79676
rect 143902 79636 143908 79648
rect 143960 79636 143966 79688
rect 143810 79608 143816 79620
rect 143598 79580 143816 79608
rect 143810 79568 143816 79580
rect 143868 79568 143874 79620
rect 143994 79568 144000 79620
rect 144052 79608 144058 79620
rect 144150 79608 144178 79840
rect 144334 79824 144362 79908
rect 144518 79824 144546 79908
rect 144334 79784 144368 79824
rect 144362 79772 144368 79784
rect 144420 79772 144426 79824
rect 144454 79772 144460 79824
rect 144512 79784 144546 79824
rect 144512 79772 144518 79784
rect 144610 79688 144638 79908
rect 144546 79636 144552 79688
rect 144604 79648 144638 79688
rect 144604 79636 144610 79648
rect 144702 79620 144730 79908
rect 144052 79580 144178 79608
rect 144052 79568 144058 79580
rect 144638 79568 144644 79620
rect 144696 79580 144730 79620
rect 144696 79568 144702 79580
rect 142798 79500 142804 79552
rect 142856 79540 142862 79552
rect 143074 79540 143080 79552
rect 142856 79512 143080 79540
rect 142856 79500 142862 79512
rect 143074 79500 143080 79512
rect 143132 79500 143138 79552
rect 144178 79500 144184 79552
rect 144236 79540 144242 79552
rect 144840 79540 144868 79908
rect 144978 79880 145006 79988
rect 144932 79852 145006 79880
rect 144932 79620 144960 79852
rect 144914 79568 144920 79620
rect 144972 79568 144978 79620
rect 144236 79512 144868 79540
rect 144236 79500 144242 79512
rect 141970 79432 141976 79484
rect 142028 79444 142062 79484
rect 145254 79472 145282 80056
rect 145622 80016 145650 80124
rect 145530 79988 145650 80016
rect 145530 79892 145558 79988
rect 146082 79960 146110 80532
rect 146064 79908 146070 79960
rect 146122 79908 146128 79960
rect 146248 79908 146254 79960
rect 146306 79908 146312 79960
rect 146340 79908 146346 79960
rect 146398 79908 146404 79960
rect 146524 79908 146530 79960
rect 146582 79908 146588 79960
rect 146616 79908 146622 79960
rect 146674 79948 146680 79960
rect 146674 79908 146708 79948
rect 145328 79840 145334 79892
rect 145386 79840 145392 79892
rect 145512 79840 145518 79892
rect 145570 79840 145576 79892
rect 145604 79840 145610 79892
rect 145662 79880 145668 79892
rect 145662 79840 145696 79880
rect 145346 79540 145374 79840
rect 145530 79756 145558 79840
rect 145530 79716 145564 79756
rect 145558 79704 145564 79716
rect 145616 79704 145622 79756
rect 145668 79608 145696 79840
rect 146064 79772 146070 79824
rect 146122 79772 146128 79824
rect 145926 79636 145932 79688
rect 145984 79676 145990 79688
rect 146082 79676 146110 79772
rect 146266 79756 146294 79908
rect 146202 79704 146208 79756
rect 146260 79716 146294 79756
rect 146260 79704 146266 79716
rect 145984 79648 146110 79676
rect 145984 79636 145990 79648
rect 146358 79620 146386 79908
rect 146432 79840 146438 79892
rect 146490 79840 146496 79892
rect 146018 79608 146024 79620
rect 145668 79580 146024 79608
rect 146018 79568 146024 79580
rect 146076 79568 146082 79620
rect 146294 79568 146300 79620
rect 146352 79580 146386 79620
rect 146352 79568 146358 79580
rect 146450 79552 146478 79840
rect 146542 79756 146570 79908
rect 146542 79716 146576 79756
rect 146570 79704 146576 79716
rect 146628 79704 146634 79756
rect 145650 79540 145656 79552
rect 145346 79512 145656 79540
rect 145650 79500 145656 79512
rect 145708 79500 145714 79552
rect 146450 79540 146484 79552
rect 146220 79512 146484 79540
rect 146220 79472 146248 79512
rect 146478 79500 146484 79512
rect 146536 79540 146542 79552
rect 146536 79512 146583 79540
rect 146536 79500 146542 79512
rect 145254 79444 146248 79472
rect 142028 79432 142034 79444
rect 146294 79432 146300 79484
rect 146352 79472 146358 79484
rect 146680 79472 146708 79908
rect 146910 79892 146938 80600
rect 153350 80220 153378 80872
rect 159514 80288 159542 81212
rect 164206 81172 164234 81212
rect 164206 81144 165614 81172
rect 165586 80968 165614 81144
rect 167748 81036 167776 81280
rect 182146 81144 187096 81172
rect 182146 81036 182174 81144
rect 186958 81104 186964 81116
rect 167748 81008 182174 81036
rect 186424 81076 186964 81104
rect 186424 80968 186452 81076
rect 186958 81064 186964 81076
rect 187016 81064 187022 81116
rect 187068 81036 187096 81144
rect 187326 81064 187332 81116
rect 187384 81104 187390 81116
rect 195146 81104 195152 81116
rect 187384 81076 195152 81104
rect 187384 81064 187390 81076
rect 195146 81064 195152 81076
rect 195204 81064 195210 81116
rect 214558 81064 214564 81116
rect 214616 81104 214622 81116
rect 214834 81104 214840 81116
rect 214616 81076 214840 81104
rect 214616 81064 214622 81076
rect 214834 81064 214840 81076
rect 214892 81064 214898 81116
rect 187068 81008 191834 81036
rect 165586 80940 166994 80968
rect 166966 80900 166994 80940
rect 169726 80940 171134 80968
rect 164206 80872 165614 80900
rect 166966 80872 168374 80900
rect 164206 80492 164234 80872
rect 165586 80696 165614 80872
rect 168346 80832 168374 80872
rect 169726 80832 169754 80940
rect 171106 80900 171134 80940
rect 172486 80940 175274 80968
rect 172486 80900 172514 80940
rect 171106 80872 172514 80900
rect 168346 80804 169754 80832
rect 175246 80832 175274 80940
rect 177776 80940 186452 80968
rect 177776 80832 177804 80940
rect 186682 80860 186688 80912
rect 186740 80900 186746 80912
rect 191806 80900 191834 81008
rect 215846 80900 215852 80912
rect 186740 80872 187280 80900
rect 191806 80872 215852 80900
rect 186740 80860 186746 80872
rect 175246 80804 177804 80832
rect 187252 80764 187280 80872
rect 215846 80860 215852 80872
rect 215904 80900 215910 80912
rect 234614 80900 234620 80912
rect 215904 80872 234620 80900
rect 215904 80860 215910 80872
rect 234614 80860 234620 80872
rect 234672 80860 234678 80912
rect 187510 80792 187516 80844
rect 187568 80832 187574 80844
rect 252554 80832 252560 80844
rect 187568 80804 252560 80832
rect 187568 80792 187574 80804
rect 252554 80792 252560 80804
rect 252612 80792 252618 80844
rect 187694 80764 187700 80776
rect 166966 80736 186452 80764
rect 187252 80736 187700 80764
rect 166966 80696 166994 80736
rect 165586 80668 166994 80696
rect 167196 80668 184244 80696
rect 153120 80192 153378 80220
rect 157444 80260 159542 80288
rect 160342 80464 164234 80492
rect 153120 80152 153148 80192
rect 150682 80124 153148 80152
rect 147002 79988 149008 80016
rect 147002 79960 147030 79988
rect 146984 79908 146990 79960
rect 147042 79908 147048 79960
rect 147278 79920 147490 79948
rect 146892 79840 146898 79892
rect 146950 79840 146956 79892
rect 147168 79840 147174 79892
rect 147226 79840 147232 79892
rect 146910 79540 146938 79840
rect 147186 79620 147214 79840
rect 147278 79676 147306 79920
rect 147462 79892 147490 79920
rect 147628 79908 147634 79960
rect 147686 79908 147692 79960
rect 148272 79908 148278 79960
rect 148330 79908 148336 79960
rect 148364 79908 148370 79960
rect 148422 79908 148428 79960
rect 147352 79840 147358 79892
rect 147410 79840 147416 79892
rect 147444 79840 147450 79892
rect 147502 79840 147508 79892
rect 147370 79744 147398 79840
rect 147646 79824 147674 79908
rect 147996 79840 148002 79892
rect 148054 79840 148060 79892
rect 147628 79772 147634 79824
rect 147686 79772 147692 79824
rect 148014 79744 148042 79840
rect 148290 79824 148318 79908
rect 148226 79772 148232 79824
rect 148284 79784 148318 79824
rect 148284 79772 148290 79784
rect 148382 79756 148410 79908
rect 148824 79772 148830 79824
rect 148882 79772 148888 79824
rect 147370 79716 147628 79744
rect 147278 79648 147536 79676
rect 147186 79580 147220 79620
rect 147214 79568 147220 79580
rect 147272 79568 147278 79620
rect 147398 79540 147404 79552
rect 146910 79512 147404 79540
rect 147398 79500 147404 79512
rect 147456 79500 147462 79552
rect 146352 79444 146708 79472
rect 146352 79432 146358 79444
rect 147030 79432 147036 79484
rect 147088 79472 147094 79484
rect 147508 79472 147536 79648
rect 147600 79552 147628 79716
rect 147830 79716 148042 79744
rect 147830 79552 147858 79716
rect 148318 79704 148324 79756
rect 148376 79716 148410 79756
rect 148376 79704 148382 79716
rect 148842 79608 148870 79772
rect 148842 79580 148916 79608
rect 147582 79500 147588 79552
rect 147640 79500 147646 79552
rect 147766 79500 147772 79552
rect 147824 79512 147858 79552
rect 147824 79500 147830 79512
rect 147088 79444 147536 79472
rect 147088 79432 147094 79444
rect 148318 79432 148324 79484
rect 148376 79472 148382 79484
rect 148778 79472 148784 79484
rect 148376 79444 148784 79472
rect 148376 79432 148382 79444
rect 148778 79432 148784 79444
rect 148836 79432 148842 79484
rect 147490 79404 147496 79416
rect 141850 79376 147496 79404
rect 147490 79364 147496 79376
rect 147548 79364 147554 79416
rect 148594 79364 148600 79416
rect 148652 79404 148658 79416
rect 148888 79404 148916 79580
rect 148980 79472 149008 79988
rect 150682 79960 150710 80124
rect 157444 80084 157472 80260
rect 153534 80056 154574 80084
rect 153534 80016 153562 80056
rect 153442 79988 153562 80016
rect 153442 79960 153470 79988
rect 149100 79908 149106 79960
rect 149158 79948 149164 79960
rect 149158 79908 149192 79948
rect 149284 79908 149290 79960
rect 149342 79908 149348 79960
rect 149744 79948 149750 79960
rect 149532 79920 149750 79948
rect 149164 79824 149192 79908
rect 149302 79880 149330 79908
rect 149256 79852 149330 79880
rect 149256 79824 149284 79852
rect 149146 79772 149152 79824
rect 149204 79772 149210 79824
rect 149238 79772 149244 79824
rect 149296 79772 149302 79824
rect 149532 79552 149560 79920
rect 149744 79908 149750 79920
rect 149802 79908 149808 79960
rect 150020 79948 150026 79960
rect 149992 79908 150026 79948
rect 150078 79908 150084 79960
rect 150388 79908 150394 79960
rect 150446 79908 150452 79960
rect 150664 79908 150670 79960
rect 150722 79908 150728 79960
rect 151492 79908 151498 79960
rect 151550 79908 151556 79960
rect 151676 79908 151682 79960
rect 151734 79908 151740 79960
rect 151768 79908 151774 79960
rect 151826 79908 151832 79960
rect 151952 79908 151958 79960
rect 152010 79908 152016 79960
rect 152044 79908 152050 79960
rect 152102 79908 152108 79960
rect 152228 79908 152234 79960
rect 152286 79948 152292 79960
rect 152286 79920 152550 79948
rect 152286 79908 152292 79920
rect 149652 79840 149658 79892
rect 149710 79840 149716 79892
rect 149836 79840 149842 79892
rect 149894 79880 149900 79892
rect 149894 79840 149928 79880
rect 149670 79608 149698 79840
rect 149900 79620 149928 79840
rect 149992 79620 150020 79908
rect 150112 79880 150118 79892
rect 150084 79840 150118 79880
rect 150170 79840 150176 79892
rect 149790 79608 149796 79620
rect 149670 79580 149796 79608
rect 149790 79568 149796 79580
rect 149848 79568 149854 79620
rect 149882 79568 149888 79620
rect 149940 79568 149946 79620
rect 149974 79568 149980 79620
rect 150032 79568 150038 79620
rect 150084 79552 150112 79840
rect 150406 79688 150434 79908
rect 150480 79840 150486 79892
rect 150538 79840 150544 79892
rect 151124 79880 151130 79892
rect 150636 79852 151130 79880
rect 150342 79636 150348 79688
rect 150400 79648 150434 79688
rect 150400 79636 150406 79648
rect 149514 79500 149520 79552
rect 149572 79500 149578 79552
rect 150066 79500 150072 79552
rect 150124 79500 150130 79552
rect 149698 79472 149704 79484
rect 148980 79444 149704 79472
rect 149698 79432 149704 79444
rect 149756 79432 149762 79484
rect 150498 79472 150526 79840
rect 150636 79824 150664 79852
rect 151124 79840 151130 79852
rect 151182 79840 151188 79892
rect 150618 79772 150624 79824
rect 150676 79772 150682 79824
rect 151510 79608 151538 79908
rect 151694 79688 151722 79908
rect 151630 79636 151636 79688
rect 151688 79648 151722 79688
rect 151786 79688 151814 79908
rect 151970 79824 151998 79908
rect 152062 79880 152090 79908
rect 152062 79852 152136 79880
rect 151970 79784 152004 79824
rect 151998 79772 152004 79784
rect 152056 79772 152062 79824
rect 151786 79648 151820 79688
rect 151688 79636 151694 79648
rect 151814 79636 151820 79648
rect 151872 79636 151878 79688
rect 152108 79620 152136 79852
rect 152320 79840 152326 79892
rect 152378 79840 152384 79892
rect 151510 79580 151768 79608
rect 151740 79484 151768 79580
rect 152090 79568 152096 79620
rect 152148 79568 152154 79620
rect 152338 79608 152366 79840
rect 152522 79744 152550 79920
rect 152596 79908 152602 79960
rect 152654 79908 152660 79960
rect 152872 79948 152878 79960
rect 152752 79920 152878 79948
rect 152614 79824 152642 79908
rect 152596 79772 152602 79824
rect 152654 79772 152660 79824
rect 152522 79716 152688 79744
rect 152660 79688 152688 79716
rect 152752 79688 152780 79920
rect 152872 79908 152878 79920
rect 152930 79908 152936 79960
rect 153240 79908 153246 79960
rect 153298 79908 153304 79960
rect 153424 79908 153430 79960
rect 153482 79908 153488 79960
rect 153516 79908 153522 79960
rect 153574 79948 153580 79960
rect 153574 79908 153608 79948
rect 153792 79908 153798 79960
rect 153850 79908 153856 79960
rect 153976 79908 153982 79960
rect 154034 79948 154040 79960
rect 154034 79920 154160 79948
rect 154034 79908 154040 79920
rect 152964 79880 152970 79892
rect 152844 79852 152970 79880
rect 152844 79688 152872 79852
rect 152964 79840 152970 79852
rect 153022 79840 153028 79892
rect 153258 79744 153286 79908
rect 153212 79716 153286 79744
rect 152642 79636 152648 79688
rect 152700 79636 152706 79688
rect 152734 79636 152740 79688
rect 152792 79636 152798 79688
rect 152826 79636 152832 79688
rect 152884 79636 152890 79688
rect 153102 79608 153108 79620
rect 152338 79580 153108 79608
rect 153102 79568 153108 79580
rect 153160 79568 153166 79620
rect 153212 79540 153240 79716
rect 153378 79636 153384 79688
rect 153436 79676 153442 79688
rect 153580 79676 153608 79908
rect 153700 79840 153706 79892
rect 153758 79840 153764 79892
rect 153718 79688 153746 79840
rect 153436 79648 153608 79676
rect 153436 79636 153442 79648
rect 153654 79636 153660 79688
rect 153712 79648 153746 79688
rect 153712 79636 153718 79648
rect 153810 79620 153838 79908
rect 153884 79840 153890 79892
rect 153942 79880 153948 79892
rect 153942 79840 153976 79880
rect 153948 79756 153976 79840
rect 153930 79704 153936 79756
rect 153988 79704 153994 79756
rect 153746 79568 153752 79620
rect 153804 79580 153838 79620
rect 153804 79568 153810 79580
rect 153654 79540 153660 79552
rect 153212 79512 153660 79540
rect 153654 79500 153660 79512
rect 153712 79500 153718 79552
rect 154132 79540 154160 79920
rect 154344 79908 154350 79960
rect 154402 79948 154408 79960
rect 154402 79908 154436 79948
rect 154298 79540 154304 79552
rect 154132 79512 154304 79540
rect 154298 79500 154304 79512
rect 154356 79500 154362 79552
rect 151446 79472 151452 79484
rect 150498 79444 151452 79472
rect 151446 79432 151452 79444
rect 151504 79432 151510 79484
rect 151722 79432 151728 79484
rect 151780 79432 151786 79484
rect 153286 79432 153292 79484
rect 153344 79472 153350 79484
rect 154408 79472 154436 79908
rect 154546 79880 154574 80056
rect 154822 80056 157472 80084
rect 154822 79960 154850 80056
rect 155098 79988 155310 80016
rect 155098 79960 155126 79988
rect 154804 79908 154810 79960
rect 154862 79908 154868 79960
rect 155080 79908 155086 79960
rect 155138 79908 155144 79960
rect 155172 79908 155178 79960
rect 155230 79908 155236 79960
rect 154546 79852 154850 79880
rect 154822 79824 154850 79852
rect 154896 79840 154902 79892
rect 154954 79840 154960 79892
rect 154712 79812 154718 79824
rect 153344 79444 154436 79472
rect 154592 79784 154718 79812
rect 154592 79472 154620 79784
rect 154712 79772 154718 79784
rect 154770 79772 154776 79824
rect 154804 79772 154810 79824
rect 154862 79772 154868 79824
rect 154914 79756 154942 79840
rect 154914 79716 154948 79756
rect 154942 79704 154948 79716
rect 155000 79704 155006 79756
rect 155190 79676 155218 79908
rect 154684 79648 155218 79676
rect 154684 79620 154712 79648
rect 154666 79568 154672 79620
rect 154724 79568 154730 79620
rect 154758 79568 154764 79620
rect 154816 79608 154822 79620
rect 155282 79608 155310 79988
rect 156018 79988 156230 80016
rect 155448 79908 155454 79960
rect 155506 79908 155512 79960
rect 155632 79908 155638 79960
rect 155690 79908 155696 79960
rect 155466 79880 155494 79908
rect 155466 79852 155540 79880
rect 155512 79824 155540 79852
rect 155650 79824 155678 79908
rect 155724 79840 155730 79892
rect 155782 79840 155788 79892
rect 155816 79840 155822 79892
rect 155874 79880 155880 79892
rect 155874 79852 155954 79880
rect 155874 79840 155880 79852
rect 155494 79772 155500 79824
rect 155552 79772 155558 79824
rect 155586 79772 155592 79824
rect 155644 79784 155678 79824
rect 155644 79772 155650 79784
rect 155742 79756 155770 79840
rect 155742 79716 155776 79756
rect 155770 79704 155776 79716
rect 155828 79704 155834 79756
rect 154816 79580 155310 79608
rect 154816 79568 154822 79580
rect 155926 79484 155954 79852
rect 156018 79552 156046 79988
rect 156202 79960 156230 79988
rect 156184 79908 156190 79960
rect 156242 79908 156248 79960
rect 156368 79908 156374 79960
rect 156426 79908 156432 79960
rect 156828 79908 156834 79960
rect 156886 79948 156892 79960
rect 157380 79948 157386 79960
rect 156886 79920 157058 79948
rect 156886 79908 156892 79920
rect 156386 79880 156414 79908
rect 156248 79852 156414 79880
rect 156248 79688 156276 79852
rect 156460 79840 156466 79892
rect 156518 79840 156524 79892
rect 156644 79840 156650 79892
rect 156702 79840 156708 79892
rect 156920 79840 156926 79892
rect 156978 79840 156984 79892
rect 156230 79636 156236 79688
rect 156288 79636 156294 79688
rect 156018 79512 156052 79552
rect 156046 79500 156052 79512
rect 156104 79500 156110 79552
rect 156138 79500 156144 79552
rect 156196 79540 156202 79552
rect 156478 79540 156506 79840
rect 156662 79620 156690 79840
rect 156598 79568 156604 79620
rect 156656 79580 156690 79620
rect 156656 79568 156662 79580
rect 156782 79568 156788 79620
rect 156840 79608 156846 79620
rect 156938 79608 156966 79840
rect 156840 79580 156966 79608
rect 156840 79568 156846 79580
rect 156196 79512 156506 79540
rect 156196 79500 156202 79512
rect 157030 79484 157058 79920
rect 157352 79908 157386 79948
rect 157438 79908 157444 79960
rect 157656 79908 157662 79960
rect 157714 79948 157720 79960
rect 157714 79920 157886 79948
rect 157714 79908 157720 79920
rect 157196 79772 157202 79824
rect 157254 79812 157260 79824
rect 157254 79772 157288 79812
rect 157260 79688 157288 79772
rect 157352 79688 157380 79908
rect 157748 79880 157754 79892
rect 157720 79840 157754 79880
rect 157806 79840 157812 79892
rect 157720 79756 157748 79840
rect 157702 79704 157708 79756
rect 157760 79704 157766 79756
rect 157242 79636 157248 79688
rect 157300 79636 157306 79688
rect 157334 79636 157340 79688
rect 157392 79636 157398 79688
rect 157610 79636 157616 79688
rect 157668 79676 157674 79688
rect 157858 79676 157886 79920
rect 157932 79908 157938 79960
rect 157990 79908 157996 79960
rect 158024 79908 158030 79960
rect 158082 79948 158088 79960
rect 158082 79908 158116 79948
rect 158208 79908 158214 79960
rect 158266 79908 158272 79960
rect 158392 79908 158398 79960
rect 158450 79908 158456 79960
rect 158484 79908 158490 79960
rect 158542 79908 158548 79960
rect 159220 79948 159226 79960
rect 159100 79920 159226 79948
rect 157950 79756 157978 79908
rect 158088 79756 158116 79908
rect 158226 79880 158254 79908
rect 158226 79852 158300 79880
rect 158162 79772 158168 79824
rect 158220 79772 158226 79824
rect 157950 79716 157984 79756
rect 157978 79704 157984 79716
rect 158036 79704 158042 79756
rect 158070 79704 158076 79756
rect 158128 79704 158134 79756
rect 158180 79688 158208 79772
rect 158272 79688 158300 79852
rect 157668 79648 157886 79676
rect 157668 79636 157674 79648
rect 158162 79636 158168 79688
rect 158220 79636 158226 79688
rect 158254 79636 158260 79688
rect 158312 79636 158318 79688
rect 157794 79500 157800 79552
rect 157852 79540 157858 79552
rect 158410 79540 158438 79908
rect 158502 79824 158530 79908
rect 158852 79840 158858 79892
rect 158910 79840 158916 79892
rect 158944 79840 158950 79892
rect 159002 79880 159008 79892
rect 159002 79840 159036 79880
rect 158502 79784 158536 79824
rect 158530 79772 158536 79784
rect 158588 79772 158594 79824
rect 158760 79772 158766 79824
rect 158818 79772 158824 79824
rect 158778 79608 158806 79772
rect 157852 79512 158438 79540
rect 158502 79580 158806 79608
rect 157852 79500 157858 79512
rect 158502 79484 158530 79580
rect 155126 79472 155132 79484
rect 154592 79444 155132 79472
rect 153344 79432 153350 79444
rect 155126 79432 155132 79444
rect 155184 79432 155190 79484
rect 155926 79444 155960 79484
rect 155954 79432 155960 79444
rect 156012 79432 156018 79484
rect 157030 79472 157064 79484
rect 156971 79444 157064 79472
rect 157058 79432 157064 79444
rect 157116 79472 157122 79484
rect 158346 79472 158352 79484
rect 157116 79444 158352 79472
rect 157116 79432 157122 79444
rect 158346 79432 158352 79444
rect 158404 79432 158410 79484
rect 158502 79444 158536 79484
rect 158530 79432 158536 79444
rect 158588 79432 158594 79484
rect 158714 79432 158720 79484
rect 158772 79472 158778 79484
rect 158870 79472 158898 79840
rect 159008 79620 159036 79840
rect 159100 79620 159128 79920
rect 159220 79908 159226 79920
rect 159278 79908 159284 79960
rect 159864 79908 159870 79960
rect 159922 79908 159928 79960
rect 159680 79840 159686 79892
rect 159738 79840 159744 79892
rect 159404 79772 159410 79824
rect 159462 79772 159468 79824
rect 159422 79744 159450 79772
rect 159376 79716 159450 79744
rect 158990 79568 158996 79620
rect 159048 79568 159054 79620
rect 159082 79568 159088 79620
rect 159140 79568 159146 79620
rect 158772 79444 158898 79472
rect 159376 79472 159404 79716
rect 159698 79676 159726 79840
rect 159468 79648 159726 79676
rect 159468 79552 159496 79648
rect 159450 79500 159456 79552
rect 159508 79500 159514 79552
rect 159882 79484 159910 79908
rect 160342 79824 160370 80464
rect 167196 80356 167224 80668
rect 182128 80628 182134 80640
rect 162688 80328 167224 80356
rect 167288 80600 182134 80628
rect 160434 79988 160922 80016
rect 160434 79960 160462 79988
rect 160416 79908 160422 79960
rect 160474 79908 160480 79960
rect 160508 79908 160514 79960
rect 160566 79908 160572 79960
rect 160600 79908 160606 79960
rect 160658 79948 160664 79960
rect 160658 79920 160830 79948
rect 160658 79908 160664 79920
rect 160342 79784 160376 79824
rect 160370 79772 160376 79784
rect 160428 79772 160434 79824
rect 160094 79568 160100 79620
rect 160152 79608 160158 79620
rect 160526 79608 160554 79908
rect 160692 79840 160698 79892
rect 160750 79840 160756 79892
rect 160152 79580 160554 79608
rect 160152 79568 160158 79580
rect 160554 79500 160560 79552
rect 160612 79540 160618 79552
rect 160710 79540 160738 79840
rect 160612 79512 160738 79540
rect 160612 79500 160618 79512
rect 159634 79472 159640 79484
rect 159376 79444 159640 79472
rect 158772 79432 158778 79444
rect 159634 79432 159640 79444
rect 159692 79432 159698 79484
rect 159818 79432 159824 79484
rect 159876 79444 159910 79484
rect 159876 79432 159882 79444
rect 160462 79432 160468 79484
rect 160520 79472 160526 79484
rect 160802 79472 160830 79920
rect 160520 79444 160830 79472
rect 160894 79484 160922 79988
rect 161152 79948 161158 79960
rect 160986 79920 161158 79948
rect 160986 79540 161014 79920
rect 161152 79908 161158 79920
rect 161210 79908 161216 79960
rect 161520 79908 161526 79960
rect 161578 79908 161584 79960
rect 161612 79908 161618 79960
rect 161670 79908 161676 79960
rect 161704 79908 161710 79960
rect 161762 79948 161768 79960
rect 161762 79920 162394 79948
rect 161762 79908 161768 79920
rect 161060 79840 161066 79892
rect 161118 79840 161124 79892
rect 161244 79840 161250 79892
rect 161302 79840 161308 79892
rect 161336 79840 161342 79892
rect 161394 79840 161400 79892
rect 161078 79688 161106 79840
rect 161078 79648 161112 79688
rect 161106 79636 161112 79648
rect 161164 79636 161170 79688
rect 161262 79608 161290 79840
rect 161354 79688 161382 79840
rect 161354 79648 161388 79688
rect 161382 79636 161388 79648
rect 161440 79636 161446 79688
rect 161538 79676 161566 79908
rect 161630 79756 161658 79908
rect 161888 79880 161894 79892
rect 161860 79840 161894 79880
rect 161946 79840 161952 79892
rect 161980 79840 161986 79892
rect 162038 79840 162044 79892
rect 161860 79756 161888 79840
rect 161630 79716 161664 79756
rect 161658 79704 161664 79716
rect 161716 79704 161722 79756
rect 161842 79704 161848 79756
rect 161900 79704 161906 79756
rect 161538 79648 161612 79676
rect 161474 79608 161480 79620
rect 161262 79580 161480 79608
rect 161474 79568 161480 79580
rect 161532 79568 161538 79620
rect 161198 79540 161204 79552
rect 160986 79512 161204 79540
rect 161198 79500 161204 79512
rect 161256 79500 161262 79552
rect 161584 79540 161612 79648
rect 161658 79568 161664 79620
rect 161716 79608 161722 79620
rect 161998 79608 162026 79840
rect 161716 79580 162026 79608
rect 161716 79568 161722 79580
rect 161750 79540 161756 79552
rect 161584 79512 161756 79540
rect 161750 79500 161756 79512
rect 161808 79500 161814 79552
rect 160894 79444 160928 79484
rect 160520 79432 160526 79444
rect 160922 79432 160928 79444
rect 160980 79432 160986 79484
rect 162366 79472 162394 79920
rect 162440 79908 162446 79960
rect 162498 79908 162504 79960
rect 162458 79688 162486 79908
rect 162458 79648 162492 79688
rect 162486 79636 162492 79648
rect 162544 79636 162550 79688
rect 162688 79552 162716 80328
rect 167288 80288 167316 80600
rect 182128 80588 182134 80600
rect 182186 80588 182192 80640
rect 178126 80560 178132 80572
rect 164206 80260 164786 80288
rect 164206 80016 164234 80260
rect 162872 79988 164234 80016
rect 162872 79620 162900 79988
rect 163360 79948 163366 79960
rect 163056 79920 163366 79948
rect 162854 79568 162860 79620
rect 162912 79568 162918 79620
rect 163056 79552 163084 79920
rect 163360 79908 163366 79920
rect 163418 79908 163424 79960
rect 164280 79908 164286 79960
rect 164338 79908 164344 79960
rect 164648 79948 164654 79960
rect 164390 79920 164654 79948
rect 163176 79840 163182 79892
rect 163234 79840 163240 79892
rect 163268 79840 163274 79892
rect 163326 79840 163332 79892
rect 163194 79552 163222 79840
rect 163286 79608 163314 79840
rect 164298 79824 164326 79908
rect 163544 79772 163550 79824
rect 163602 79772 163608 79824
rect 164280 79772 164286 79824
rect 164338 79772 164344 79824
rect 163562 79676 163590 79772
rect 163562 79648 164096 79676
rect 164068 79620 164096 79648
rect 163498 79608 163504 79620
rect 163286 79580 163504 79608
rect 163498 79568 163504 79580
rect 163556 79568 163562 79620
rect 164050 79568 164056 79620
rect 164108 79568 164114 79620
rect 162670 79500 162676 79552
rect 162728 79500 162734 79552
rect 163038 79500 163044 79552
rect 163096 79500 163102 79552
rect 163194 79512 163228 79552
rect 163222 79500 163228 79512
rect 163280 79500 163286 79552
rect 164234 79500 164240 79552
rect 164292 79540 164298 79552
rect 164390 79540 164418 79920
rect 164648 79908 164654 79920
rect 164706 79908 164712 79960
rect 164758 79880 164786 80260
rect 164850 80260 167316 80288
rect 169726 80532 172514 80560
rect 164850 79960 164878 80260
rect 169726 80152 169754 80532
rect 172486 80492 172514 80532
rect 173866 80532 178132 80560
rect 173866 80492 173894 80532
rect 178126 80520 178132 80532
rect 178184 80520 178190 80572
rect 172486 80464 173894 80492
rect 184216 80492 184244 80668
rect 186424 80628 186452 80736
rect 187694 80724 187700 80736
rect 187752 80764 187758 80776
rect 270494 80764 270500 80776
rect 187752 80736 270500 80764
rect 187752 80724 187758 80736
rect 270494 80724 270500 80736
rect 270552 80724 270558 80776
rect 186958 80656 186964 80708
rect 187016 80696 187022 80708
rect 189258 80696 189264 80708
rect 187016 80668 189264 80696
rect 187016 80656 187022 80668
rect 189258 80656 189264 80668
rect 189316 80696 189322 80708
rect 288434 80696 288440 80708
rect 189316 80668 288440 80696
rect 189316 80656 189322 80668
rect 288434 80656 288440 80668
rect 288492 80656 288498 80708
rect 186682 80628 186688 80640
rect 186424 80600 186688 80628
rect 186682 80588 186688 80600
rect 186740 80588 186746 80640
rect 184382 80520 184388 80572
rect 184440 80560 184446 80572
rect 187326 80560 187332 80572
rect 184440 80532 187332 80560
rect 184440 80520 184446 80532
rect 187326 80520 187332 80532
rect 187384 80520 187390 80572
rect 187510 80492 187516 80504
rect 184216 80464 187516 80492
rect 187510 80452 187516 80464
rect 187568 80452 187574 80504
rect 178586 80424 178592 80436
rect 172992 80396 178592 80424
rect 169542 80124 169754 80152
rect 171014 80260 171134 80288
rect 164942 80056 167454 80084
rect 164832 79908 164838 79960
rect 164890 79908 164896 79960
rect 164942 79880 164970 80056
rect 167426 80016 167454 80056
rect 169542 80016 169570 80124
rect 166322 79988 167362 80016
rect 167426 79988 169570 80016
rect 166322 79960 166350 79988
rect 165752 79908 165758 79960
rect 165810 79908 165816 79960
rect 165844 79908 165850 79960
rect 165902 79908 165908 79960
rect 165936 79908 165942 79960
rect 165994 79948 166000 79960
rect 165994 79920 166120 79948
rect 165994 79908 166000 79920
rect 164758 79852 164970 79880
rect 165384 79840 165390 79892
rect 165442 79840 165448 79892
rect 165568 79840 165574 79892
rect 165626 79840 165632 79892
rect 165770 79880 165798 79908
rect 165724 79852 165798 79880
rect 164602 79636 164608 79688
rect 164660 79676 164666 79688
rect 165402 79676 165430 79840
rect 164660 79648 165430 79676
rect 164660 79636 164666 79648
rect 165586 79608 165614 79840
rect 165724 79676 165752 79852
rect 165862 79756 165890 79908
rect 165798 79704 165804 79756
rect 165856 79716 165890 79756
rect 165856 79704 165862 79716
rect 165724 79648 165890 79676
rect 165706 79608 165712 79620
rect 165586 79580 165712 79608
rect 165706 79568 165712 79580
rect 165764 79568 165770 79620
rect 164292 79512 164418 79540
rect 165862 79540 165890 79648
rect 165982 79568 165988 79620
rect 166040 79608 166046 79620
rect 166092 79608 166120 79920
rect 166212 79908 166218 79960
rect 166270 79908 166276 79960
rect 166304 79908 166310 79960
rect 166362 79908 166368 79960
rect 166396 79908 166402 79960
rect 166454 79908 166460 79960
rect 166488 79908 166494 79960
rect 166546 79908 166552 79960
rect 166580 79908 166586 79960
rect 166638 79908 166644 79960
rect 167040 79908 167046 79960
rect 167098 79908 167104 79960
rect 166230 79756 166258 79908
rect 166414 79880 166442 79908
rect 166368 79852 166442 79880
rect 166230 79716 166264 79756
rect 166258 79704 166264 79716
rect 166316 79704 166322 79756
rect 166040 79580 166120 79608
rect 166040 79568 166046 79580
rect 166166 79540 166172 79552
rect 165862 79512 166172 79540
rect 164292 79500 164298 79512
rect 166166 79500 166172 79512
rect 166224 79500 166230 79552
rect 165246 79472 165252 79484
rect 162366 79444 165252 79472
rect 165246 79432 165252 79444
rect 165304 79432 165310 79484
rect 165614 79432 165620 79484
rect 165672 79472 165678 79484
rect 166368 79472 166396 79852
rect 166506 79812 166534 79908
rect 166460 79784 166534 79812
rect 166460 79540 166488 79784
rect 166598 79756 166626 79908
rect 166764 79772 166770 79824
rect 166822 79772 166828 79824
rect 166534 79704 166540 79756
rect 166592 79716 166626 79756
rect 166592 79704 166598 79716
rect 166782 79552 166810 79772
rect 166902 79704 166908 79756
rect 166960 79704 166966 79756
rect 166920 79552 166948 79704
rect 167058 79608 167086 79908
rect 167334 79688 167362 79988
rect 171014 79960 171042 80260
rect 167408 79908 167414 79960
rect 167466 79908 167472 79960
rect 168328 79908 168334 79960
rect 168386 79908 168392 79960
rect 168420 79908 168426 79960
rect 168478 79908 168484 79960
rect 168512 79908 168518 79960
rect 168570 79948 168576 79960
rect 169340 79948 169346 79960
rect 168570 79908 168604 79948
rect 167426 79744 167454 79908
rect 168346 79812 168374 79908
rect 168438 79880 168466 79908
rect 168438 79852 168512 79880
rect 168346 79784 168420 79812
rect 168282 79744 168288 79756
rect 167426 79716 168288 79744
rect 168282 79704 168288 79716
rect 168340 79704 168346 79756
rect 167334 79648 167368 79688
rect 167362 79636 167368 79648
rect 167420 79636 167426 79688
rect 167638 79608 167644 79620
rect 167058 79580 167644 79608
rect 167638 79568 167644 79580
rect 167696 79568 167702 79620
rect 166626 79540 166632 79552
rect 166460 79512 166632 79540
rect 166626 79500 166632 79512
rect 166684 79500 166690 79552
rect 166782 79512 166816 79552
rect 166810 79500 166816 79512
rect 166868 79500 166874 79552
rect 166902 79500 166908 79552
rect 166960 79500 166966 79552
rect 165672 79444 166396 79472
rect 165672 79432 165678 79444
rect 167730 79432 167736 79484
rect 167788 79472 167794 79484
rect 168392 79472 168420 79784
rect 168484 79688 168512 79852
rect 168576 79688 168604 79908
rect 168668 79920 169346 79948
rect 168466 79636 168472 79688
rect 168524 79636 168530 79688
rect 168558 79636 168564 79688
rect 168616 79636 168622 79688
rect 168668 79620 168696 79920
rect 169340 79908 169346 79920
rect 169398 79908 169404 79960
rect 169892 79948 169898 79960
rect 169864 79908 169898 79948
rect 169950 79908 169956 79960
rect 169984 79908 169990 79960
rect 170042 79908 170048 79960
rect 170076 79908 170082 79960
rect 170134 79908 170140 79960
rect 170444 79908 170450 79960
rect 170502 79908 170508 79960
rect 170904 79948 170910 79960
rect 170738 79920 170910 79948
rect 169064 79840 169070 79892
rect 169122 79840 169128 79892
rect 168788 79772 168794 79824
rect 168846 79772 168852 79824
rect 168806 79676 168834 79772
rect 168926 79676 168932 79688
rect 168806 79648 168932 79676
rect 168926 79636 168932 79648
rect 168984 79636 168990 79688
rect 168650 79568 168656 79620
rect 168708 79568 168714 79620
rect 167788 79444 168420 79472
rect 169082 79472 169110 79840
rect 169386 79744 169392 79756
rect 169220 79716 169392 79744
rect 169220 79620 169248 79716
rect 169386 79704 169392 79716
rect 169444 79704 169450 79756
rect 169202 79568 169208 79620
rect 169260 79568 169266 79620
rect 169864 79540 169892 79908
rect 170002 79880 170030 79908
rect 169956 79852 170030 79880
rect 169956 79756 169984 79852
rect 170094 79824 170122 79908
rect 170030 79772 170036 79824
rect 170088 79784 170122 79824
rect 170088 79772 170094 79784
rect 170260 79772 170266 79824
rect 170318 79772 170324 79824
rect 169938 79704 169944 79756
rect 169996 79704 170002 79756
rect 170278 79688 170306 79772
rect 170462 79756 170490 79908
rect 170462 79716 170496 79756
rect 170490 79704 170496 79716
rect 170548 79704 170554 79756
rect 170214 79636 170220 79688
rect 170272 79648 170306 79688
rect 170272 79636 170278 79648
rect 170738 79620 170766 79920
rect 170904 79908 170910 79920
rect 170962 79908 170968 79960
rect 170996 79908 171002 79960
rect 171054 79908 171060 79960
rect 170812 79840 170818 79892
rect 170870 79840 170876 79892
rect 170830 79676 170858 79840
rect 170950 79676 170956 79688
rect 170830 79648 170956 79676
rect 170950 79636 170956 79648
rect 171008 79636 171014 79688
rect 171106 79620 171134 80260
rect 172992 80152 173020 80396
rect 178586 80384 178592 80396
rect 178644 80384 178650 80436
rect 182174 80384 182180 80436
rect 182232 80424 182238 80436
rect 191098 80424 191104 80436
rect 182232 80396 191104 80424
rect 182232 80384 182238 80396
rect 191098 80384 191104 80396
rect 191156 80384 191162 80436
rect 177758 80248 177764 80300
rect 177816 80288 177822 80300
rect 177816 80260 180794 80288
rect 177816 80248 177822 80260
rect 179506 80220 179512 80232
rect 171934 80124 173020 80152
rect 173176 80192 179512 80220
rect 171934 79960 171962 80124
rect 173176 80084 173204 80192
rect 179506 80180 179512 80192
rect 179564 80180 179570 80232
rect 177758 80152 177764 80164
rect 172486 80056 173204 80084
rect 173314 80124 177764 80152
rect 171364 79908 171370 79960
rect 171422 79908 171428 79960
rect 171640 79908 171646 79960
rect 171698 79908 171704 79960
rect 171732 79908 171738 79960
rect 171790 79908 171796 79960
rect 171916 79908 171922 79960
rect 171974 79908 171980 79960
rect 172376 79908 172382 79960
rect 172434 79908 172440 79960
rect 171382 79880 171410 79908
rect 171336 79852 171410 79880
rect 171336 79824 171364 79852
rect 171318 79772 171324 79824
rect 171376 79772 171382 79824
rect 170738 79580 170772 79620
rect 170766 79568 170772 79580
rect 170824 79568 170830 79620
rect 171106 79580 171140 79620
rect 171134 79568 171140 79580
rect 171192 79568 171198 79620
rect 170582 79540 170588 79552
rect 169864 79512 170588 79540
rect 170582 79500 170588 79512
rect 170640 79500 170646 79552
rect 171658 79540 171686 79908
rect 171750 79620 171778 79908
rect 172008 79880 172014 79892
rect 171980 79840 172014 79880
rect 172066 79840 172072 79892
rect 171980 79620 172008 79840
rect 172394 79756 172422 79908
rect 172486 79824 172514 80056
rect 172578 79988 172974 80016
rect 172578 79960 172606 79988
rect 172560 79908 172566 79960
rect 172618 79908 172624 79960
rect 172652 79908 172658 79960
rect 172710 79908 172716 79960
rect 172744 79908 172750 79960
rect 172802 79908 172808 79960
rect 172486 79784 172520 79824
rect 172514 79772 172520 79784
rect 172572 79772 172578 79824
rect 172394 79716 172428 79756
rect 172422 79704 172428 79716
rect 172480 79704 172486 79756
rect 171750 79580 171784 79620
rect 171778 79568 171784 79580
rect 171836 79568 171842 79620
rect 171962 79568 171968 79620
rect 172020 79568 172026 79620
rect 172514 79568 172520 79620
rect 172572 79608 172578 79620
rect 172670 79608 172698 79908
rect 172762 79676 172790 79908
rect 172946 79744 172974 79988
rect 173314 79960 173342 80124
rect 177758 80112 177764 80124
rect 177816 80112 177822 80164
rect 178034 80084 178040 80096
rect 173498 80056 178040 80084
rect 173020 79908 173026 79960
rect 173078 79908 173084 79960
rect 173296 79908 173302 79960
rect 173354 79908 173360 79960
rect 173038 79880 173066 79908
rect 173498 79880 173526 80056
rect 178034 80044 178040 80056
rect 178092 80044 178098 80096
rect 178218 80016 178224 80028
rect 175246 79988 178224 80016
rect 175246 79960 175274 79988
rect 178218 79976 178224 79988
rect 178276 79976 178282 80028
rect 180766 80016 180794 80260
rect 201218 80084 201224 80096
rect 182146 80056 201224 80084
rect 182146 80016 182174 80056
rect 201218 80044 201224 80056
rect 201276 80084 201282 80096
rect 525794 80084 525800 80096
rect 201276 80056 525800 80084
rect 201276 80044 201282 80056
rect 525794 80044 525800 80056
rect 525852 80044 525858 80096
rect 180766 79988 182174 80016
rect 173572 79908 173578 79960
rect 173630 79908 173636 79960
rect 173940 79908 173946 79960
rect 173998 79948 174004 79960
rect 174768 79948 174774 79960
rect 173998 79920 174630 79948
rect 173998 79908 174004 79920
rect 173038 79852 173526 79880
rect 173388 79772 173394 79824
rect 173446 79772 173452 79824
rect 172946 79716 173204 79744
rect 173066 79676 173072 79688
rect 172762 79648 173072 79676
rect 173066 79636 173072 79648
rect 173124 79636 173130 79688
rect 173176 79620 173204 79716
rect 173406 79620 173434 79772
rect 172572 79580 172698 79608
rect 172572 79568 172578 79580
rect 173158 79568 173164 79620
rect 173216 79568 173222 79620
rect 173406 79580 173440 79620
rect 173434 79568 173440 79580
rect 173492 79568 173498 79620
rect 172146 79540 172152 79552
rect 171658 79512 172152 79540
rect 172146 79500 172152 79512
rect 172204 79500 172210 79552
rect 171870 79472 171876 79484
rect 169082 79444 171876 79472
rect 167788 79432 167794 79444
rect 171870 79432 171876 79444
rect 171928 79432 171934 79484
rect 172606 79432 172612 79484
rect 172664 79472 172670 79484
rect 173590 79472 173618 79908
rect 173756 79840 173762 79892
rect 173814 79840 173820 79892
rect 174216 79880 174222 79892
rect 174188 79840 174222 79880
rect 174274 79840 174280 79892
rect 174492 79880 174498 79892
rect 174464 79840 174498 79880
rect 174550 79840 174556 79892
rect 173774 79688 173802 79840
rect 173710 79636 173716 79688
rect 173768 79648 173802 79688
rect 173768 79636 173774 79648
rect 174188 79608 174216 79840
rect 172664 79444 173618 79472
rect 173820 79580 174216 79608
rect 173820 79472 173848 79580
rect 173894 79500 173900 79552
rect 173952 79540 173958 79552
rect 174464 79540 174492 79840
rect 174602 79620 174630 79920
rect 174538 79568 174544 79620
rect 174596 79580 174630 79620
rect 174740 79908 174774 79948
rect 174826 79908 174832 79960
rect 175044 79908 175050 79960
rect 175102 79908 175108 79960
rect 175136 79908 175142 79960
rect 175194 79908 175200 79960
rect 175228 79908 175234 79960
rect 175286 79908 175292 79960
rect 175412 79908 175418 79960
rect 175470 79908 175476 79960
rect 175504 79908 175510 79960
rect 175562 79908 175568 79960
rect 175964 79908 175970 79960
rect 176022 79908 176028 79960
rect 176976 79908 176982 79960
rect 177034 79908 177040 79960
rect 174740 79608 174768 79908
rect 174952 79880 174958 79892
rect 174832 79852 174958 79880
rect 174832 79756 174860 79852
rect 174952 79840 174958 79852
rect 175010 79840 175016 79892
rect 175062 79756 175090 79908
rect 174814 79704 174820 79756
rect 174872 79704 174878 79756
rect 174998 79704 175004 79756
rect 175056 79716 175090 79756
rect 175154 79756 175182 79908
rect 175154 79716 175188 79756
rect 175056 79704 175062 79716
rect 175182 79704 175188 79716
rect 175240 79704 175246 79756
rect 175274 79608 175280 79620
rect 174740 79580 175280 79608
rect 174596 79568 174602 79580
rect 175274 79568 175280 79580
rect 175332 79568 175338 79620
rect 173952 79512 174492 79540
rect 173952 79500 173958 79512
rect 175430 79484 175458 79908
rect 175522 79552 175550 79908
rect 175780 79840 175786 79892
rect 175838 79840 175844 79892
rect 175798 79608 175826 79840
rect 175982 79676 176010 79908
rect 176240 79840 176246 79892
rect 176298 79840 176304 79892
rect 176332 79840 176338 79892
rect 176390 79840 176396 79892
rect 176516 79840 176522 79892
rect 176574 79840 176580 79892
rect 176258 79688 176286 79840
rect 176350 79744 176378 79840
rect 176350 79716 176424 79744
rect 176396 79688 176424 79716
rect 176534 79688 176562 79840
rect 176102 79676 176108 79688
rect 175982 79648 176108 79676
rect 176102 79636 176108 79648
rect 176160 79636 176166 79688
rect 176194 79636 176200 79688
rect 176252 79648 176286 79688
rect 176252 79636 176258 79648
rect 176378 79636 176384 79688
rect 176436 79636 176442 79688
rect 176534 79648 176568 79688
rect 176562 79636 176568 79648
rect 176620 79636 176626 79688
rect 176838 79636 176844 79688
rect 176896 79676 176902 79688
rect 176994 79676 177022 79908
rect 177068 79840 177074 79892
rect 177126 79880 177132 79892
rect 177758 79880 177764 79892
rect 177126 79852 177764 79880
rect 177126 79840 177132 79852
rect 177758 79840 177764 79852
rect 177816 79840 177822 79892
rect 176896 79648 177022 79676
rect 176896 79636 176902 79648
rect 175798 79580 176148 79608
rect 175522 79512 175556 79552
rect 175550 79500 175556 79512
rect 175608 79500 175614 79552
rect 173986 79472 173992 79484
rect 173820 79444 173992 79472
rect 172664 79432 172670 79444
rect 173986 79432 173992 79444
rect 174044 79432 174050 79484
rect 175430 79444 175464 79484
rect 175458 79432 175464 79444
rect 175516 79432 175522 79484
rect 175918 79432 175924 79484
rect 175976 79472 175982 79484
rect 176120 79472 176148 79580
rect 178126 79568 178132 79620
rect 178184 79608 178190 79620
rect 191190 79608 191196 79620
rect 178184 79580 191196 79608
rect 178184 79568 178190 79580
rect 191190 79568 191196 79580
rect 191248 79568 191254 79620
rect 178310 79500 178316 79552
rect 178368 79540 178374 79552
rect 192570 79540 192576 79552
rect 178368 79512 192576 79540
rect 178368 79500 178374 79512
rect 192570 79500 192576 79512
rect 192628 79500 192634 79552
rect 217134 79500 217140 79552
rect 217192 79540 217198 79552
rect 217410 79540 217416 79552
rect 217192 79512 217416 79540
rect 217192 79500 217198 79512
rect 217410 79500 217416 79512
rect 217468 79500 217474 79552
rect 175976 79444 176148 79472
rect 175976 79432 175982 79444
rect 178954 79432 178960 79484
rect 179012 79472 179018 79484
rect 187142 79472 187148 79484
rect 179012 79444 187148 79472
rect 179012 79432 179018 79444
rect 187142 79432 187148 79444
rect 187200 79432 187206 79484
rect 194502 79432 194508 79484
rect 194560 79472 194566 79484
rect 340874 79472 340880 79484
rect 194560 79444 340880 79472
rect 194560 79432 194566 79444
rect 340874 79432 340880 79444
rect 340932 79432 340938 79484
rect 162118 79404 162124 79416
rect 148652 79376 148916 79404
rect 148980 79376 162124 79404
rect 148652 79364 148658 79376
rect 120534 79296 120540 79348
rect 120592 79336 120598 79348
rect 147766 79336 147772 79348
rect 120592 79308 147772 79336
rect 120592 79296 120598 79308
rect 147766 79296 147772 79308
rect 147824 79296 147830 79348
rect 119154 79228 119160 79280
rect 119212 79268 119218 79280
rect 146294 79268 146300 79280
rect 119212 79240 146300 79268
rect 119212 79228 119218 79240
rect 146294 79228 146300 79240
rect 146352 79228 146358 79280
rect 146386 79228 146392 79280
rect 146444 79268 146450 79280
rect 148980 79268 149008 79376
rect 162118 79364 162124 79376
rect 162176 79364 162182 79416
rect 174354 79404 174360 79416
rect 164896 79376 174360 79404
rect 149238 79296 149244 79348
rect 149296 79336 149302 79348
rect 149296 79308 157334 79336
rect 149296 79296 149302 79308
rect 146444 79240 149008 79268
rect 146444 79228 146450 79240
rect 153930 79228 153936 79280
rect 153988 79268 153994 79280
rect 154114 79268 154120 79280
rect 153988 79240 154120 79268
rect 153988 79228 153994 79240
rect 154114 79228 154120 79240
rect 154172 79228 154178 79280
rect 116302 79160 116308 79212
rect 116360 79200 116366 79212
rect 146404 79200 146432 79228
rect 116360 79172 146432 79200
rect 116360 79160 116366 79172
rect 152090 79160 152096 79212
rect 152148 79200 152154 79212
rect 157306 79200 157334 79308
rect 158346 79296 158352 79348
rect 158404 79336 158410 79348
rect 162854 79336 162860 79348
rect 158404 79308 162860 79336
rect 158404 79296 158410 79308
rect 162854 79296 162860 79308
rect 162912 79296 162918 79348
rect 164896 79200 164924 79376
rect 174354 79364 174360 79376
rect 174412 79364 174418 79416
rect 179138 79364 179144 79416
rect 179196 79404 179202 79416
rect 207750 79404 207756 79416
rect 179196 79376 207756 79404
rect 179196 79364 179202 79376
rect 207750 79364 207756 79376
rect 207808 79364 207814 79416
rect 376754 79404 376760 79416
rect 211448 79376 376760 79404
rect 211448 79348 211476 79376
rect 376754 79364 376760 79376
rect 376812 79364 376818 79416
rect 165246 79296 165252 79348
rect 165304 79336 165310 79348
rect 211430 79336 211436 79348
rect 165304 79308 211436 79336
rect 165304 79296 165310 79308
rect 211430 79296 211436 79308
rect 211488 79296 211494 79348
rect 214374 79296 214380 79348
rect 214432 79336 214438 79348
rect 448514 79336 448520 79348
rect 214432 79308 448520 79336
rect 214432 79296 214438 79308
rect 448514 79296 448520 79308
rect 448572 79296 448578 79348
rect 170858 79228 170864 79280
rect 170916 79268 170922 79280
rect 193122 79268 193128 79280
rect 170916 79240 193128 79268
rect 170916 79228 170922 79240
rect 193122 79228 193128 79240
rect 193180 79228 193186 79280
rect 152148 79172 154574 79200
rect 157306 79172 164924 79200
rect 152148 79160 152154 79172
rect 115566 79092 115572 79144
rect 115624 79132 115630 79144
rect 142246 79132 142252 79144
rect 115624 79104 142252 79132
rect 115624 79092 115630 79104
rect 142246 79092 142252 79104
rect 142304 79092 142310 79144
rect 142798 79092 142804 79144
rect 142856 79132 142862 79144
rect 143534 79132 143540 79144
rect 142856 79104 143540 79132
rect 142856 79092 142862 79104
rect 143534 79092 143540 79104
rect 143592 79092 143598 79144
rect 144914 79092 144920 79144
rect 144972 79132 144978 79144
rect 146018 79132 146024 79144
rect 144972 79104 146024 79132
rect 144972 79092 144978 79104
rect 146018 79092 146024 79104
rect 146076 79092 146082 79144
rect 118050 79024 118056 79076
rect 118108 79064 118114 79076
rect 148686 79064 148692 79076
rect 118108 79036 148692 79064
rect 118108 79024 118114 79036
rect 148686 79024 148692 79036
rect 148744 79024 148750 79076
rect 112714 78956 112720 79008
rect 112772 78996 112778 79008
rect 144730 78996 144736 79008
rect 112772 78968 144736 78996
rect 112772 78956 112778 78968
rect 144730 78956 144736 78968
rect 144788 78956 144794 79008
rect 154546 78996 154574 79172
rect 171226 79160 171232 79212
rect 171284 79200 171290 79212
rect 171284 79172 180932 79200
rect 171284 79160 171290 79172
rect 157794 79092 157800 79144
rect 157852 79132 157858 79144
rect 158070 79132 158076 79144
rect 157852 79104 158076 79132
rect 157852 79092 157858 79104
rect 158070 79092 158076 79104
rect 158128 79132 158134 79144
rect 162118 79132 162124 79144
rect 158128 79104 162124 79132
rect 158128 79092 158134 79104
rect 162118 79092 162124 79104
rect 162176 79092 162182 79144
rect 166166 79092 166172 79144
rect 166224 79132 166230 79144
rect 179046 79132 179052 79144
rect 166224 79104 179052 79132
rect 166224 79092 166230 79104
rect 179046 79092 179052 79104
rect 179104 79092 179110 79144
rect 180904 79132 180932 79172
rect 180978 79160 180984 79212
rect 181036 79200 181042 79212
rect 198182 79200 198188 79212
rect 181036 79172 198188 79200
rect 181036 79160 181042 79172
rect 198182 79160 198188 79172
rect 198240 79160 198246 79212
rect 206186 79160 206192 79212
rect 206244 79200 206250 79212
rect 206554 79200 206560 79212
rect 206244 79172 206560 79200
rect 206244 79160 206250 79172
rect 206554 79160 206560 79172
rect 206612 79160 206618 79212
rect 204622 79132 204628 79144
rect 180904 79104 204628 79132
rect 204622 79092 204628 79104
rect 204680 79092 204686 79144
rect 156046 79024 156052 79076
rect 156104 79064 156110 79076
rect 156690 79064 156696 79076
rect 156104 79036 156696 79064
rect 156104 79024 156110 79036
rect 156690 79024 156696 79036
rect 156748 79024 156754 79076
rect 158990 79024 158996 79076
rect 159048 79064 159054 79076
rect 193858 79064 193864 79076
rect 159048 79036 193864 79064
rect 159048 79024 159054 79036
rect 193858 79024 193864 79036
rect 193916 79064 193922 79076
rect 194502 79064 194508 79076
rect 193916 79036 194508 79064
rect 193916 79024 193922 79036
rect 194502 79024 194508 79036
rect 194560 79024 194566 79076
rect 162670 78996 162676 79008
rect 154546 78968 162676 78996
rect 162670 78956 162676 78968
rect 162728 78956 162734 79008
rect 167730 78956 167736 79008
rect 167788 78996 167794 79008
rect 201678 78996 201684 79008
rect 167788 78968 201684 78996
rect 167788 78956 167794 78968
rect 201678 78956 201684 78968
rect 201736 78956 201742 79008
rect 115198 78888 115204 78940
rect 115256 78928 115262 78940
rect 147674 78928 147680 78940
rect 115256 78900 147680 78928
rect 115256 78888 115262 78900
rect 147674 78888 147680 78900
rect 147732 78888 147738 78940
rect 169754 78888 169760 78940
rect 169812 78928 169818 78940
rect 204898 78928 204904 78940
rect 169812 78900 204904 78928
rect 169812 78888 169818 78900
rect 204898 78888 204904 78900
rect 204956 78888 204962 78940
rect 112438 78820 112444 78872
rect 112496 78860 112502 78872
rect 146110 78860 146116 78872
rect 112496 78832 146116 78860
rect 112496 78820 112502 78832
rect 146110 78820 146116 78832
rect 146168 78820 146174 78872
rect 167270 78820 167276 78872
rect 167328 78860 167334 78872
rect 214374 78860 214380 78872
rect 167328 78832 214380 78860
rect 167328 78820 167334 78832
rect 214374 78820 214380 78832
rect 214432 78820 214438 78872
rect 130286 78752 130292 78804
rect 130344 78792 130350 78804
rect 185578 78792 185584 78804
rect 130344 78764 141096 78792
rect 130344 78752 130350 78764
rect 113910 78724 113916 78736
rect 106246 78696 113916 78724
rect 100294 78548 100300 78600
rect 100352 78588 100358 78600
rect 106246 78588 106274 78696
rect 113910 78684 113916 78696
rect 113968 78684 113974 78736
rect 138198 78684 138204 78736
rect 138256 78724 138262 78736
rect 138566 78724 138572 78736
rect 138256 78696 138572 78724
rect 138256 78684 138262 78696
rect 138566 78684 138572 78696
rect 138624 78684 138630 78736
rect 141068 78724 141096 78764
rect 169864 78764 185584 78792
rect 143626 78724 143632 78736
rect 141068 78696 143632 78724
rect 143626 78684 143632 78696
rect 143684 78724 143690 78736
rect 144270 78724 144276 78736
rect 143684 78696 144276 78724
rect 143684 78684 143690 78696
rect 144270 78684 144276 78696
rect 144328 78684 144334 78736
rect 144546 78684 144552 78736
rect 144604 78724 144610 78736
rect 144914 78724 144920 78736
rect 144604 78696 144920 78724
rect 144604 78684 144610 78696
rect 144914 78684 144920 78696
rect 144972 78684 144978 78736
rect 157150 78684 157156 78736
rect 157208 78724 157214 78736
rect 160738 78724 160744 78736
rect 157208 78696 160744 78724
rect 157208 78684 157214 78696
rect 160738 78684 160744 78696
rect 160796 78684 160802 78736
rect 138658 78656 138664 78668
rect 100352 78560 106274 78588
rect 111076 78628 138664 78656
rect 100352 78548 100358 78560
rect 105262 78480 105268 78532
rect 105320 78520 105326 78532
rect 111076 78520 111104 78628
rect 138658 78616 138664 78628
rect 138716 78616 138722 78668
rect 139946 78616 139952 78668
rect 140004 78656 140010 78668
rect 140130 78656 140136 78668
rect 140004 78628 140136 78656
rect 140004 78616 140010 78628
rect 140130 78616 140136 78628
rect 140188 78616 140194 78668
rect 140498 78616 140504 78668
rect 140556 78656 140562 78668
rect 145006 78656 145012 78668
rect 140556 78628 145012 78656
rect 140556 78616 140562 78628
rect 145006 78616 145012 78628
rect 145064 78616 145070 78668
rect 147950 78616 147956 78668
rect 148008 78656 148014 78668
rect 148318 78656 148324 78668
rect 148008 78628 148324 78656
rect 148008 78616 148014 78628
rect 148318 78616 148324 78628
rect 148376 78616 148382 78668
rect 157426 78616 157432 78668
rect 157484 78656 157490 78668
rect 157886 78656 157892 78668
rect 157484 78628 157892 78656
rect 157484 78616 157490 78628
rect 157886 78616 157892 78628
rect 157944 78616 157950 78668
rect 158162 78616 158168 78668
rect 158220 78656 158226 78668
rect 158346 78656 158352 78668
rect 158220 78628 158352 78656
rect 158220 78616 158226 78628
rect 158346 78616 158352 78628
rect 158404 78616 158410 78668
rect 159266 78616 159272 78668
rect 159324 78656 159330 78668
rect 159450 78656 159456 78668
rect 159324 78628 159456 78656
rect 159324 78616 159330 78628
rect 159450 78616 159456 78628
rect 159508 78616 159514 78668
rect 113910 78548 113916 78600
rect 113968 78588 113974 78600
rect 113968 78560 139532 78588
rect 113968 78548 113974 78560
rect 105320 78492 111104 78520
rect 105320 78480 105326 78492
rect 122190 78480 122196 78532
rect 122248 78520 122254 78532
rect 122248 78492 139440 78520
rect 122248 78480 122254 78492
rect 105538 78412 105544 78464
rect 105596 78452 105602 78464
rect 105722 78452 105728 78464
rect 105596 78424 105728 78452
rect 105596 78412 105602 78424
rect 105722 78412 105728 78424
rect 105780 78452 105786 78464
rect 136910 78452 136916 78464
rect 105780 78424 136916 78452
rect 105780 78412 105786 78424
rect 136910 78412 136916 78424
rect 136968 78412 136974 78464
rect 107194 78384 107200 78396
rect 103486 78356 107200 78384
rect 60734 78276 60740 78328
rect 60792 78316 60798 78328
rect 103486 78316 103514 78356
rect 107194 78344 107200 78356
rect 107252 78384 107258 78396
rect 137186 78384 137192 78396
rect 107252 78356 137192 78384
rect 107252 78344 107258 78356
rect 137186 78344 137192 78356
rect 137244 78344 137250 78396
rect 136266 78316 136272 78328
rect 60792 78288 103514 78316
rect 107948 78288 136272 78316
rect 60792 78276 60798 78288
rect 75914 78208 75920 78260
rect 75972 78248 75978 78260
rect 105722 78248 105728 78260
rect 75972 78220 105728 78248
rect 75972 78208 75978 78220
rect 105722 78208 105728 78220
rect 105780 78208 105786 78260
rect 57974 78072 57980 78124
rect 58032 78112 58038 78124
rect 107286 78112 107292 78124
rect 58032 78084 107292 78112
rect 58032 78072 58038 78084
rect 107286 78072 107292 78084
rect 107344 78112 107350 78124
rect 107948 78112 107976 78288
rect 136266 78276 136272 78288
rect 136324 78276 136330 78328
rect 139412 78316 139440 78492
rect 139504 78452 139532 78560
rect 161474 78548 161480 78600
rect 161532 78588 161538 78600
rect 161658 78588 161664 78600
rect 161532 78560 161664 78588
rect 161532 78548 161538 78560
rect 161658 78548 161664 78560
rect 161716 78548 161722 78600
rect 169864 78588 169892 78764
rect 185578 78752 185584 78764
rect 185636 78752 185642 78804
rect 209222 78752 209228 78804
rect 209280 78792 209286 78804
rect 480254 78792 480260 78804
rect 209280 78764 480260 78792
rect 209280 78752 209286 78764
rect 480254 78752 480260 78764
rect 480312 78752 480318 78804
rect 171042 78684 171048 78736
rect 171100 78724 171106 78736
rect 174722 78724 174728 78736
rect 171100 78696 174728 78724
rect 171100 78684 171106 78696
rect 174722 78684 174728 78696
rect 174780 78684 174786 78736
rect 211798 78684 211804 78736
rect 211856 78724 211862 78736
rect 483014 78724 483020 78736
rect 211856 78696 483020 78724
rect 211856 78684 211862 78696
rect 483014 78684 483020 78696
rect 483072 78684 483078 78736
rect 169938 78616 169944 78668
rect 169996 78656 170002 78668
rect 169996 78628 178034 78656
rect 169996 78616 170002 78628
rect 169864 78560 169984 78588
rect 169956 78532 169984 78560
rect 171502 78548 171508 78600
rect 171560 78588 171566 78600
rect 172238 78588 172244 78600
rect 171560 78560 172244 78588
rect 171560 78548 171566 78560
rect 172238 78548 172244 78560
rect 172296 78548 172302 78600
rect 178006 78588 178034 78628
rect 179046 78616 179052 78668
rect 179104 78656 179110 78668
rect 179230 78656 179236 78668
rect 179104 78628 179236 78656
rect 179104 78616 179110 78628
rect 179230 78616 179236 78628
rect 179288 78656 179294 78668
rect 200942 78656 200948 78668
rect 179288 78628 200948 78656
rect 179288 78616 179294 78628
rect 200942 78616 200948 78628
rect 201000 78616 201006 78668
rect 211798 78588 211804 78600
rect 178006 78560 211804 78588
rect 211798 78548 211804 78560
rect 211856 78548 211862 78600
rect 169938 78480 169944 78532
rect 169996 78480 170002 78532
rect 199102 78520 199108 78532
rect 170048 78492 199108 78520
rect 153930 78452 153936 78464
rect 139504 78424 153936 78452
rect 153930 78412 153936 78424
rect 153988 78412 153994 78464
rect 161658 78412 161664 78464
rect 161716 78452 161722 78464
rect 162486 78452 162492 78464
rect 161716 78424 162492 78452
rect 161716 78412 161722 78424
rect 162486 78412 162492 78424
rect 162544 78412 162550 78464
rect 165154 78412 165160 78464
rect 165212 78452 165218 78464
rect 170048 78452 170076 78492
rect 199102 78480 199108 78492
rect 199160 78520 199166 78532
rect 199562 78520 199568 78532
rect 199160 78492 199568 78520
rect 199160 78480 199166 78492
rect 199562 78480 199568 78492
rect 199620 78480 199626 78532
rect 197630 78452 197636 78464
rect 165212 78424 170076 78452
rect 170140 78424 197636 78452
rect 165212 78412 165218 78424
rect 139578 78344 139584 78396
rect 139636 78384 139642 78396
rect 140406 78384 140412 78396
rect 139636 78356 140412 78384
rect 139636 78344 139642 78356
rect 140406 78344 140412 78356
rect 140464 78344 140470 78396
rect 147950 78344 147956 78396
rect 148008 78384 148014 78396
rect 149146 78384 149152 78396
rect 148008 78356 149152 78384
rect 148008 78344 148014 78356
rect 149146 78344 149152 78356
rect 149204 78344 149210 78396
rect 163130 78344 163136 78396
rect 163188 78384 163194 78396
rect 170140 78384 170168 78424
rect 197630 78412 197636 78424
rect 197688 78412 197694 78464
rect 198734 78384 198740 78396
rect 163188 78356 170168 78384
rect 170232 78356 198740 78384
rect 163188 78344 163194 78356
rect 143534 78316 143540 78328
rect 139412 78288 143540 78316
rect 143534 78276 143540 78288
rect 143592 78276 143598 78328
rect 136542 78248 136548 78260
rect 107344 78084 107976 78112
rect 108040 78220 136548 78248
rect 107344 78072 107350 78084
rect 53834 78004 53840 78056
rect 53892 78044 53898 78056
rect 106918 78044 106924 78056
rect 53892 78016 106924 78044
rect 53892 78004 53898 78016
rect 106918 78004 106924 78016
rect 106976 78044 106982 78056
rect 108040 78044 108068 78220
rect 136542 78208 136548 78220
rect 136600 78208 136606 78260
rect 145834 78208 145840 78260
rect 145892 78208 145898 78260
rect 160738 78208 160744 78260
rect 160796 78248 160802 78260
rect 162486 78248 162492 78260
rect 160796 78220 162492 78248
rect 160796 78208 160802 78220
rect 162486 78208 162492 78220
rect 162544 78208 162550 78260
rect 164234 78208 164240 78260
rect 164292 78248 164298 78260
rect 170232 78248 170260 78356
rect 198734 78344 198740 78356
rect 198792 78344 198798 78396
rect 171134 78276 171140 78328
rect 171192 78316 171198 78328
rect 203518 78316 203524 78328
rect 171192 78288 203524 78316
rect 171192 78276 171198 78288
rect 203518 78276 203524 78288
rect 203576 78276 203582 78328
rect 164292 78220 170260 78248
rect 164292 78208 164298 78220
rect 172422 78208 172428 78260
rect 172480 78248 172486 78260
rect 180058 78248 180064 78260
rect 172480 78220 180064 78248
rect 172480 78208 172486 78220
rect 180058 78208 180064 78220
rect 180116 78208 180122 78260
rect 135254 78180 135260 78192
rect 106976 78016 108068 78044
rect 108132 78152 135260 78180
rect 106976 78004 106982 78016
rect 46934 77936 46940 77988
rect 46992 77976 46998 77988
rect 107010 77976 107016 77988
rect 46992 77948 107016 77976
rect 46992 77936 46998 77948
rect 107010 77936 107016 77948
rect 107068 77976 107074 77988
rect 108132 77976 108160 78152
rect 135254 78140 135260 78152
rect 135312 78140 135318 78192
rect 136726 78140 136732 78192
rect 136784 78180 136790 78192
rect 137278 78180 137284 78192
rect 136784 78152 137284 78180
rect 136784 78140 136790 78152
rect 137278 78140 137284 78152
rect 137336 78140 137342 78192
rect 140130 78140 140136 78192
rect 140188 78180 140194 78192
rect 140774 78180 140780 78192
rect 140188 78152 140780 78180
rect 140188 78140 140194 78152
rect 140774 78140 140780 78152
rect 140832 78140 140838 78192
rect 142246 78140 142252 78192
rect 142304 78180 142310 78192
rect 145282 78180 145288 78192
rect 142304 78152 145288 78180
rect 142304 78140 142310 78152
rect 145282 78140 145288 78152
rect 145340 78180 145346 78192
rect 145852 78180 145880 78208
rect 145340 78152 145880 78180
rect 145340 78140 145346 78152
rect 152918 78140 152924 78192
rect 152976 78180 152982 78192
rect 156230 78180 156236 78192
rect 152976 78152 156236 78180
rect 152976 78140 152982 78152
rect 156230 78140 156236 78152
rect 156288 78140 156294 78192
rect 164142 78140 164148 78192
rect 164200 78180 164206 78192
rect 178770 78180 178776 78192
rect 164200 78152 178776 78180
rect 164200 78140 164206 78152
rect 178770 78140 178776 78152
rect 178828 78180 178834 78192
rect 179138 78180 179144 78192
rect 178828 78152 179144 78180
rect 178828 78140 178834 78152
rect 179138 78140 179144 78152
rect 179196 78140 179202 78192
rect 179322 78140 179328 78192
rect 179380 78180 179386 78192
rect 213086 78180 213092 78192
rect 179380 78152 213092 78180
rect 179380 78140 179386 78152
rect 213086 78140 213092 78152
rect 213144 78140 213150 78192
rect 120718 78072 120724 78124
rect 120776 78112 120782 78124
rect 145650 78112 145656 78124
rect 120776 78084 145656 78112
rect 120776 78072 120782 78084
rect 145650 78072 145656 78084
rect 145708 78072 145714 78124
rect 164234 78072 164240 78124
rect 164292 78112 164298 78124
rect 164786 78112 164792 78124
rect 164292 78084 164792 78112
rect 164292 78072 164298 78084
rect 164786 78072 164792 78084
rect 164844 78072 164850 78124
rect 169386 78072 169392 78124
rect 169444 78112 169450 78124
rect 169570 78112 169576 78124
rect 169444 78084 169576 78112
rect 169444 78072 169450 78084
rect 169570 78072 169576 78084
rect 169628 78112 169634 78124
rect 171134 78112 171140 78124
rect 169628 78084 171140 78112
rect 169628 78072 169634 78084
rect 171134 78072 171140 78084
rect 171192 78072 171198 78124
rect 171318 78072 171324 78124
rect 171376 78112 171382 78124
rect 187694 78112 187700 78124
rect 171376 78084 187700 78112
rect 171376 78072 171382 78084
rect 187694 78072 187700 78084
rect 187752 78072 187758 78124
rect 197630 78072 197636 78124
rect 197688 78112 197694 78124
rect 198458 78112 198464 78124
rect 197688 78084 198464 78112
rect 197688 78072 197694 78084
rect 198458 78072 198464 78084
rect 198516 78112 198522 78124
rect 393314 78112 393320 78124
rect 198516 78084 393320 78112
rect 198516 78072 198522 78084
rect 393314 78072 393320 78084
rect 393372 78072 393378 78124
rect 108298 78004 108304 78056
rect 108356 78044 108362 78056
rect 129826 78044 129832 78056
rect 108356 78016 129832 78044
rect 108356 78004 108362 78016
rect 129826 78004 129832 78016
rect 129884 78044 129890 78056
rect 130654 78044 130660 78056
rect 129884 78016 130660 78044
rect 129884 78004 129890 78016
rect 130654 78004 130660 78016
rect 130712 78004 130718 78056
rect 130746 78004 130752 78056
rect 130804 78044 130810 78056
rect 142062 78044 142068 78056
rect 130804 78016 142068 78044
rect 130804 78004 130810 78016
rect 142062 78004 142068 78016
rect 142120 78004 142126 78056
rect 152918 78004 152924 78056
rect 152976 78044 152982 78056
rect 153194 78044 153200 78056
rect 152976 78016 153200 78044
rect 152976 78004 152982 78016
rect 153194 78004 153200 78016
rect 153252 78004 153258 78056
rect 158438 78004 158444 78056
rect 158496 78044 158502 78056
rect 162210 78044 162216 78056
rect 158496 78016 162216 78044
rect 158496 78004 158502 78016
rect 162210 78004 162216 78016
rect 162268 78004 162274 78056
rect 164050 78004 164056 78056
rect 164108 78044 164114 78056
rect 178678 78044 178684 78056
rect 164108 78016 178684 78044
rect 164108 78004 164114 78016
rect 178678 78004 178684 78016
rect 178736 78044 178742 78056
rect 178954 78044 178960 78056
rect 178736 78016 178960 78044
rect 178736 78004 178742 78016
rect 178954 78004 178960 78016
rect 179012 78004 179018 78056
rect 198734 78004 198740 78056
rect 198792 78044 198798 78056
rect 199470 78044 199476 78056
rect 198792 78016 199476 78044
rect 198792 78004 198798 78016
rect 199470 78004 199476 78016
rect 199528 78044 199534 78056
rect 415486 78044 415492 78056
rect 199528 78016 415492 78044
rect 199528 78004 199534 78016
rect 415486 78004 415492 78016
rect 415544 78004 415550 78056
rect 107068 77948 108160 77976
rect 107068 77936 107074 77948
rect 108390 77936 108396 77988
rect 108448 77976 108454 77988
rect 131206 77976 131212 77988
rect 108448 77948 131212 77976
rect 108448 77936 108454 77948
rect 131206 77936 131212 77948
rect 131264 77976 131270 77988
rect 142522 77976 142528 77988
rect 131264 77948 142528 77976
rect 131264 77936 131270 77948
rect 142522 77936 142528 77948
rect 142580 77936 142586 77988
rect 156506 77936 156512 77988
rect 156564 77976 156570 77988
rect 156874 77976 156880 77988
rect 156564 77948 156880 77976
rect 156564 77936 156570 77948
rect 156874 77936 156880 77948
rect 156932 77936 156938 77988
rect 166902 77936 166908 77988
rect 166960 77976 166966 77988
rect 170490 77976 170496 77988
rect 166960 77948 170496 77976
rect 166960 77936 166966 77948
rect 170490 77936 170496 77948
rect 170548 77936 170554 77988
rect 175550 77936 175556 77988
rect 175608 77976 175614 77988
rect 176102 77976 176108 77988
rect 175608 77948 176108 77976
rect 175608 77936 175614 77948
rect 176102 77936 176108 77948
rect 176160 77936 176166 77988
rect 177942 77936 177948 77988
rect 178000 77976 178006 77988
rect 181990 77976 181996 77988
rect 178000 77948 181996 77976
rect 178000 77936 178006 77948
rect 181990 77936 181996 77948
rect 182048 77936 182054 77988
rect 199102 77936 199108 77988
rect 199160 77976 199166 77988
rect 422294 77976 422300 77988
rect 199160 77948 422300 77976
rect 199160 77936 199166 77948
rect 422294 77936 422300 77948
rect 422352 77936 422358 77988
rect 109494 77868 109500 77920
rect 109552 77908 109558 77920
rect 129734 77908 129740 77920
rect 109552 77880 129740 77908
rect 109552 77868 109558 77880
rect 129734 77868 129740 77880
rect 129792 77868 129798 77920
rect 130654 77868 130660 77920
rect 130712 77908 130718 77920
rect 137370 77908 137376 77920
rect 130712 77880 137376 77908
rect 130712 77868 130718 77880
rect 137370 77868 137376 77880
rect 137428 77868 137434 77920
rect 138750 77868 138756 77920
rect 138808 77908 138814 77920
rect 139302 77908 139308 77920
rect 138808 77880 139308 77908
rect 138808 77868 138814 77880
rect 139302 77868 139308 77880
rect 139360 77868 139366 77920
rect 143810 77868 143816 77920
rect 143868 77908 143874 77920
rect 144454 77908 144460 77920
rect 143868 77880 144460 77908
rect 143868 77868 143874 77880
rect 144454 77868 144460 77880
rect 144512 77868 144518 77920
rect 168282 77868 168288 77920
rect 168340 77908 168346 77920
rect 180610 77908 180616 77920
rect 168340 77880 180616 77908
rect 168340 77868 168346 77880
rect 180610 77868 180616 77880
rect 180668 77908 180674 77920
rect 201770 77908 201776 77920
rect 180668 77880 201776 77908
rect 180668 77868 180674 77880
rect 201770 77868 201776 77880
rect 201828 77868 201834 77920
rect 108114 77800 108120 77852
rect 108172 77840 108178 77852
rect 128538 77840 128544 77852
rect 108172 77812 128544 77840
rect 108172 77800 108178 77812
rect 128538 77800 128544 77812
rect 128596 77800 128602 77852
rect 129918 77800 129924 77852
rect 129976 77840 129982 77852
rect 133874 77840 133880 77852
rect 129976 77812 133880 77840
rect 129976 77800 129982 77812
rect 133874 77800 133880 77812
rect 133932 77800 133938 77852
rect 134518 77800 134524 77852
rect 134576 77840 134582 77852
rect 142246 77840 142252 77852
rect 134576 77812 142252 77840
rect 134576 77800 134582 77812
rect 142246 77800 142252 77812
rect 142304 77800 142310 77852
rect 170490 77800 170496 77852
rect 170548 77840 170554 77852
rect 179138 77840 179144 77852
rect 170548 77812 179144 77840
rect 170548 77800 170554 77812
rect 179138 77800 179144 77812
rect 179196 77840 179202 77852
rect 179322 77840 179328 77852
rect 179196 77812 179328 77840
rect 179196 77800 179202 77812
rect 179322 77800 179328 77812
rect 179380 77800 179386 77852
rect 179966 77800 179972 77852
rect 180024 77840 180030 77852
rect 191282 77840 191288 77852
rect 180024 77812 191288 77840
rect 180024 77800 180030 77812
rect 191282 77800 191288 77812
rect 191340 77800 191346 77852
rect 99834 77732 99840 77784
rect 99892 77772 99898 77784
rect 99892 77744 122834 77772
rect 99892 77732 99898 77744
rect 122806 77636 122834 77744
rect 130930 77732 130936 77784
rect 130988 77772 130994 77784
rect 139486 77772 139492 77784
rect 130988 77744 139492 77772
rect 130988 77732 130994 77744
rect 139486 77732 139492 77744
rect 139544 77732 139550 77784
rect 162394 77732 162400 77784
rect 162452 77772 162458 77784
rect 162762 77772 162768 77784
rect 162452 77744 162768 77772
rect 162452 77732 162458 77744
rect 162762 77732 162768 77744
rect 162820 77732 162826 77784
rect 167178 77732 167184 77784
rect 167236 77772 167242 77784
rect 179046 77772 179052 77784
rect 167236 77744 179052 77772
rect 167236 77732 167242 77744
rect 179046 77732 179052 77744
rect 179104 77732 179110 77784
rect 130654 77664 130660 77716
rect 130712 77704 130718 77716
rect 131022 77704 131028 77716
rect 130712 77676 131028 77704
rect 130712 77664 130718 77676
rect 131022 77664 131028 77676
rect 131080 77704 131086 77716
rect 144086 77704 144092 77716
rect 131080 77676 144092 77704
rect 131080 77664 131086 77676
rect 144086 77664 144092 77676
rect 144144 77664 144150 77716
rect 148410 77664 148416 77716
rect 148468 77704 148474 77716
rect 207842 77704 207848 77716
rect 148468 77676 207848 77704
rect 148468 77664 148474 77676
rect 207842 77664 207848 77676
rect 207900 77664 207906 77716
rect 132862 77636 132868 77648
rect 122806 77608 132868 77636
rect 132862 77596 132868 77608
rect 132920 77596 132926 77648
rect 133874 77596 133880 77648
rect 133932 77636 133938 77648
rect 134334 77636 134340 77648
rect 133932 77608 134340 77636
rect 133932 77596 133938 77608
rect 134334 77596 134340 77608
rect 134392 77596 134398 77648
rect 140406 77596 140412 77648
rect 140464 77636 140470 77648
rect 140682 77636 140688 77648
rect 140464 77608 140688 77636
rect 140464 77596 140470 77608
rect 140682 77596 140688 77608
rect 140740 77596 140746 77648
rect 150894 77596 150900 77648
rect 150952 77636 150958 77648
rect 169938 77636 169944 77648
rect 150952 77608 169944 77636
rect 150952 77596 150958 77608
rect 169938 77596 169944 77608
rect 169996 77596 170002 77648
rect 175734 77596 175740 77648
rect 175792 77636 175798 77648
rect 176194 77636 176200 77648
rect 175792 77608 176200 77636
rect 175792 77596 175798 77608
rect 176194 77596 176200 77608
rect 176252 77596 176258 77648
rect 176654 77596 176660 77648
rect 176712 77636 176718 77648
rect 176838 77636 176844 77648
rect 176712 77608 176844 77636
rect 176712 77596 176718 77608
rect 176838 77596 176844 77608
rect 176896 77596 176902 77648
rect 177758 77596 177764 77648
rect 177816 77636 177822 77648
rect 211706 77636 211712 77648
rect 177816 77608 211712 77636
rect 177816 77596 177822 77608
rect 211706 77596 211712 77608
rect 211764 77596 211770 77648
rect 145006 77528 145012 77580
rect 145064 77568 145070 77580
rect 145558 77568 145564 77580
rect 145064 77540 145564 77568
rect 145064 77528 145070 77540
rect 145558 77528 145564 77540
rect 145616 77528 145622 77580
rect 157518 77528 157524 77580
rect 157576 77568 157582 77580
rect 170858 77568 170864 77580
rect 157576 77540 170864 77568
rect 157576 77528 157582 77540
rect 170858 77528 170864 77540
rect 170916 77528 170922 77580
rect 174354 77528 174360 77580
rect 174412 77568 174418 77580
rect 178862 77568 178868 77580
rect 174412 77540 178868 77568
rect 174412 77528 174418 77540
rect 178862 77528 178868 77540
rect 178920 77528 178926 77580
rect 146294 77460 146300 77512
rect 146352 77500 146358 77512
rect 146846 77500 146852 77512
rect 146352 77472 146852 77500
rect 146352 77460 146358 77472
rect 146846 77460 146852 77472
rect 146904 77460 146910 77512
rect 148686 77460 148692 77512
rect 148744 77500 148750 77512
rect 148962 77500 148968 77512
rect 148744 77472 148968 77500
rect 148744 77460 148750 77472
rect 148962 77460 148968 77472
rect 149020 77460 149026 77512
rect 161842 77460 161848 77512
rect 161900 77500 161906 77512
rect 162394 77500 162400 77512
rect 161900 77472 162400 77500
rect 161900 77460 161906 77472
rect 162394 77460 162400 77472
rect 162452 77460 162458 77512
rect 167362 77460 167368 77512
rect 167420 77500 167426 77512
rect 178494 77500 178500 77512
rect 167420 77472 178500 77500
rect 167420 77460 167426 77472
rect 178494 77460 178500 77472
rect 178552 77460 178558 77512
rect 133046 77432 133052 77444
rect 132604 77404 133052 77432
rect 132604 77376 132632 77404
rect 133046 77392 133052 77404
rect 133104 77392 133110 77444
rect 146018 77392 146024 77444
rect 146076 77432 146082 77444
rect 146938 77432 146944 77444
rect 146076 77404 146944 77432
rect 146076 77392 146082 77404
rect 146938 77392 146944 77404
rect 146996 77392 147002 77444
rect 169938 77392 169944 77444
rect 169996 77432 170002 77444
rect 170674 77432 170680 77444
rect 169996 77404 170680 77432
rect 169996 77392 170002 77404
rect 170674 77392 170680 77404
rect 170732 77392 170738 77444
rect 132586 77324 132592 77376
rect 132644 77324 132650 77376
rect 132770 77324 132776 77376
rect 132828 77364 132834 77376
rect 133230 77364 133236 77376
rect 132828 77336 133236 77364
rect 132828 77324 132834 77336
rect 133230 77324 133236 77336
rect 133288 77324 133294 77376
rect 135622 77324 135628 77376
rect 135680 77364 135686 77376
rect 136266 77364 136272 77376
rect 135680 77336 136272 77364
rect 135680 77324 135686 77336
rect 136266 77324 136272 77336
rect 136324 77324 136330 77376
rect 175826 77324 175832 77376
rect 175884 77364 175890 77376
rect 176562 77364 176568 77376
rect 175884 77336 176568 77364
rect 175884 77324 175890 77336
rect 176562 77324 176568 77336
rect 176620 77324 176626 77376
rect 109034 77256 109040 77308
rect 109092 77296 109098 77308
rect 109494 77296 109500 77308
rect 109092 77268 109500 77296
rect 109092 77256 109098 77268
rect 109494 77256 109500 77268
rect 109552 77256 109558 77308
rect 132494 77256 132500 77308
rect 132552 77296 132558 77308
rect 133414 77296 133420 77308
rect 132552 77268 133420 77296
rect 132552 77256 132558 77268
rect 133414 77256 133420 77268
rect 133472 77256 133478 77308
rect 135806 77256 135812 77308
rect 135864 77296 135870 77308
rect 136174 77296 136180 77308
rect 135864 77268 136180 77296
rect 135864 77256 135870 77268
rect 136174 77256 136180 77268
rect 136232 77256 136238 77308
rect 138290 77256 138296 77308
rect 138348 77296 138354 77308
rect 138474 77296 138480 77308
rect 138348 77268 138480 77296
rect 138348 77256 138354 77268
rect 138474 77256 138480 77268
rect 138532 77256 138538 77308
rect 154942 77256 154948 77308
rect 155000 77296 155006 77308
rect 164878 77296 164884 77308
rect 155000 77268 164884 77296
rect 155000 77256 155006 77268
rect 164878 77256 164884 77268
rect 164936 77256 164942 77308
rect 174170 77256 174176 77308
rect 174228 77296 174234 77308
rect 177574 77296 177580 77308
rect 174228 77268 177580 77296
rect 174228 77256 174234 77268
rect 177574 77256 177580 77268
rect 177632 77256 177638 77308
rect 187694 77256 187700 77308
rect 187752 77296 187758 77308
rect 500954 77296 500960 77308
rect 187752 77268 500960 77296
rect 187752 77256 187758 77268
rect 500954 77256 500960 77268
rect 501012 77256 501018 77308
rect 111242 77188 111248 77240
rect 111300 77228 111306 77240
rect 145098 77228 145104 77240
rect 111300 77200 145104 77228
rect 111300 77188 111306 77200
rect 145098 77188 145104 77200
rect 145156 77228 145162 77240
rect 146018 77228 146024 77240
rect 145156 77200 146024 77228
rect 145156 77188 145162 77200
rect 146018 77188 146024 77200
rect 146076 77188 146082 77240
rect 155494 77188 155500 77240
rect 155552 77228 155558 77240
rect 217134 77228 217140 77240
rect 155552 77200 217140 77228
rect 155552 77188 155558 77200
rect 217134 77188 217140 77200
rect 217192 77188 217198 77240
rect 124858 77120 124864 77172
rect 124916 77160 124922 77172
rect 125594 77160 125600 77172
rect 124916 77132 125600 77160
rect 124916 77120 124922 77132
rect 125594 77120 125600 77132
rect 125652 77160 125658 77172
rect 141878 77160 141884 77172
rect 125652 77132 141884 77160
rect 125652 77120 125658 77132
rect 141878 77120 141884 77132
rect 141936 77120 141942 77172
rect 145926 77120 145932 77172
rect 145984 77160 145990 77172
rect 148318 77160 148324 77172
rect 145984 77132 148324 77160
rect 145984 77120 145990 77132
rect 148318 77120 148324 77132
rect 148376 77120 148382 77172
rect 213178 77160 213184 77172
rect 160066 77132 213184 77160
rect 102134 77052 102140 77104
rect 102192 77092 102198 77104
rect 102870 77092 102876 77104
rect 102192 77064 102876 77092
rect 102192 77052 102198 77064
rect 102870 77052 102876 77064
rect 102928 77092 102934 77104
rect 137462 77092 137468 77104
rect 102928 77064 137468 77092
rect 102928 77052 102934 77064
rect 137462 77052 137468 77064
rect 137520 77052 137526 77104
rect 114462 76984 114468 77036
rect 114520 77024 114526 77036
rect 147122 77024 147128 77036
rect 114520 76996 147128 77024
rect 114520 76984 114526 76996
rect 147122 76984 147128 76996
rect 147180 76984 147186 77036
rect 114278 76916 114284 76968
rect 114336 76956 114342 76968
rect 146754 76956 146760 76968
rect 114336 76928 146760 76956
rect 114336 76916 114342 76928
rect 146754 76916 146760 76928
rect 146812 76916 146818 76968
rect 115290 76848 115296 76900
rect 115348 76888 115354 76900
rect 149698 76888 149704 76900
rect 115348 76860 149704 76888
rect 115348 76848 115354 76860
rect 149698 76848 149704 76860
rect 149756 76848 149762 76900
rect 152182 76848 152188 76900
rect 152240 76888 152246 76900
rect 160066 76888 160094 77132
rect 213178 77120 213184 77132
rect 213236 77160 213242 77172
rect 213236 77132 219434 77160
rect 213236 77120 213242 77132
rect 164878 77052 164884 77104
rect 164936 77092 164942 77104
rect 164936 77064 215524 77092
rect 164936 77052 164942 77064
rect 170030 76984 170036 77036
rect 170088 77024 170094 77036
rect 170766 77024 170772 77036
rect 170088 76996 170772 77024
rect 170088 76984 170094 76996
rect 170766 76984 170772 76996
rect 170824 76984 170830 77036
rect 171226 76984 171232 77036
rect 171284 77024 171290 77036
rect 171410 77024 171416 77036
rect 171284 76996 171416 77024
rect 171284 76984 171290 76996
rect 171410 76984 171416 76996
rect 171468 76984 171474 77036
rect 174170 76984 174176 77036
rect 174228 77024 174234 77036
rect 174906 77024 174912 77036
rect 174228 76996 174912 77024
rect 174228 76984 174234 76996
rect 174906 76984 174912 76996
rect 174964 76984 174970 77036
rect 175458 76984 175464 77036
rect 175516 77024 175522 77036
rect 210510 77024 210516 77036
rect 175516 76996 210516 77024
rect 175516 76984 175522 76996
rect 210510 76984 210516 76996
rect 210568 76984 210574 77036
rect 165338 76916 165344 76968
rect 165396 76956 165402 76968
rect 199378 76956 199384 76968
rect 165396 76928 199384 76956
rect 165396 76916 165402 76928
rect 199378 76916 199384 76928
rect 199436 76916 199442 76968
rect 152240 76860 160094 76888
rect 152240 76848 152246 76860
rect 160186 76848 160192 76900
rect 160244 76888 160250 76900
rect 160738 76888 160744 76900
rect 160244 76860 160744 76888
rect 160244 76848 160250 76860
rect 160738 76848 160744 76860
rect 160796 76848 160802 76900
rect 161566 76848 161572 76900
rect 161624 76888 161630 76900
rect 164142 76888 164148 76900
rect 161624 76860 164148 76888
rect 161624 76848 161630 76860
rect 164142 76848 164148 76860
rect 164200 76848 164206 76900
rect 165798 76848 165804 76900
rect 165856 76888 165862 76900
rect 166166 76888 166172 76900
rect 165856 76860 166172 76888
rect 165856 76848 165862 76860
rect 166166 76848 166172 76860
rect 166224 76848 166230 76900
rect 169846 76848 169852 76900
rect 169904 76888 169910 76900
rect 170306 76888 170312 76900
rect 169904 76860 170312 76888
rect 169904 76848 169910 76860
rect 170306 76848 170312 76860
rect 170364 76848 170370 76900
rect 172698 76848 172704 76900
rect 172756 76888 172762 76900
rect 173526 76888 173532 76900
rect 172756 76860 173532 76888
rect 172756 76848 172762 76860
rect 173526 76848 173532 76860
rect 173584 76848 173590 76900
rect 175458 76848 175464 76900
rect 175516 76888 175522 76900
rect 176378 76888 176384 76900
rect 175516 76860 176384 76888
rect 175516 76848 175522 76860
rect 176378 76848 176384 76860
rect 176436 76848 176442 76900
rect 177850 76848 177856 76900
rect 177908 76888 177914 76900
rect 210418 76888 210424 76900
rect 177908 76860 210424 76888
rect 177908 76848 177914 76860
rect 210418 76848 210424 76860
rect 210476 76848 210482 76900
rect 112990 76780 112996 76832
rect 113048 76820 113054 76832
rect 144362 76820 144368 76832
rect 113048 76792 144368 76820
rect 113048 76780 113054 76792
rect 144362 76780 144368 76792
rect 144420 76780 144426 76832
rect 153286 76780 153292 76832
rect 153344 76820 153350 76832
rect 154022 76820 154028 76832
rect 153344 76792 154028 76820
rect 153344 76780 153350 76792
rect 154022 76780 154028 76792
rect 154080 76780 154086 76832
rect 189258 76820 189264 76832
rect 160066 76792 189264 76820
rect 114370 76712 114376 76764
rect 114428 76752 114434 76764
rect 145742 76752 145748 76764
rect 114428 76724 145748 76752
rect 114428 76712 114434 76724
rect 145742 76712 145748 76724
rect 145800 76752 145806 76764
rect 152550 76752 152556 76764
rect 145800 76724 152556 76752
rect 145800 76712 145806 76724
rect 152550 76712 152556 76724
rect 152608 76712 152614 76764
rect 99374 76644 99380 76696
rect 99432 76684 99438 76696
rect 110874 76684 110880 76696
rect 99432 76656 110880 76684
rect 99432 76644 99438 76656
rect 110874 76644 110880 76656
rect 110932 76684 110938 76696
rect 140038 76684 140044 76696
rect 110932 76656 140044 76684
rect 110932 76644 110938 76656
rect 140038 76644 140044 76656
rect 140096 76644 140102 76696
rect 140958 76644 140964 76696
rect 141016 76684 141022 76696
rect 141234 76684 141240 76696
rect 141016 76656 141240 76684
rect 141016 76644 141022 76656
rect 141234 76644 141240 76656
rect 141292 76644 141298 76696
rect 150526 76644 150532 76696
rect 150584 76684 150590 76696
rect 151630 76684 151636 76696
rect 150584 76656 151636 76684
rect 150584 76644 150590 76656
rect 151630 76644 151636 76656
rect 151688 76644 151694 76696
rect 151906 76644 151912 76696
rect 151964 76684 151970 76696
rect 152458 76684 152464 76696
rect 151964 76656 152464 76684
rect 151964 76644 151970 76656
rect 152458 76644 152464 76656
rect 152516 76644 152522 76696
rect 159818 76644 159824 76696
rect 159876 76684 159882 76696
rect 160066 76684 160094 76792
rect 189258 76780 189264 76792
rect 189316 76780 189322 76832
rect 193122 76780 193128 76832
rect 193180 76820 193186 76832
rect 214558 76820 214564 76832
rect 193180 76792 214564 76820
rect 193180 76780 193186 76792
rect 214558 76780 214564 76792
rect 214616 76820 214622 76832
rect 215496 76820 215524 77064
rect 219406 76888 219434 77132
rect 247678 76888 247684 76900
rect 219406 76860 247684 76888
rect 247678 76848 247684 76860
rect 247736 76848 247742 76900
rect 217318 76820 217324 76832
rect 214616 76792 215294 76820
rect 215496 76792 217324 76820
rect 214616 76780 214622 76792
rect 162854 76712 162860 76764
rect 162912 76752 162918 76764
rect 163682 76752 163688 76764
rect 162912 76724 163688 76752
rect 162912 76712 162918 76724
rect 163682 76712 163688 76724
rect 163740 76712 163746 76764
rect 164326 76712 164332 76764
rect 164384 76752 164390 76764
rect 164786 76752 164792 76764
rect 164384 76724 164792 76752
rect 164384 76712 164390 76724
rect 164786 76712 164792 76724
rect 164844 76712 164850 76764
rect 167362 76712 167368 76764
rect 167420 76752 167426 76764
rect 167546 76752 167552 76764
rect 167420 76724 167552 76752
rect 167420 76712 167426 76724
rect 167546 76712 167552 76724
rect 167604 76712 167610 76764
rect 174262 76712 174268 76764
rect 174320 76752 174326 76764
rect 175182 76752 175188 76764
rect 174320 76724 175188 76752
rect 174320 76712 174326 76724
rect 175182 76712 175188 76724
rect 175240 76712 175246 76764
rect 176010 76712 176016 76764
rect 176068 76752 176074 76764
rect 176194 76752 176200 76764
rect 176068 76724 176200 76752
rect 176068 76712 176074 76724
rect 176194 76712 176200 76724
rect 176252 76712 176258 76764
rect 177206 76712 177212 76764
rect 177264 76752 177270 76764
rect 206646 76752 206652 76764
rect 177264 76724 206652 76752
rect 177264 76712 177270 76724
rect 206646 76712 206652 76724
rect 206704 76712 206710 76764
rect 159876 76656 160094 76684
rect 159876 76644 159882 76656
rect 160186 76644 160192 76696
rect 160244 76684 160250 76696
rect 160370 76684 160376 76696
rect 160244 76656 160376 76684
rect 160244 76644 160250 76656
rect 160370 76644 160376 76656
rect 160428 76644 160434 76696
rect 160830 76644 160836 76696
rect 160888 76684 160894 76696
rect 161290 76684 161296 76696
rect 160888 76656 161296 76684
rect 160888 76644 160894 76656
rect 161290 76644 161296 76656
rect 161348 76644 161354 76696
rect 161566 76644 161572 76696
rect 161624 76684 161630 76696
rect 161934 76684 161940 76696
rect 161624 76656 161940 76684
rect 161624 76644 161630 76656
rect 161934 76644 161940 76656
rect 161992 76644 161998 76696
rect 163222 76644 163228 76696
rect 163280 76684 163286 76696
rect 163406 76684 163412 76696
rect 163280 76656 163412 76684
rect 163280 76644 163286 76656
rect 163406 76644 163412 76656
rect 163464 76644 163470 76696
rect 164694 76644 164700 76696
rect 164752 76684 164758 76696
rect 165062 76684 165068 76696
rect 164752 76656 165068 76684
rect 164752 76644 164758 76656
rect 165062 76644 165068 76656
rect 165120 76644 165126 76696
rect 165890 76644 165896 76696
rect 165948 76684 165954 76696
rect 166074 76684 166080 76696
rect 165948 76656 166080 76684
rect 165948 76644 165954 76656
rect 166074 76644 166080 76656
rect 166132 76644 166138 76696
rect 167178 76644 167184 76696
rect 167236 76684 167242 76696
rect 167454 76684 167460 76696
rect 167236 76656 167460 76684
rect 167236 76644 167242 76656
rect 167454 76644 167460 76656
rect 167512 76644 167518 76696
rect 168558 76644 168564 76696
rect 168616 76684 168622 76696
rect 169110 76684 169116 76696
rect 168616 76656 169116 76684
rect 168616 76644 168622 76656
rect 169110 76644 169116 76656
rect 169168 76644 169174 76696
rect 171134 76644 171140 76696
rect 171192 76684 171198 76696
rect 171962 76684 171968 76696
rect 171192 76656 171968 76684
rect 171192 76644 171198 76656
rect 171962 76644 171968 76656
rect 172020 76644 172026 76696
rect 172422 76644 172428 76696
rect 172480 76684 172486 76696
rect 198090 76684 198096 76696
rect 172480 76656 198096 76684
rect 172480 76644 172486 76656
rect 198090 76644 198096 76656
rect 198148 76644 198154 76696
rect 215266 76684 215294 76792
rect 217318 76780 217324 76792
rect 217376 76820 217382 76832
rect 289814 76820 289820 76832
rect 217376 76792 289820 76820
rect 217376 76780 217382 76792
rect 289814 76780 289820 76792
rect 289872 76780 289878 76832
rect 217134 76712 217140 76764
rect 217192 76752 217198 76764
rect 296714 76752 296720 76764
rect 217192 76724 296720 76752
rect 217192 76712 217198 76724
rect 296714 76712 296720 76724
rect 296772 76712 296778 76764
rect 324314 76684 324320 76696
rect 215266 76656 324320 76684
rect 324314 76644 324320 76656
rect 324372 76644 324378 76696
rect 66254 76576 66260 76628
rect 66312 76616 66318 76628
rect 102134 76616 102140 76628
rect 66312 76588 102140 76616
rect 66312 76576 66318 76588
rect 102134 76576 102140 76588
rect 102192 76576 102198 76628
rect 113818 76576 113824 76628
rect 113876 76616 113882 76628
rect 141142 76616 141148 76628
rect 113876 76588 141148 76616
rect 113876 76576 113882 76588
rect 141142 76576 141148 76588
rect 141200 76576 141206 76628
rect 147306 76576 147312 76628
rect 147364 76616 147370 76628
rect 181438 76616 181444 76628
rect 147364 76588 181444 76616
rect 147364 76576 147370 76588
rect 181438 76576 181444 76588
rect 181496 76576 181502 76628
rect 189258 76576 189264 76628
rect 189316 76616 189322 76628
rect 189718 76616 189724 76628
rect 189316 76588 189724 76616
rect 189316 76576 189322 76588
rect 189718 76576 189724 76588
rect 189776 76616 189782 76628
rect 353294 76616 353300 76628
rect 189776 76588 353300 76616
rect 189776 76576 189782 76588
rect 353294 76576 353300 76588
rect 353352 76576 353358 76628
rect 59354 76508 59360 76560
rect 59412 76548 59418 76560
rect 102962 76548 102968 76560
rect 59412 76520 102968 76548
rect 59412 76508 59418 76520
rect 102962 76508 102968 76520
rect 103020 76548 103026 76560
rect 103020 76520 103514 76548
rect 103020 76508 103026 76520
rect 103486 76344 103514 76520
rect 114554 76508 114560 76560
rect 114612 76548 114618 76560
rect 132770 76548 132776 76560
rect 114612 76520 132776 76548
rect 114612 76508 114618 76520
rect 132770 76508 132776 76520
rect 132828 76508 132834 76560
rect 132954 76508 132960 76560
rect 133012 76548 133018 76560
rect 133782 76548 133788 76560
rect 133012 76520 133788 76548
rect 133012 76508 133018 76520
rect 133782 76508 133788 76520
rect 133840 76508 133846 76560
rect 135622 76508 135628 76560
rect 135680 76548 135686 76560
rect 136082 76548 136088 76560
rect 135680 76520 136088 76548
rect 135680 76508 135686 76520
rect 136082 76508 136088 76520
rect 136140 76508 136146 76560
rect 136634 76508 136640 76560
rect 136692 76548 136698 76560
rect 137462 76548 137468 76560
rect 136692 76520 137468 76548
rect 136692 76508 136698 76520
rect 137462 76508 137468 76520
rect 137520 76508 137526 76560
rect 146754 76508 146760 76560
rect 146812 76548 146818 76560
rect 184934 76548 184940 76560
rect 146812 76520 184940 76548
rect 146812 76508 146818 76520
rect 184934 76508 184940 76520
rect 184992 76508 184998 76560
rect 367094 76548 367100 76560
rect 190426 76520 367100 76548
rect 111702 76440 111708 76492
rect 111760 76480 111766 76492
rect 137646 76480 137652 76492
rect 111760 76452 137652 76480
rect 111760 76440 111766 76452
rect 137646 76440 137652 76452
rect 137704 76440 137710 76492
rect 154942 76440 154948 76492
rect 155000 76480 155006 76492
rect 155402 76480 155408 76492
rect 155000 76452 155408 76480
rect 155000 76440 155006 76452
rect 155402 76440 155408 76452
rect 155460 76440 155466 76492
rect 155954 76440 155960 76492
rect 156012 76480 156018 76492
rect 157058 76480 157064 76492
rect 156012 76452 157064 76480
rect 156012 76440 156018 76452
rect 157058 76440 157064 76452
rect 157116 76440 157122 76492
rect 158714 76440 158720 76492
rect 158772 76480 158778 76492
rect 159082 76480 159088 76492
rect 158772 76452 159088 76480
rect 158772 76440 158778 76452
rect 159082 76440 159088 76452
rect 159140 76440 159146 76492
rect 163222 76440 163228 76492
rect 163280 76480 163286 76492
rect 163958 76480 163964 76492
rect 163280 76452 163964 76480
rect 163280 76440 163286 76452
rect 163958 76440 163964 76452
rect 164016 76440 164022 76492
rect 164326 76440 164332 76492
rect 164384 76480 164390 76492
rect 164510 76480 164516 76492
rect 164384 76452 164516 76480
rect 164384 76440 164390 76452
rect 164510 76440 164516 76452
rect 164568 76440 164574 76492
rect 178586 76440 178592 76492
rect 178644 76480 178650 76492
rect 187694 76480 187700 76492
rect 178644 76452 187700 76480
rect 178644 76440 178650 76452
rect 187694 76440 187700 76452
rect 187752 76440 187758 76492
rect 110966 76372 110972 76424
rect 111024 76412 111030 76424
rect 126974 76412 126980 76424
rect 111024 76384 126980 76412
rect 111024 76372 111030 76384
rect 126974 76372 126980 76384
rect 127032 76372 127038 76424
rect 134334 76372 134340 76424
rect 134392 76412 134398 76424
rect 135162 76412 135168 76424
rect 134392 76384 135168 76412
rect 134392 76372 134398 76384
rect 135162 76372 135168 76384
rect 135220 76372 135226 76424
rect 135438 76372 135444 76424
rect 135496 76412 135502 76424
rect 136082 76412 136088 76424
rect 135496 76384 136088 76412
rect 135496 76372 135502 76384
rect 136082 76372 136088 76384
rect 136140 76372 136146 76424
rect 150434 76372 150440 76424
rect 150492 76412 150498 76424
rect 151262 76412 151268 76424
rect 150492 76384 151268 76412
rect 150492 76372 150498 76384
rect 151262 76372 151268 76384
rect 151320 76372 151326 76424
rect 163774 76372 163780 76424
rect 163832 76412 163838 76424
rect 166350 76412 166356 76424
rect 163832 76384 166356 76412
rect 163832 76372 163838 76384
rect 166350 76372 166356 76384
rect 166408 76372 166414 76424
rect 136818 76344 136824 76356
rect 103486 76316 136824 76344
rect 136818 76304 136824 76316
rect 136876 76304 136882 76356
rect 161014 76304 161020 76356
rect 161072 76344 161078 76356
rect 187418 76344 187424 76356
rect 161072 76316 187424 76344
rect 161072 76304 161078 76316
rect 187418 76304 187424 76316
rect 187476 76344 187482 76356
rect 190426 76344 190454 76520
rect 367094 76508 367100 76520
rect 367152 76508 367158 76560
rect 187476 76316 190454 76344
rect 187476 76304 187482 76316
rect 164510 76236 164516 76288
rect 164568 76276 164574 76288
rect 165430 76276 165436 76288
rect 164568 76248 165436 76276
rect 164568 76236 164574 76248
rect 165430 76236 165436 76248
rect 165488 76236 165494 76288
rect 166074 76236 166080 76288
rect 166132 76276 166138 76288
rect 166810 76276 166816 76288
rect 166132 76248 166816 76276
rect 166132 76236 166138 76248
rect 166810 76236 166816 76248
rect 166868 76236 166874 76288
rect 132770 76168 132776 76220
rect 132828 76208 132834 76220
rect 140866 76208 140872 76220
rect 132828 76180 140872 76208
rect 132828 76168 132834 76180
rect 140866 76168 140872 76180
rect 140924 76168 140930 76220
rect 171778 76100 171784 76152
rect 171836 76140 171842 76152
rect 172422 76140 172428 76152
rect 171836 76112 172428 76140
rect 171836 76100 171842 76112
rect 172422 76100 172428 76112
rect 172480 76100 172486 76152
rect 132770 76032 132776 76084
rect 132828 76072 132834 76084
rect 133598 76072 133604 76084
rect 132828 76044 133604 76072
rect 132828 76032 132834 76044
rect 133598 76032 133604 76044
rect 133656 76032 133662 76084
rect 144362 75964 144368 76016
rect 144420 76004 144426 76016
rect 146294 76004 146300 76016
rect 144420 75976 146300 76004
rect 144420 75964 144426 75976
rect 146294 75964 146300 75976
rect 146352 75964 146358 76016
rect 173342 75896 173348 75948
rect 173400 75936 173406 75948
rect 173618 75936 173624 75948
rect 173400 75908 173624 75936
rect 173400 75896 173406 75908
rect 173618 75896 173624 75908
rect 173676 75896 173682 75948
rect 177206 75896 177212 75948
rect 177264 75936 177270 75948
rect 177666 75936 177672 75948
rect 177264 75908 177672 75936
rect 177264 75896 177270 75908
rect 177666 75896 177672 75908
rect 177724 75896 177730 75948
rect 210510 75896 210516 75948
rect 210568 75936 210574 75948
rect 553394 75936 553400 75948
rect 210568 75908 553400 75936
rect 210568 75896 210574 75908
rect 553394 75896 553400 75908
rect 553452 75896 553458 75948
rect 103054 75828 103060 75880
rect 103112 75868 103118 75880
rect 103112 75840 139992 75868
rect 103112 75828 103118 75840
rect 103882 75760 103888 75812
rect 103940 75800 103946 75812
rect 104066 75800 104072 75812
rect 103940 75772 104072 75800
rect 103940 75760 103946 75772
rect 104066 75760 104072 75772
rect 104124 75800 104130 75812
rect 138934 75800 138940 75812
rect 104124 75772 138940 75800
rect 104124 75760 104130 75772
rect 138934 75760 138940 75772
rect 138992 75760 138998 75812
rect 139964 75800 139992 75840
rect 140038 75828 140044 75880
rect 140096 75868 140102 75880
rect 140222 75868 140228 75880
rect 140096 75840 140228 75868
rect 140096 75828 140102 75840
rect 140222 75828 140228 75840
rect 140280 75828 140286 75880
rect 166626 75828 166632 75880
rect 166684 75868 166690 75880
rect 200758 75868 200764 75880
rect 166684 75840 200764 75868
rect 166684 75828 166690 75840
rect 200758 75828 200764 75840
rect 200816 75828 200822 75880
rect 144822 75800 144828 75812
rect 139964 75772 144828 75800
rect 144822 75760 144828 75772
rect 144880 75760 144886 75812
rect 157306 75772 169754 75800
rect 111886 75692 111892 75744
rect 111944 75732 111950 75744
rect 111944 75704 138014 75732
rect 111944 75692 111950 75704
rect 100754 75624 100760 75676
rect 100812 75664 100818 75676
rect 101214 75664 101220 75676
rect 100812 75636 101220 75664
rect 100812 75624 100818 75636
rect 101214 75624 101220 75636
rect 101272 75664 101278 75676
rect 135070 75664 135076 75676
rect 101272 75636 135076 75664
rect 101272 75624 101278 75636
rect 135070 75624 135076 75636
rect 135128 75624 135134 75676
rect 135346 75624 135352 75676
rect 135404 75664 135410 75676
rect 135898 75664 135904 75676
rect 135404 75636 135904 75664
rect 135404 75624 135410 75636
rect 135898 75624 135904 75636
rect 135956 75624 135962 75676
rect 104434 75556 104440 75608
rect 104492 75596 104498 75608
rect 137554 75596 137560 75608
rect 104492 75568 137560 75596
rect 104492 75556 104498 75568
rect 137554 75556 137560 75568
rect 137612 75556 137618 75608
rect 137986 75596 138014 75704
rect 138198 75692 138204 75744
rect 138256 75732 138262 75744
rect 139210 75732 139216 75744
rect 138256 75704 139216 75732
rect 138256 75692 138262 75704
rect 139210 75692 139216 75704
rect 139268 75692 139274 75744
rect 139762 75692 139768 75744
rect 139820 75732 139826 75744
rect 140222 75732 140228 75744
rect 139820 75704 140228 75732
rect 139820 75692 139826 75704
rect 140222 75692 140228 75704
rect 140280 75692 140286 75744
rect 142522 75624 142528 75676
rect 142580 75664 142586 75676
rect 142798 75664 142804 75676
rect 142580 75636 142804 75664
rect 142580 75624 142586 75636
rect 142798 75624 142804 75636
rect 142856 75624 142862 75676
rect 137986 75568 144224 75596
rect 93854 75488 93860 75540
rect 93912 75528 93918 75540
rect 105262 75528 105268 75540
rect 93912 75500 105268 75528
rect 93912 75488 93918 75500
rect 105262 75488 105268 75500
rect 105320 75488 105326 75540
rect 116578 75488 116584 75540
rect 116636 75528 116642 75540
rect 116636 75500 142844 75528
rect 116636 75488 116642 75500
rect 104250 75420 104256 75472
rect 104308 75460 104314 75472
rect 131022 75460 131028 75472
rect 104308 75432 131028 75460
rect 104308 75420 104314 75432
rect 131022 75420 131028 75432
rect 131080 75420 131086 75472
rect 131114 75420 131120 75472
rect 131172 75460 131178 75472
rect 132586 75460 132592 75472
rect 131172 75432 132592 75460
rect 131172 75420 131178 75432
rect 132586 75420 132592 75432
rect 132644 75420 132650 75472
rect 85574 75352 85580 75404
rect 85632 75392 85638 75404
rect 103882 75392 103888 75404
rect 85632 75364 103888 75392
rect 85632 75352 85638 75364
rect 103882 75352 103888 75364
rect 103940 75352 103946 75404
rect 117222 75352 117228 75404
rect 117280 75392 117286 75404
rect 142816 75392 142844 75500
rect 144196 75460 144224 75568
rect 146478 75556 146484 75608
rect 146536 75596 146542 75608
rect 157306 75596 157334 75772
rect 146536 75568 157334 75596
rect 146536 75556 146542 75568
rect 158622 75556 158628 75608
rect 158680 75596 158686 75608
rect 169726 75596 169754 75772
rect 175090 75760 175096 75812
rect 175148 75800 175154 75812
rect 204898 75800 204904 75812
rect 175148 75772 204904 75800
rect 175148 75760 175154 75772
rect 204898 75760 204904 75772
rect 204956 75760 204962 75812
rect 172974 75692 172980 75744
rect 173032 75732 173038 75744
rect 207566 75732 207572 75744
rect 173032 75704 207572 75732
rect 173032 75692 173038 75704
rect 207566 75692 207572 75704
rect 207624 75732 207630 75744
rect 208302 75732 208308 75744
rect 207624 75704 208308 75732
rect 207624 75692 207630 75704
rect 208302 75692 208308 75704
rect 208360 75692 208366 75744
rect 170582 75624 170588 75676
rect 170640 75664 170646 75676
rect 171042 75664 171048 75676
rect 170640 75636 171048 75664
rect 170640 75624 170646 75636
rect 171042 75624 171048 75636
rect 171100 75664 171106 75676
rect 204714 75664 204720 75676
rect 171100 75636 204720 75664
rect 171100 75624 171106 75636
rect 204714 75624 204720 75636
rect 204772 75624 204778 75676
rect 180794 75596 180800 75608
rect 158680 75568 160094 75596
rect 169726 75568 180800 75596
rect 158680 75556 158686 75568
rect 144822 75488 144828 75540
rect 144880 75528 144886 75540
rect 147030 75528 147036 75540
rect 144880 75500 147036 75528
rect 144880 75488 144886 75500
rect 147030 75488 147036 75500
rect 147088 75488 147094 75540
rect 154574 75488 154580 75540
rect 154632 75528 154638 75540
rect 155494 75528 155500 75540
rect 154632 75500 155500 75528
rect 154632 75488 154638 75500
rect 155494 75488 155500 75500
rect 155552 75488 155558 75540
rect 156138 75488 156144 75540
rect 156196 75528 156202 75540
rect 156782 75528 156788 75540
rect 156196 75500 156788 75528
rect 156196 75488 156202 75500
rect 156782 75488 156788 75500
rect 156840 75488 156846 75540
rect 160066 75528 160094 75568
rect 180794 75556 180800 75568
rect 180852 75556 180858 75608
rect 179966 75528 179972 75540
rect 160066 75500 179972 75528
rect 179966 75488 179972 75500
rect 180024 75488 180030 75540
rect 180702 75488 180708 75540
rect 180760 75528 180766 75540
rect 216674 75528 216680 75540
rect 180760 75500 216680 75528
rect 180760 75488 180766 75500
rect 216674 75488 216680 75500
rect 216732 75488 216738 75540
rect 146662 75460 146668 75472
rect 144196 75432 146668 75460
rect 146662 75420 146668 75432
rect 146720 75460 146726 75472
rect 176746 75460 176752 75472
rect 146720 75432 176752 75460
rect 146720 75420 146726 75432
rect 176746 75420 176752 75432
rect 176804 75420 176810 75472
rect 176930 75420 176936 75472
rect 176988 75460 176994 75472
rect 177114 75460 177120 75472
rect 176988 75432 177120 75460
rect 176988 75420 176994 75432
rect 177114 75420 177120 75432
rect 177172 75420 177178 75472
rect 117280 75364 138014 75392
rect 142816 75364 145880 75392
rect 117280 75352 117286 75364
rect 99006 75284 99012 75336
rect 99064 75324 99070 75336
rect 131114 75324 131120 75336
rect 99064 75296 131120 75324
rect 99064 75284 99070 75296
rect 131114 75284 131120 75296
rect 131172 75284 131178 75336
rect 137002 75284 137008 75336
rect 137060 75324 137066 75336
rect 137186 75324 137192 75336
rect 137060 75296 137192 75324
rect 137060 75284 137066 75296
rect 137186 75284 137192 75296
rect 137244 75284 137250 75336
rect 137986 75324 138014 75364
rect 145466 75324 145472 75336
rect 137986 75296 145472 75324
rect 145466 75284 145472 75296
rect 145524 75284 145530 75336
rect 71038 75216 71044 75268
rect 71096 75256 71102 75268
rect 104434 75256 104440 75268
rect 71096 75228 104440 75256
rect 71096 75216 71102 75228
rect 104434 75216 104440 75228
rect 104492 75216 104498 75268
rect 118602 75216 118608 75268
rect 118660 75256 118666 75268
rect 138014 75256 138020 75268
rect 118660 75228 138020 75256
rect 118660 75216 118666 75228
rect 138014 75216 138020 75228
rect 138072 75216 138078 75268
rect 138106 75216 138112 75268
rect 138164 75256 138170 75268
rect 138474 75256 138480 75268
rect 138164 75228 138480 75256
rect 138164 75216 138170 75228
rect 138474 75216 138480 75228
rect 138532 75216 138538 75268
rect 141234 75216 141240 75268
rect 141292 75256 141298 75268
rect 141602 75256 141608 75268
rect 141292 75228 141608 75256
rect 141292 75216 141298 75228
rect 141602 75216 141608 75228
rect 141660 75216 141666 75268
rect 142890 75216 142896 75268
rect 142948 75256 142954 75268
rect 143350 75256 143356 75268
rect 142948 75228 143356 75256
rect 142948 75216 142954 75228
rect 143350 75216 143356 75228
rect 143408 75216 143414 75268
rect 143902 75216 143908 75268
rect 143960 75256 143966 75268
rect 144086 75256 144092 75268
rect 143960 75228 144092 75256
rect 143960 75216 143966 75228
rect 144086 75216 144092 75228
rect 144144 75216 144150 75268
rect 145190 75216 145196 75268
rect 145248 75256 145254 75268
rect 145742 75256 145748 75268
rect 145248 75228 145748 75256
rect 145248 75216 145254 75228
rect 145742 75216 145748 75228
rect 145800 75216 145806 75268
rect 35894 75148 35900 75200
rect 35952 75188 35958 75200
rect 100754 75188 100760 75200
rect 35952 75160 100760 75188
rect 35952 75148 35958 75160
rect 100754 75148 100760 75160
rect 100812 75148 100818 75200
rect 112438 75148 112444 75200
rect 112496 75188 112502 75200
rect 112496 75160 138336 75188
rect 112496 75148 112502 75160
rect 97902 75080 97908 75132
rect 97960 75120 97966 75132
rect 114554 75120 114560 75132
rect 97960 75092 114560 75120
rect 97960 75080 97966 75092
rect 114554 75080 114560 75092
rect 114612 75080 114618 75132
rect 121086 75080 121092 75132
rect 121144 75120 121150 75132
rect 138308 75120 138336 75160
rect 141142 75148 141148 75200
rect 141200 75188 141206 75200
rect 141970 75188 141976 75200
rect 141200 75160 141976 75188
rect 141200 75148 141206 75160
rect 141970 75148 141976 75160
rect 142028 75148 142034 75200
rect 142706 75148 142712 75200
rect 142764 75188 142770 75200
rect 143166 75188 143172 75200
rect 142764 75160 143172 75188
rect 142764 75148 142770 75160
rect 143166 75148 143172 75160
rect 143224 75148 143230 75200
rect 145852 75188 145880 75364
rect 151078 75352 151084 75404
rect 151136 75392 151142 75404
rect 216674 75392 216680 75404
rect 151136 75364 216680 75392
rect 151136 75352 151142 75364
rect 216674 75352 216680 75364
rect 216732 75352 216738 75404
rect 149698 75284 149704 75336
rect 149756 75324 149762 75336
rect 187694 75324 187700 75336
rect 149756 75296 187700 75324
rect 149756 75284 149762 75296
rect 187694 75284 187700 75296
rect 187752 75284 187758 75336
rect 191742 75284 191748 75336
rect 191800 75324 191806 75336
rect 304994 75324 305000 75336
rect 191800 75296 305000 75324
rect 191800 75284 191806 75296
rect 304994 75284 305000 75296
rect 305052 75284 305058 75336
rect 147490 75216 147496 75268
rect 147548 75256 147554 75268
rect 193858 75256 193864 75268
rect 147548 75228 193864 75256
rect 147548 75216 147554 75228
rect 193858 75216 193864 75228
rect 193916 75216 193922 75268
rect 204898 75216 204904 75268
rect 204956 75256 204962 75268
rect 442258 75256 442264 75268
rect 204956 75228 442264 75256
rect 204956 75216 204962 75228
rect 442258 75216 442264 75228
rect 442316 75216 442322 75268
rect 148042 75188 148048 75200
rect 145852 75160 148048 75188
rect 148042 75148 148048 75160
rect 148100 75188 148106 75200
rect 148100 75160 150894 75188
rect 148100 75148 148106 75160
rect 140958 75120 140964 75132
rect 121144 75092 138014 75120
rect 138308 75092 140964 75120
rect 121144 75080 121150 75092
rect 108574 75012 108580 75064
rect 108632 75052 108638 75064
rect 108632 75024 128354 75052
rect 108632 75012 108638 75024
rect 128326 74984 128354 75024
rect 130562 75012 130568 75064
rect 130620 75052 130626 75064
rect 130930 75052 130936 75064
rect 130620 75024 130936 75052
rect 130620 75012 130626 75024
rect 130930 75012 130936 75024
rect 130988 75012 130994 75064
rect 137986 75052 138014 75092
rect 140958 75080 140964 75092
rect 141016 75080 141022 75132
rect 142430 75080 142436 75132
rect 142488 75120 142494 75132
rect 143258 75120 143264 75132
rect 142488 75092 143264 75120
rect 142488 75080 142494 75092
rect 143258 75080 143264 75092
rect 143316 75080 143322 75132
rect 149330 75080 149336 75132
rect 149388 75120 149394 75132
rect 149974 75120 149980 75132
rect 149388 75092 149980 75120
rect 149388 75080 149394 75092
rect 149974 75080 149980 75092
rect 150032 75080 150038 75132
rect 150866 75120 150894 75160
rect 151998 75148 152004 75200
rect 152056 75188 152062 75200
rect 153010 75188 153016 75200
rect 152056 75160 153016 75188
rect 152056 75148 152062 75160
rect 153010 75148 153016 75160
rect 153068 75148 153074 75200
rect 156046 75148 156052 75200
rect 156104 75188 156110 75200
rect 156966 75188 156972 75200
rect 156104 75160 156972 75188
rect 156104 75148 156110 75160
rect 156966 75148 156972 75160
rect 157024 75148 157030 75200
rect 201678 75188 201684 75200
rect 157306 75160 201684 75188
rect 157306 75120 157334 75160
rect 201678 75148 201684 75160
rect 201736 75148 201742 75200
rect 208302 75148 208308 75200
rect 208360 75188 208366 75200
rect 521654 75188 521660 75200
rect 208360 75160 521660 75188
rect 208360 75148 208366 75160
rect 521654 75148 521660 75160
rect 521712 75148 521718 75200
rect 150866 75092 157334 75120
rect 158714 75080 158720 75132
rect 158772 75120 158778 75132
rect 160002 75120 160008 75132
rect 158772 75092 160008 75120
rect 158772 75080 158778 75092
rect 160002 75080 160008 75092
rect 160060 75080 160066 75132
rect 165706 75080 165712 75132
rect 165764 75120 165770 75132
rect 189626 75120 189632 75132
rect 165764 75092 189632 75120
rect 165764 75080 165770 75092
rect 189626 75080 189632 75092
rect 189684 75080 189690 75132
rect 146570 75052 146576 75064
rect 137986 75024 146576 75052
rect 146570 75012 146576 75024
rect 146628 75012 146634 75064
rect 151630 75012 151636 75064
rect 151688 75052 151694 75064
rect 151814 75052 151820 75064
rect 151688 75024 151820 75052
rect 151688 75012 151694 75024
rect 151814 75012 151820 75024
rect 151872 75012 151878 75064
rect 154666 75012 154672 75064
rect 154724 75052 154730 75064
rect 155586 75052 155592 75064
rect 154724 75024 155592 75052
rect 154724 75012 154730 75024
rect 155586 75012 155592 75024
rect 155644 75012 155650 75064
rect 158898 75012 158904 75064
rect 158956 75052 158962 75064
rect 159910 75052 159916 75064
rect 158956 75024 159916 75052
rect 158956 75012 158962 75024
rect 159910 75012 159916 75024
rect 159968 75012 159974 75064
rect 191374 75052 191380 75064
rect 160066 75024 191380 75052
rect 131298 74984 131304 74996
rect 128326 74956 131304 74984
rect 131298 74944 131304 74956
rect 131356 74984 131362 74996
rect 131356 74956 136220 74984
rect 131356 74944 131362 74956
rect 136192 74916 136220 74956
rect 137002 74944 137008 74996
rect 137060 74984 137066 74996
rect 137738 74984 137744 74996
rect 137060 74956 137744 74984
rect 137060 74944 137066 74956
rect 137738 74944 137744 74956
rect 137796 74944 137802 74996
rect 138014 74944 138020 74996
rect 138072 74984 138078 74996
rect 145190 74984 145196 74996
rect 138072 74956 145196 74984
rect 138072 74944 138078 74956
rect 145190 74944 145196 74956
rect 145248 74944 145254 74996
rect 139302 74916 139308 74928
rect 136192 74888 139308 74916
rect 139302 74876 139308 74888
rect 139360 74876 139366 74928
rect 143718 74876 143724 74928
rect 143776 74916 143782 74928
rect 144730 74916 144736 74928
rect 143776 74888 144736 74916
rect 143776 74876 143782 74888
rect 144730 74876 144736 74888
rect 144788 74876 144794 74928
rect 131022 74808 131028 74860
rect 131080 74848 131086 74860
rect 135346 74848 135352 74860
rect 131080 74820 135352 74848
rect 131080 74808 131086 74820
rect 135346 74808 135352 74820
rect 135404 74808 135410 74860
rect 156322 74808 156328 74860
rect 156380 74848 156386 74860
rect 160066 74848 160094 75024
rect 191374 75012 191380 75024
rect 191432 75052 191438 75064
rect 191742 75052 191748 75064
rect 191432 75024 191748 75052
rect 191432 75012 191438 75024
rect 191742 75012 191748 75024
rect 191800 75012 191806 75064
rect 173158 74944 173164 74996
rect 173216 74984 173222 74996
rect 173526 74984 173532 74996
rect 173216 74956 173532 74984
rect 173216 74944 173222 74956
rect 173526 74944 173532 74956
rect 173584 74944 173590 74996
rect 176746 74944 176752 74996
rect 176804 74984 176810 74996
rect 185026 74984 185032 74996
rect 176804 74956 185032 74984
rect 176804 74944 176810 74956
rect 185026 74944 185032 74956
rect 185084 74944 185090 74996
rect 210786 74984 210792 74996
rect 185136 74956 210792 74984
rect 181990 74876 181996 74928
rect 182048 74916 182054 74928
rect 185136 74916 185164 74956
rect 210786 74944 210792 74956
rect 210844 74944 210850 74996
rect 211338 74916 211344 74928
rect 182048 74888 185164 74916
rect 186286 74888 211344 74916
rect 182048 74876 182054 74888
rect 156380 74820 160094 74848
rect 156380 74808 156386 74820
rect 173066 74808 173072 74860
rect 173124 74848 173130 74860
rect 177942 74848 177948 74860
rect 173124 74820 177948 74848
rect 173124 74808 173130 74820
rect 177942 74808 177948 74820
rect 178000 74848 178006 74860
rect 186286 74848 186314 74888
rect 211338 74876 211344 74888
rect 211396 74876 211402 74928
rect 178000 74820 186314 74848
rect 178000 74808 178006 74820
rect 161750 74740 161756 74792
rect 161808 74780 161814 74792
rect 162670 74780 162676 74792
rect 161808 74752 162676 74780
rect 161808 74740 161814 74752
rect 162670 74740 162676 74752
rect 162728 74740 162734 74792
rect 130654 74672 130660 74724
rect 130712 74712 130718 74724
rect 131022 74712 131028 74724
rect 130712 74684 131028 74712
rect 130712 74672 130718 74684
rect 131022 74672 131028 74684
rect 131080 74672 131086 74724
rect 167086 74536 167092 74588
rect 167144 74576 167150 74588
rect 167730 74576 167736 74588
rect 167144 74548 167736 74576
rect 167144 74536 167150 74548
rect 167730 74536 167736 74548
rect 167788 74536 167794 74588
rect 128538 74468 128544 74520
rect 128596 74508 128602 74520
rect 139578 74508 139584 74520
rect 128596 74480 139584 74508
rect 128596 74468 128602 74480
rect 139578 74468 139584 74480
rect 139636 74468 139642 74520
rect 142246 74468 142252 74520
rect 142304 74508 142310 74520
rect 143074 74508 143080 74520
rect 142304 74480 143080 74508
rect 142304 74468 142310 74480
rect 143074 74468 143080 74480
rect 143132 74468 143138 74520
rect 152642 74468 152648 74520
rect 152700 74508 152706 74520
rect 218330 74508 218336 74520
rect 152700 74480 218336 74508
rect 152700 74468 152706 74480
rect 218330 74468 218336 74480
rect 218388 74468 218394 74520
rect 119430 74400 119436 74452
rect 119488 74440 119494 74452
rect 153838 74440 153844 74452
rect 119488 74412 153844 74440
rect 119488 74400 119494 74412
rect 153838 74400 153844 74412
rect 153896 74400 153902 74452
rect 159634 74400 159640 74452
rect 159692 74440 159698 74452
rect 218146 74440 218152 74452
rect 159692 74412 218152 74440
rect 159692 74400 159698 74412
rect 218146 74400 218152 74412
rect 218204 74400 218210 74452
rect 106734 74332 106740 74384
rect 106792 74372 106798 74384
rect 140590 74372 140596 74384
rect 106792 74344 140596 74372
rect 106792 74332 106798 74344
rect 140590 74332 140596 74344
rect 140648 74332 140654 74384
rect 153746 74332 153752 74384
rect 153804 74372 153810 74384
rect 154482 74372 154488 74384
rect 153804 74344 154488 74372
rect 153804 74332 153810 74344
rect 154482 74332 154488 74344
rect 154540 74332 154546 74384
rect 156230 74332 156236 74384
rect 156288 74372 156294 74384
rect 188522 74372 188528 74384
rect 156288 74344 188528 74372
rect 156288 74332 156294 74344
rect 188522 74332 188528 74344
rect 188580 74332 188586 74384
rect 115382 74264 115388 74316
rect 115440 74304 115446 74316
rect 147858 74304 147864 74316
rect 115440 74276 147864 74304
rect 115440 74264 115446 74276
rect 147858 74264 147864 74276
rect 147916 74304 147922 74316
rect 148686 74304 148692 74316
rect 147916 74276 148692 74304
rect 147916 74264 147922 74276
rect 148686 74264 148692 74276
rect 148744 74264 148750 74316
rect 165062 74264 165068 74316
rect 165120 74304 165126 74316
rect 165706 74304 165712 74316
rect 165120 74276 165712 74304
rect 165120 74264 165126 74276
rect 165706 74264 165712 74276
rect 165764 74264 165770 74316
rect 168282 74264 168288 74316
rect 168340 74304 168346 74316
rect 202322 74304 202328 74316
rect 168340 74276 202328 74304
rect 168340 74264 168346 74276
rect 202322 74264 202328 74276
rect 202380 74264 202386 74316
rect 109954 74196 109960 74248
rect 110012 74236 110018 74248
rect 142522 74236 142528 74248
rect 110012 74208 142528 74236
rect 110012 74196 110018 74208
rect 142522 74196 142528 74208
rect 142580 74196 142586 74248
rect 153838 74196 153844 74248
rect 153896 74236 153902 74248
rect 154390 74236 154396 74248
rect 153896 74208 154396 74236
rect 153896 74196 153902 74208
rect 154390 74196 154396 74208
rect 154448 74196 154454 74248
rect 155862 74196 155868 74248
rect 155920 74236 155926 74248
rect 156966 74236 156972 74248
rect 155920 74208 156972 74236
rect 155920 74196 155926 74208
rect 156966 74196 156972 74208
rect 157024 74236 157030 74248
rect 157024 74208 157334 74236
rect 157024 74196 157030 74208
rect 108482 74128 108488 74180
rect 108540 74168 108546 74180
rect 140406 74168 140412 74180
rect 108540 74140 140412 74168
rect 108540 74128 108546 74140
rect 140406 74128 140412 74140
rect 140464 74128 140470 74180
rect 149146 74128 149152 74180
rect 149204 74168 149210 74180
rect 156782 74168 156788 74180
rect 149204 74140 156788 74168
rect 149204 74128 149210 74140
rect 156782 74128 156788 74140
rect 156840 74128 156846 74180
rect 157306 74168 157334 74208
rect 159450 74196 159456 74248
rect 159508 74236 159514 74248
rect 194042 74236 194048 74248
rect 159508 74208 194048 74236
rect 159508 74196 159514 74208
rect 194042 74196 194048 74208
rect 194100 74196 194106 74248
rect 189074 74168 189080 74180
rect 157306 74140 189080 74168
rect 189074 74128 189080 74140
rect 189132 74128 189138 74180
rect 218238 74128 218244 74180
rect 218296 74168 218302 74180
rect 218606 74168 218612 74180
rect 218296 74140 218612 74168
rect 218296 74128 218302 74140
rect 218606 74128 218612 74140
rect 218664 74128 218670 74180
rect 121178 74060 121184 74112
rect 121236 74100 121242 74112
rect 152918 74100 152924 74112
rect 121236 74072 152924 74100
rect 121236 74060 121242 74072
rect 152918 74060 152924 74072
rect 152976 74060 152982 74112
rect 163130 74060 163136 74112
rect 163188 74100 163194 74112
rect 163866 74100 163872 74112
rect 163188 74072 163872 74100
rect 163188 74060 163194 74072
rect 163866 74060 163872 74072
rect 163924 74060 163930 74112
rect 165706 74060 165712 74112
rect 165764 74100 165770 74112
rect 166534 74100 166540 74112
rect 165764 74072 166540 74100
rect 165764 74060 165770 74072
rect 166534 74060 166540 74072
rect 166592 74060 166598 74112
rect 167270 74060 167276 74112
rect 167328 74100 167334 74112
rect 168190 74100 168196 74112
rect 167328 74072 168196 74100
rect 167328 74060 167334 74072
rect 168190 74060 168196 74072
rect 168248 74060 168254 74112
rect 196986 74100 196992 74112
rect 169726 74072 196992 74100
rect 119062 73992 119068 74044
rect 119120 74032 119126 74044
rect 151630 74032 151636 74044
rect 119120 74004 151636 74032
rect 119120 73992 119126 74004
rect 151630 73992 151636 74004
rect 151688 73992 151694 74044
rect 159726 73992 159732 74044
rect 159784 74032 159790 74044
rect 159910 74032 159916 74044
rect 159784 74004 159916 74032
rect 159784 73992 159790 74004
rect 159910 73992 159916 74004
rect 159968 73992 159974 74044
rect 164142 73992 164148 74044
rect 164200 74032 164206 74044
rect 169726 74032 169754 74072
rect 196986 74060 196992 74072
rect 197044 74060 197050 74112
rect 164200 74004 169754 74032
rect 164200 73992 164206 74004
rect 175274 73992 175280 74044
rect 175332 74032 175338 74044
rect 206370 74032 206376 74044
rect 175332 74004 206376 74032
rect 175332 73992 175338 74004
rect 206370 73992 206376 74004
rect 206428 73992 206434 74044
rect 218330 73992 218336 74044
rect 218388 74032 218394 74044
rect 255314 74032 255320 74044
rect 218388 74004 255320 74032
rect 218388 73992 218394 74004
rect 255314 73992 255320 74004
rect 255372 73992 255378 74044
rect 111334 73924 111340 73976
rect 111392 73964 111398 73976
rect 142246 73964 142252 73976
rect 111392 73936 142252 73964
rect 111392 73924 111398 73936
rect 142246 73924 142252 73936
rect 142304 73924 142310 73976
rect 158530 73924 158536 73976
rect 158588 73964 158594 73976
rect 159818 73964 159824 73976
rect 158588 73936 159824 73964
rect 158588 73924 158594 73936
rect 159818 73924 159824 73936
rect 159876 73924 159882 73976
rect 163498 73924 163504 73976
rect 163556 73964 163562 73976
rect 168190 73964 168196 73976
rect 163556 73936 168196 73964
rect 163556 73924 163562 73936
rect 168190 73924 168196 73936
rect 168248 73924 168254 73976
rect 170214 73924 170220 73976
rect 170272 73964 170278 73976
rect 180518 73964 180524 73976
rect 170272 73936 180524 73964
rect 170272 73924 170278 73936
rect 180518 73924 180524 73936
rect 180576 73924 180582 73976
rect 188522 73924 188528 73976
rect 188580 73964 188586 73976
rect 261478 73964 261484 73976
rect 188580 73936 261484 73964
rect 188580 73924 188586 73936
rect 261478 73924 261484 73936
rect 261536 73924 261542 73976
rect 89714 73856 89720 73908
rect 89772 73896 89778 73908
rect 89772 73868 103514 73896
rect 89772 73856 89778 73868
rect 8938 73788 8944 73840
rect 8996 73828 9002 73840
rect 8996 73800 84194 73828
rect 8996 73788 9002 73800
rect 84166 73692 84194 73800
rect 103486 73760 103514 73868
rect 119338 73856 119344 73908
rect 119396 73896 119402 73908
rect 149238 73896 149244 73908
rect 119396 73868 149244 73896
rect 119396 73856 119402 73868
rect 149238 73856 149244 73868
rect 149296 73896 149302 73908
rect 149974 73896 149980 73908
rect 149296 73868 149980 73896
rect 149296 73856 149302 73868
rect 149974 73856 149980 73868
rect 150032 73856 150038 73908
rect 173710 73856 173716 73908
rect 173768 73896 173774 73908
rect 203610 73896 203616 73908
rect 173768 73868 203616 73896
rect 173768 73856 173774 73868
rect 203610 73856 203616 73868
rect 203668 73856 203674 73908
rect 218146 73856 218152 73908
rect 218204 73896 218210 73908
rect 347774 73896 347780 73908
rect 218204 73868 347780 73896
rect 218204 73856 218210 73868
rect 347774 73856 347780 73868
rect 347832 73856 347838 73908
rect 107194 73788 107200 73840
rect 107252 73828 107258 73840
rect 136358 73828 136364 73840
rect 107252 73800 136364 73828
rect 107252 73788 107258 73800
rect 136358 73788 136364 73800
rect 136416 73788 136422 73840
rect 159358 73788 159364 73840
rect 159416 73828 159422 73840
rect 160002 73828 160008 73840
rect 159416 73800 160008 73828
rect 159416 73788 159422 73800
rect 160002 73788 160008 73800
rect 160060 73788 160066 73840
rect 162210 73788 162216 73840
rect 162268 73828 162274 73840
rect 192938 73828 192944 73840
rect 162268 73800 192944 73828
rect 162268 73788 162274 73800
rect 192938 73788 192944 73800
rect 192996 73828 193002 73840
rect 322934 73828 322940 73840
rect 192996 73800 322940 73828
rect 192996 73788 193002 73800
rect 322934 73788 322940 73800
rect 322992 73788 322998 73840
rect 104342 73760 104348 73772
rect 103486 73732 104348 73760
rect 104342 73720 104348 73732
rect 104400 73760 104406 73772
rect 139118 73760 139124 73772
rect 104400 73732 139124 73760
rect 104400 73720 104406 73732
rect 139118 73720 139124 73732
rect 139176 73720 139182 73772
rect 157978 73720 157984 73772
rect 158036 73760 158042 73772
rect 158530 73760 158536 73772
rect 158036 73732 158536 73760
rect 158036 73720 158042 73732
rect 158530 73720 158536 73732
rect 158588 73720 158594 73772
rect 180518 73720 180524 73772
rect 180576 73760 180582 73772
rect 208854 73760 208860 73772
rect 180576 73732 208860 73760
rect 180576 73720 180582 73732
rect 208854 73720 208860 73732
rect 208912 73720 208918 73772
rect 105906 73692 105912 73704
rect 84166 73664 105912 73692
rect 105906 73652 105912 73664
rect 105964 73692 105970 73704
rect 132402 73692 132408 73704
rect 105964 73664 132408 73692
rect 105964 73652 105970 73664
rect 132402 73652 132408 73664
rect 132460 73652 132466 73704
rect 179046 73652 179052 73704
rect 179104 73692 179110 73704
rect 201494 73692 201500 73704
rect 179104 73664 201500 73692
rect 179104 73652 179110 73664
rect 201494 73652 201500 73664
rect 201552 73652 201558 73704
rect 122006 73584 122012 73636
rect 122064 73624 122070 73636
rect 128446 73624 128452 73636
rect 122064 73596 128452 73624
rect 122064 73584 122070 73596
rect 128446 73584 128452 73596
rect 128504 73624 128510 73636
rect 129642 73624 129648 73636
rect 128504 73596 129648 73624
rect 128504 73584 128510 73596
rect 129642 73584 129648 73596
rect 129700 73584 129706 73636
rect 152274 73584 152280 73636
rect 152332 73624 152338 73636
rect 153010 73624 153016 73636
rect 152332 73596 153016 73624
rect 152332 73584 152338 73596
rect 153010 73584 153016 73596
rect 153068 73584 153074 73636
rect 162118 73584 162124 73636
rect 162176 73624 162182 73636
rect 167914 73624 167920 73636
rect 162176 73596 167920 73624
rect 162176 73584 162182 73596
rect 167914 73584 167920 73596
rect 167972 73584 167978 73636
rect 106274 73176 106280 73228
rect 106332 73216 106338 73228
rect 106734 73216 106740 73228
rect 106332 73188 106740 73216
rect 106332 73176 106338 73188
rect 106734 73176 106740 73188
rect 106792 73176 106798 73228
rect 107654 73176 107660 73228
rect 107712 73216 107718 73228
rect 108482 73216 108488 73228
rect 107712 73188 108488 73216
rect 107712 73176 107718 73188
rect 108482 73176 108488 73188
rect 108540 73176 108546 73228
rect 121362 73108 121368 73160
rect 121420 73148 121426 73160
rect 149606 73148 149612 73160
rect 121420 73120 149612 73148
rect 121420 73108 121426 73120
rect 149606 73108 149612 73120
rect 149664 73148 149670 73160
rect 149882 73148 149888 73160
rect 149664 73120 149888 73148
rect 149664 73108 149670 73120
rect 149882 73108 149888 73120
rect 149940 73108 149946 73160
rect 161106 73108 161112 73160
rect 161164 73148 161170 73160
rect 195238 73148 195244 73160
rect 161164 73120 195244 73148
rect 161164 73108 161170 73120
rect 195238 73108 195244 73120
rect 195296 73108 195302 73160
rect 327718 73108 327724 73160
rect 327776 73148 327782 73160
rect 579614 73148 579620 73160
rect 327776 73120 579620 73148
rect 327776 73108 327782 73120
rect 579614 73108 579620 73120
rect 579672 73108 579678 73160
rect 121270 73040 121276 73092
rect 121328 73080 121334 73092
rect 129918 73080 129924 73092
rect 121328 73052 129924 73080
rect 121328 73040 121334 73052
rect 129918 73040 129924 73052
rect 129976 73080 129982 73092
rect 130746 73080 130752 73092
rect 129976 73052 130752 73080
rect 129976 73040 129982 73052
rect 130746 73040 130752 73052
rect 130804 73040 130810 73092
rect 131390 73040 131396 73092
rect 131448 73080 131454 73092
rect 132494 73080 132500 73092
rect 131448 73052 132500 73080
rect 131448 73040 131454 73052
rect 132494 73040 132500 73052
rect 132552 73040 132558 73092
rect 142338 73040 142344 73092
rect 142396 73080 142402 73092
rect 143442 73080 143448 73092
rect 142396 73052 143448 73080
rect 142396 73040 142402 73052
rect 143442 73040 143448 73052
rect 143500 73040 143506 73092
rect 159082 73040 159088 73092
rect 159140 73080 159146 73092
rect 194134 73080 194140 73092
rect 159140 73052 194140 73080
rect 159140 73040 159146 73052
rect 194134 73040 194140 73052
rect 194192 73040 194198 73092
rect 115658 72972 115664 73024
rect 115716 73012 115722 73024
rect 147858 73012 147864 73024
rect 115716 72984 147864 73012
rect 115716 72972 115722 72984
rect 147858 72972 147864 72984
rect 147916 73012 147922 73024
rect 148502 73012 148508 73024
rect 147916 72984 148508 73012
rect 147916 72972 147922 72984
rect 148502 72972 148508 72984
rect 148560 72972 148566 73024
rect 156690 72972 156696 73024
rect 156748 73012 156754 73024
rect 157150 73012 157156 73024
rect 156748 72984 157156 73012
rect 156748 72972 156754 72984
rect 157150 72972 157156 72984
rect 157208 73012 157214 73024
rect 210326 73012 210332 73024
rect 157208 72984 210332 73012
rect 157208 72972 157214 72984
rect 210326 72972 210332 72984
rect 210384 72972 210390 73024
rect 102594 72944 102600 72956
rect 84166 72916 102600 72944
rect 52454 72564 52460 72616
rect 52512 72604 52518 72616
rect 84166 72604 84194 72916
rect 102594 72904 102600 72916
rect 102652 72944 102658 72956
rect 136450 72944 136456 72956
rect 102652 72916 136456 72944
rect 102652 72904 102658 72916
rect 136450 72904 136456 72916
rect 136508 72904 136514 72956
rect 157242 72904 157248 72956
rect 157300 72944 157306 72956
rect 191006 72944 191012 72956
rect 157300 72916 191012 72944
rect 157300 72904 157306 72916
rect 191006 72904 191012 72916
rect 191064 72944 191070 72956
rect 191064 72916 200114 72944
rect 191064 72904 191070 72916
rect 107102 72836 107108 72888
rect 107160 72876 107166 72888
rect 140314 72876 140320 72888
rect 107160 72848 140320 72876
rect 107160 72836 107166 72848
rect 140314 72836 140320 72848
rect 140372 72836 140378 72888
rect 157702 72836 157708 72888
rect 157760 72876 157766 72888
rect 192478 72876 192484 72888
rect 157760 72848 192484 72876
rect 157760 72836 157766 72848
rect 192478 72836 192484 72848
rect 192536 72836 192542 72888
rect 110230 72768 110236 72820
rect 110288 72808 110294 72820
rect 142154 72808 142160 72820
rect 110288 72780 142160 72808
rect 110288 72768 110294 72780
rect 142154 72768 142160 72780
rect 142212 72768 142218 72820
rect 158254 72768 158260 72820
rect 158312 72808 158318 72820
rect 191834 72808 191840 72820
rect 158312 72780 191840 72808
rect 158312 72768 158318 72780
rect 191834 72768 191840 72780
rect 191892 72768 191898 72820
rect 117130 72700 117136 72752
rect 117188 72740 117194 72752
rect 148410 72740 148416 72752
rect 117188 72712 148416 72740
rect 117188 72700 117194 72712
rect 148410 72700 148416 72712
rect 148468 72740 148474 72752
rect 150894 72740 150900 72752
rect 148468 72712 150900 72740
rect 148468 72700 148474 72712
rect 150894 72700 150900 72712
rect 150952 72700 150958 72752
rect 154482 72700 154488 72752
rect 154540 72740 154546 72752
rect 187234 72740 187240 72752
rect 154540 72712 187240 72740
rect 154540 72700 154546 72712
rect 187234 72700 187240 72712
rect 187292 72700 187298 72752
rect 200086 72740 200114 72916
rect 218146 72836 218152 72888
rect 218204 72876 218210 72888
rect 218606 72876 218612 72888
rect 218204 72848 218612 72876
rect 218204 72836 218210 72848
rect 218606 72836 218612 72848
rect 218664 72876 218670 72888
rect 229738 72876 229744 72888
rect 218664 72848 229744 72876
rect 218664 72836 218670 72848
rect 229738 72836 229744 72848
rect 229796 72836 229802 72888
rect 216950 72768 216956 72820
rect 217008 72808 217014 72820
rect 342898 72808 342904 72820
rect 217008 72780 342904 72808
rect 217008 72768 217014 72780
rect 342898 72768 342904 72780
rect 342956 72768 342962 72820
rect 318794 72740 318800 72752
rect 200086 72712 318800 72740
rect 318794 72700 318800 72712
rect 318852 72700 318858 72752
rect 96614 72632 96620 72684
rect 96672 72672 96678 72684
rect 107102 72672 107108 72684
rect 96672 72644 107108 72672
rect 96672 72632 96678 72644
rect 107102 72632 107108 72644
rect 107160 72632 107166 72684
rect 111518 72632 111524 72684
rect 111576 72672 111582 72684
rect 142338 72672 142344 72684
rect 111576 72644 142344 72672
rect 111576 72632 111582 72644
rect 142338 72632 142344 72644
rect 142396 72632 142402 72684
rect 155862 72632 155868 72684
rect 155920 72672 155926 72684
rect 188338 72672 188344 72684
rect 155920 72644 188344 72672
rect 155920 72632 155926 72644
rect 188338 72632 188344 72644
rect 188396 72632 188402 72684
rect 192478 72632 192484 72684
rect 192536 72672 192542 72684
rect 323578 72672 323584 72684
rect 192536 72644 323584 72672
rect 192536 72632 192542 72644
rect 323578 72632 323584 72644
rect 323636 72632 323642 72684
rect 52512 72576 84194 72604
rect 52512 72564 52518 72576
rect 118510 72564 118516 72616
rect 118568 72604 118574 72616
rect 148134 72604 148140 72616
rect 118568 72576 148140 72604
rect 118568 72564 118574 72576
rect 148134 72564 148140 72576
rect 148192 72604 148198 72616
rect 148594 72604 148600 72616
rect 148192 72576 148600 72604
rect 148192 72564 148198 72576
rect 148594 72564 148600 72576
rect 148652 72564 148658 72616
rect 158346 72564 158352 72616
rect 158404 72604 158410 72616
rect 188154 72604 188160 72616
rect 158404 72576 188160 72604
rect 158404 72564 158410 72576
rect 188154 72564 188160 72576
rect 188212 72604 188218 72616
rect 332594 72604 332600 72616
rect 188212 72576 332600 72604
rect 188212 72564 188218 72576
rect 332594 72564 332600 72576
rect 332652 72564 332658 72616
rect 9674 72496 9680 72548
rect 9732 72536 9738 72548
rect 98822 72536 98828 72548
rect 9732 72508 98828 72536
rect 9732 72496 9738 72508
rect 98822 72496 98828 72508
rect 98880 72496 98886 72548
rect 99098 72496 99104 72548
rect 99156 72536 99162 72548
rect 131390 72536 131396 72548
rect 99156 72508 131396 72536
rect 99156 72496 99162 72508
rect 131390 72496 131396 72508
rect 131448 72496 131454 72548
rect 156414 72496 156420 72548
rect 156472 72536 156478 72548
rect 157150 72536 157156 72548
rect 156472 72508 157156 72536
rect 156472 72496 156478 72508
rect 157150 72496 157156 72508
rect 157208 72536 157214 72548
rect 190270 72536 190276 72548
rect 157208 72508 190276 72536
rect 157208 72496 157214 72508
rect 190270 72496 190276 72508
rect 190328 72496 190334 72548
rect 194134 72496 194140 72548
rect 194192 72536 194198 72548
rect 340966 72536 340972 72548
rect 194192 72508 340972 72536
rect 194192 72496 194198 72508
rect 340966 72496 340972 72508
rect 341024 72496 341030 72548
rect 4154 72428 4160 72480
rect 4212 72468 4218 72480
rect 99190 72468 99196 72480
rect 4212 72440 99196 72468
rect 4212 72428 4218 72440
rect 99190 72428 99196 72440
rect 99248 72428 99254 72480
rect 109678 72428 109684 72480
rect 109736 72468 109742 72480
rect 138198 72468 138204 72480
rect 109736 72440 138204 72468
rect 109736 72428 109742 72440
rect 138198 72428 138204 72440
rect 138256 72428 138262 72480
rect 146570 72428 146576 72480
rect 146628 72468 146634 72480
rect 182174 72468 182180 72480
rect 146628 72440 182180 72468
rect 146628 72428 146634 72440
rect 182174 72428 182180 72440
rect 182232 72428 182238 72480
rect 195238 72428 195244 72480
rect 195296 72468 195302 72480
rect 368474 72468 368480 72480
rect 195296 72440 368480 72468
rect 195296 72428 195302 72440
rect 368474 72428 368480 72440
rect 368532 72428 368538 72480
rect 109770 72360 109776 72412
rect 109828 72400 109834 72412
rect 121454 72400 121460 72412
rect 109828 72372 121460 72400
rect 109828 72360 109834 72372
rect 121454 72360 121460 72372
rect 121512 72400 121518 72412
rect 141510 72400 141516 72412
rect 121512 72372 141516 72400
rect 121512 72360 121518 72372
rect 141510 72360 141516 72372
rect 141568 72360 141574 72412
rect 161382 72360 161388 72412
rect 161440 72400 161446 72412
rect 194226 72400 194232 72412
rect 161440 72372 194232 72400
rect 161440 72360 161446 72372
rect 194226 72360 194232 72372
rect 194284 72360 194290 72412
rect 98822 72292 98828 72344
rect 98880 72332 98886 72344
rect 133138 72332 133144 72344
rect 98880 72304 133144 72332
rect 98880 72292 98886 72304
rect 133138 72292 133144 72304
rect 133196 72292 133202 72344
rect 159174 72292 159180 72344
rect 159232 72332 159238 72344
rect 216950 72332 216956 72344
rect 159232 72304 216956 72332
rect 159232 72292 159238 72304
rect 216950 72292 216956 72304
rect 217008 72292 217014 72344
rect 99190 72224 99196 72276
rect 99248 72264 99254 72276
rect 132586 72264 132592 72276
rect 99248 72236 132592 72264
rect 99248 72224 99254 72236
rect 132586 72224 132592 72236
rect 132644 72224 132650 72276
rect 155678 72224 155684 72276
rect 155736 72264 155742 72276
rect 218146 72264 218152 72276
rect 155736 72236 218152 72264
rect 155736 72224 155742 72236
rect 218146 72224 218152 72236
rect 218204 72224 218210 72276
rect 3510 71680 3516 71732
rect 3568 71720 3574 71732
rect 13078 71720 13084 71732
rect 3568 71692 13084 71720
rect 3568 71680 3574 71692
rect 13078 71680 13084 71692
rect 13136 71680 13142 71732
rect 121914 71680 121920 71732
rect 121972 71720 121978 71732
rect 149790 71720 149796 71732
rect 121972 71692 149796 71720
rect 121972 71680 121978 71692
rect 149790 71680 149796 71692
rect 149848 71680 149854 71732
rect 161106 71680 161112 71732
rect 161164 71720 161170 71732
rect 192294 71720 192300 71732
rect 161164 71692 192300 71720
rect 161164 71680 161170 71692
rect 192294 71680 192300 71692
rect 192352 71680 192358 71732
rect 105814 71612 105820 71664
rect 105872 71652 105878 71664
rect 140038 71652 140044 71664
rect 105872 71624 140044 71652
rect 105872 71612 105878 71624
rect 140038 71612 140044 71624
rect 140096 71612 140102 71664
rect 157518 71612 157524 71664
rect 157576 71652 157582 71664
rect 158254 71652 158260 71664
rect 157576 71624 158260 71652
rect 157576 71612 157582 71624
rect 158254 71612 158260 71624
rect 158312 71612 158318 71664
rect 159910 71612 159916 71664
rect 159968 71652 159974 71664
rect 193766 71652 193772 71664
rect 159968 71624 193772 71652
rect 159968 71612 159974 71624
rect 193766 71612 193772 71624
rect 193824 71612 193830 71664
rect 104526 71544 104532 71596
rect 104584 71584 104590 71596
rect 137922 71584 137928 71596
rect 104584 71556 137928 71584
rect 104584 71544 104590 71556
rect 137922 71544 137928 71556
rect 137980 71544 137986 71596
rect 158272 71584 158300 71612
rect 192386 71584 192392 71596
rect 158272 71556 192392 71584
rect 192386 71544 192392 71556
rect 192444 71544 192450 71596
rect 118142 71476 118148 71528
rect 118200 71516 118206 71528
rect 147950 71516 147956 71528
rect 118200 71488 147956 71516
rect 118200 71476 118206 71488
rect 147950 71476 147956 71488
rect 148008 71516 148014 71528
rect 150158 71516 150164 71528
rect 148008 71488 150164 71516
rect 148008 71476 148014 71488
rect 150158 71476 150164 71488
rect 150216 71476 150222 71528
rect 157334 71476 157340 71528
rect 157392 71516 157398 71528
rect 158438 71516 158444 71528
rect 157392 71488 158444 71516
rect 157392 71476 157398 71488
rect 158438 71476 158444 71488
rect 158496 71476 158502 71528
rect 160738 71476 160744 71528
rect 160796 71516 160802 71528
rect 195054 71516 195060 71528
rect 160796 71488 195060 71516
rect 160796 71476 160802 71488
rect 195054 71476 195060 71488
rect 195112 71476 195118 71528
rect 116854 71408 116860 71460
rect 116912 71448 116918 71460
rect 148226 71448 148232 71460
rect 116912 71420 148232 71448
rect 116912 71408 116918 71420
rect 148226 71408 148232 71420
rect 148284 71448 148290 71460
rect 148502 71448 148508 71460
rect 148284 71420 148508 71448
rect 148284 71408 148290 71420
rect 148502 71408 148508 71420
rect 148560 71408 148566 71460
rect 159818 71408 159824 71460
rect 159876 71448 159882 71460
rect 193674 71448 193680 71460
rect 159876 71420 193680 71448
rect 159876 71408 159882 71420
rect 193674 71408 193680 71420
rect 193732 71408 193738 71460
rect 134978 71380 134984 71392
rect 109006 71352 134984 71380
rect 109006 71312 109034 71352
rect 134978 71340 134984 71352
rect 135036 71340 135042 71392
rect 157334 71340 157340 71392
rect 157392 71380 157398 71392
rect 157794 71380 157800 71392
rect 157392 71352 157800 71380
rect 157392 71340 157398 71352
rect 157794 71340 157800 71352
rect 157852 71340 157858 71392
rect 158438 71340 158444 71392
rect 158496 71380 158502 71392
rect 161106 71380 161112 71392
rect 158496 71352 161112 71380
rect 158496 71340 158502 71352
rect 161106 71340 161112 71352
rect 161164 71340 161170 71392
rect 162762 71340 162768 71392
rect 162820 71380 162826 71392
rect 196526 71380 196532 71392
rect 162820 71352 196532 71380
rect 162820 71340 162826 71352
rect 196526 71340 196532 71352
rect 196584 71340 196590 71392
rect 108316 71284 109034 71312
rect 71774 71136 71780 71188
rect 71832 71176 71838 71188
rect 104526 71176 104532 71188
rect 71832 71148 104532 71176
rect 71832 71136 71838 71148
rect 104526 71136 104532 71148
rect 104584 71136 104590 71188
rect 35158 71068 35164 71120
rect 35216 71108 35222 71120
rect 103238 71108 103244 71120
rect 35216 71080 103244 71108
rect 35216 71068 35222 71080
rect 103238 71068 103244 71080
rect 103296 71108 103302 71120
rect 108316 71108 108344 71284
rect 119614 71272 119620 71324
rect 119672 71312 119678 71324
rect 150066 71312 150072 71324
rect 119672 71284 150072 71312
rect 119672 71272 119678 71284
rect 150066 71272 150072 71284
rect 150124 71272 150130 71324
rect 166258 71272 166264 71324
rect 166316 71312 166322 71324
rect 166902 71312 166908 71324
rect 166316 71284 166908 71312
rect 166316 71272 166322 71284
rect 166902 71272 166908 71284
rect 166960 71312 166966 71324
rect 200666 71312 200672 71324
rect 166960 71284 200672 71312
rect 166960 71272 166966 71284
rect 200666 71272 200672 71284
rect 200724 71272 200730 71324
rect 112070 71204 112076 71256
rect 112128 71244 112134 71256
rect 142798 71244 142804 71256
rect 112128 71216 142804 71244
rect 112128 71204 112134 71216
rect 142798 71204 142804 71216
rect 142856 71204 142862 71256
rect 160922 71204 160928 71256
rect 160980 71244 160986 71256
rect 195514 71244 195520 71256
rect 160980 71216 195520 71244
rect 160980 71204 160986 71216
rect 195514 71204 195520 71216
rect 195572 71204 195578 71256
rect 122098 71136 122104 71188
rect 122156 71176 122162 71188
rect 151446 71176 151452 71188
rect 122156 71148 151452 71176
rect 122156 71136 122162 71148
rect 151446 71136 151452 71148
rect 151504 71136 151510 71188
rect 153562 71136 153568 71188
rect 153620 71176 153626 71188
rect 187050 71176 187056 71188
rect 153620 71148 187056 71176
rect 153620 71136 153626 71148
rect 187050 71136 187056 71148
rect 187108 71136 187114 71188
rect 133414 71108 133420 71120
rect 103296 71080 108344 71108
rect 108408 71080 133420 71108
rect 103296 71068 103302 71080
rect 27614 71000 27620 71052
rect 27672 71040 27678 71052
rect 99926 71040 99932 71052
rect 27672 71012 99932 71040
rect 27672 71000 27678 71012
rect 99926 71000 99932 71012
rect 99984 71040 99990 71052
rect 99984 71012 103514 71040
rect 99984 71000 99990 71012
rect 103486 70972 103514 71012
rect 107378 71000 107384 71052
rect 107436 71040 107442 71052
rect 108408 71040 108436 71080
rect 133414 71068 133420 71080
rect 133472 71068 133478 71120
rect 147122 71068 147128 71120
rect 147180 71108 147186 71120
rect 184198 71108 184204 71120
rect 147180 71080 184204 71108
rect 147180 71068 147186 71080
rect 184198 71068 184204 71080
rect 184256 71068 184262 71120
rect 107436 71012 108436 71040
rect 107436 71000 107442 71012
rect 111702 71000 111708 71052
rect 111760 71040 111766 71052
rect 128354 71040 128360 71052
rect 111760 71012 128360 71040
rect 111760 71000 111766 71012
rect 128354 71000 128360 71012
rect 128412 71040 128418 71052
rect 129550 71040 129556 71052
rect 128412 71012 129556 71040
rect 128412 71000 128418 71012
rect 129550 71000 129556 71012
rect 129608 71000 129614 71052
rect 150894 71000 150900 71052
rect 150952 71040 150958 71052
rect 200114 71040 200120 71052
rect 150952 71012 200120 71040
rect 150952 71000 150958 71012
rect 200114 71000 200120 71012
rect 200172 71000 200178 71052
rect 134426 70972 134432 70984
rect 103486 70944 134432 70972
rect 134426 70932 134432 70944
rect 134484 70932 134490 70984
rect 160002 70932 160008 70984
rect 160060 70972 160066 70984
rect 192846 70972 192852 70984
rect 160060 70944 192852 70972
rect 160060 70932 160066 70944
rect 192846 70932 192852 70944
rect 192904 70932 192910 70984
rect 157058 70864 157064 70916
rect 157116 70904 157122 70916
rect 188614 70904 188620 70916
rect 157116 70876 188620 70904
rect 157116 70864 157122 70876
rect 188614 70864 188620 70876
rect 188672 70864 188678 70916
rect 158530 70796 158536 70848
rect 158588 70836 158594 70848
rect 188062 70836 188068 70848
rect 158588 70808 188068 70836
rect 158588 70796 158594 70808
rect 188062 70796 188068 70808
rect 188120 70796 188126 70848
rect 169202 70728 169208 70780
rect 169260 70768 169266 70780
rect 169386 70768 169392 70780
rect 169260 70740 169392 70768
rect 169260 70728 169266 70740
rect 169386 70728 169392 70740
rect 169444 70728 169450 70780
rect 149790 70592 149796 70644
rect 149848 70632 149854 70644
rect 150250 70632 150256 70644
rect 149848 70604 150256 70632
rect 149848 70592 149854 70604
rect 150250 70592 150256 70604
rect 150308 70592 150314 70644
rect 103514 70388 103520 70440
rect 103572 70428 103578 70440
rect 105814 70428 105820 70440
rect 103572 70400 105820 70428
rect 103572 70388 103578 70400
rect 105814 70388 105820 70400
rect 105872 70388 105878 70440
rect 113174 70388 113180 70440
rect 113232 70428 113238 70440
rect 115106 70428 115112 70440
rect 113232 70400 115112 70428
rect 113232 70388 113238 70400
rect 115106 70388 115112 70400
rect 115164 70388 115170 70440
rect 100754 70320 100760 70372
rect 100812 70360 100818 70372
rect 101306 70360 101312 70372
rect 100812 70332 101312 70360
rect 100812 70320 100818 70332
rect 101306 70320 101312 70332
rect 101364 70360 101370 70372
rect 135990 70360 135996 70372
rect 101364 70332 135996 70360
rect 101364 70320 101370 70332
rect 135990 70320 135996 70332
rect 136048 70320 136054 70372
rect 168006 70320 168012 70372
rect 168064 70360 168070 70372
rect 214282 70360 214288 70372
rect 168064 70332 214288 70360
rect 168064 70320 168070 70332
rect 214282 70320 214288 70332
rect 214340 70320 214346 70372
rect 118878 70252 118884 70304
rect 118936 70292 118942 70304
rect 152090 70292 152096 70304
rect 118936 70264 152096 70292
rect 118936 70252 118942 70264
rect 152090 70252 152096 70264
rect 152148 70292 152154 70304
rect 152642 70292 152648 70304
rect 152148 70264 152648 70292
rect 152148 70252 152154 70264
rect 152642 70252 152648 70264
rect 152700 70252 152706 70304
rect 164050 70252 164056 70304
rect 164108 70292 164114 70304
rect 204990 70292 204996 70304
rect 164108 70264 204996 70292
rect 164108 70252 164114 70264
rect 204990 70252 204996 70264
rect 205048 70252 205054 70304
rect 104158 70184 104164 70236
rect 104216 70224 104222 70236
rect 137186 70224 137192 70236
rect 104216 70196 137192 70224
rect 104216 70184 104222 70196
rect 137186 70184 137192 70196
rect 137244 70184 137250 70236
rect 161842 70184 161848 70236
rect 161900 70224 161906 70236
rect 196618 70224 196624 70236
rect 161900 70196 196624 70224
rect 161900 70184 161906 70196
rect 196618 70184 196624 70196
rect 196676 70184 196682 70236
rect 105998 70156 106004 70168
rect 103486 70128 106004 70156
rect 85666 69776 85672 69828
rect 85724 69816 85730 69828
rect 103486 69816 103514 70128
rect 105998 70116 106004 70128
rect 106056 70156 106062 70168
rect 139026 70156 139032 70168
rect 106056 70128 139032 70156
rect 106056 70116 106062 70128
rect 139026 70116 139032 70128
rect 139084 70116 139090 70168
rect 162302 70116 162308 70168
rect 162360 70156 162366 70168
rect 196710 70156 196716 70168
rect 162360 70128 196716 70156
rect 162360 70116 162366 70128
rect 196710 70116 196716 70128
rect 196768 70116 196774 70168
rect 108390 70048 108396 70100
rect 108448 70088 108454 70100
rect 108666 70088 108672 70100
rect 108448 70060 108672 70088
rect 108448 70048 108454 70060
rect 108666 70048 108672 70060
rect 108724 70088 108730 70100
rect 139946 70088 139952 70100
rect 108724 70060 139952 70088
rect 108724 70048 108730 70060
rect 139946 70048 139952 70060
rect 140004 70048 140010 70100
rect 160462 70048 160468 70100
rect 160520 70088 160526 70100
rect 161198 70088 161204 70100
rect 160520 70060 161204 70088
rect 160520 70048 160526 70060
rect 161198 70048 161204 70060
rect 161256 70088 161262 70100
rect 194962 70088 194968 70100
rect 161256 70060 194968 70088
rect 161256 70048 161262 70060
rect 194962 70048 194968 70060
rect 195020 70048 195026 70100
rect 120810 69980 120816 70032
rect 120868 70020 120874 70032
rect 150986 70020 150992 70032
rect 120868 69992 150992 70020
rect 120868 69980 120874 69992
rect 150986 69980 150992 69992
rect 151044 69980 151050 70032
rect 163958 69980 163964 70032
rect 164016 70020 164022 70032
rect 197906 70020 197912 70032
rect 164016 69992 197912 70020
rect 164016 69980 164022 69992
rect 197906 69980 197912 69992
rect 197964 69980 197970 70032
rect 111978 69912 111984 69964
rect 112036 69952 112042 69964
rect 142430 69952 142436 69964
rect 112036 69924 142436 69952
rect 112036 69912 112042 69924
rect 142430 69912 142436 69924
rect 142488 69912 142494 69964
rect 163314 69912 163320 69964
rect 163372 69952 163378 69964
rect 164050 69952 164056 69964
rect 163372 69924 164056 69952
rect 163372 69912 163378 69924
rect 164050 69912 164056 69924
rect 164108 69912 164114 69964
rect 165154 69912 165160 69964
rect 165212 69952 165218 69964
rect 199286 69952 199292 69964
rect 165212 69924 199292 69952
rect 165212 69912 165218 69924
rect 199286 69912 199292 69924
rect 199344 69912 199350 69964
rect 113542 69844 113548 69896
rect 113600 69884 113606 69896
rect 142982 69884 142988 69896
rect 113600 69856 142988 69884
rect 113600 69844 113606 69856
rect 142982 69844 142988 69856
rect 143040 69844 143046 69896
rect 151354 69844 151360 69896
rect 151412 69884 151418 69896
rect 242158 69884 242164 69896
rect 151412 69856 242164 69884
rect 151412 69844 151418 69856
rect 242158 69844 242164 69856
rect 242216 69844 242222 69896
rect 85724 69788 103514 69816
rect 85724 69776 85730 69788
rect 115106 69776 115112 69828
rect 115164 69816 115170 69828
rect 141326 69816 141332 69828
rect 115164 69788 141332 69816
rect 115164 69776 115170 69788
rect 141326 69776 141332 69788
rect 141384 69776 141390 69828
rect 150986 69776 150992 69828
rect 151044 69816 151050 69828
rect 151538 69816 151544 69828
rect 151044 69788 151544 69816
rect 151044 69776 151050 69788
rect 151538 69776 151544 69788
rect 151596 69776 151602 69828
rect 160370 69776 160376 69828
rect 160428 69816 160434 69828
rect 194686 69816 194692 69828
rect 160428 69788 194692 69816
rect 160428 69776 160434 69788
rect 194686 69776 194692 69788
rect 194744 69816 194750 69828
rect 362954 69816 362960 69828
rect 194744 69788 362960 69816
rect 194744 69776 194750 69788
rect 362954 69776 362960 69788
rect 363012 69776 363018 69828
rect 60826 69708 60832 69760
rect 60884 69748 60890 69760
rect 104158 69748 104164 69760
rect 60884 69720 104164 69748
rect 60884 69708 60890 69720
rect 104158 69708 104164 69720
rect 104216 69708 104222 69760
rect 117314 69708 117320 69760
rect 117372 69748 117378 69760
rect 117774 69748 117780 69760
rect 117372 69720 117780 69748
rect 117372 69708 117378 69720
rect 117774 69708 117780 69720
rect 117832 69748 117838 69760
rect 141050 69748 141056 69760
rect 117832 69720 141056 69748
rect 117832 69708 117838 69720
rect 141050 69708 141056 69720
rect 141108 69708 141114 69760
rect 163406 69708 163412 69760
rect 163464 69748 163470 69760
rect 163958 69748 163964 69760
rect 163464 69720 163964 69748
rect 163464 69708 163470 69720
rect 163958 69708 163964 69720
rect 164016 69708 164022 69760
rect 164786 69708 164792 69760
rect 164844 69748 164850 69760
rect 165154 69748 165160 69760
rect 164844 69720 165160 69748
rect 164844 69708 164850 69720
rect 165154 69708 165160 69720
rect 165212 69708 165218 69760
rect 166166 69708 166172 69760
rect 166224 69748 166230 69760
rect 166224 69720 200114 69748
rect 166224 69708 166230 69720
rect 45554 69640 45560 69692
rect 45612 69680 45618 69692
rect 100754 69680 100760 69692
rect 45612 69652 100760 69680
rect 45612 69640 45618 69652
rect 100754 69640 100760 69652
rect 100812 69640 100818 69692
rect 102870 69640 102876 69692
rect 102928 69680 102934 69692
rect 108390 69680 108396 69692
rect 102928 69652 108396 69680
rect 102928 69640 102934 69652
rect 108390 69640 108396 69652
rect 108448 69640 108454 69692
rect 148594 69640 148600 69692
rect 148652 69680 148658 69692
rect 189718 69680 189724 69692
rect 148652 69652 189724 69680
rect 148652 69640 148658 69652
rect 189718 69640 189724 69652
rect 189776 69640 189782 69692
rect 200086 69680 200114 69720
rect 214282 69708 214288 69760
rect 214340 69748 214346 69760
rect 397454 69748 397460 69760
rect 214340 69720 397460 69748
rect 214340 69708 214346 69720
rect 397454 69708 397460 69720
rect 397512 69708 397518 69760
rect 201126 69680 201132 69692
rect 200086 69652 201132 69680
rect 201126 69640 201132 69652
rect 201184 69680 201190 69692
rect 430574 69680 430580 69692
rect 201184 69652 430580 69680
rect 201184 69640 201190 69652
rect 430574 69640 430580 69652
rect 430632 69640 430638 69692
rect 161934 69572 161940 69624
rect 161992 69612 161998 69624
rect 162670 69612 162676 69624
rect 161992 69584 162676 69612
rect 161992 69572 161998 69584
rect 162670 69572 162676 69584
rect 162728 69572 162734 69624
rect 166074 69572 166080 69624
rect 166132 69612 166138 69624
rect 166718 69612 166724 69624
rect 166132 69584 166724 69612
rect 166132 69572 166138 69584
rect 166718 69572 166724 69584
rect 166776 69572 166782 69624
rect 194778 69612 194784 69624
rect 171106 69584 194784 69612
rect 162688 69544 162716 69572
rect 171106 69544 171134 69584
rect 194778 69572 194784 69584
rect 194836 69572 194842 69624
rect 162688 69516 171134 69544
rect 178862 69504 178868 69556
rect 178920 69544 178926 69556
rect 210326 69544 210332 69556
rect 178920 69516 210332 69544
rect 178920 69504 178926 69516
rect 210326 69504 210332 69516
rect 210384 69544 210390 69556
rect 210694 69544 210700 69556
rect 210384 69516 210700 69544
rect 210384 69504 210390 69516
rect 210694 69504 210700 69516
rect 210752 69504 210758 69556
rect 166718 69436 166724 69488
rect 166776 69476 166782 69488
rect 186866 69476 186872 69488
rect 166776 69448 186872 69476
rect 166776 69436 166782 69448
rect 186866 69436 186872 69448
rect 186924 69436 186930 69488
rect 140038 69028 140044 69080
rect 140096 69068 140102 69080
rect 142154 69068 142160 69080
rect 140096 69040 142160 69068
rect 140096 69028 140102 69040
rect 142154 69028 142160 69040
rect 142212 69028 142218 69080
rect 110046 68960 110052 69012
rect 110104 69000 110110 69012
rect 143902 69000 143908 69012
rect 110104 68972 143908 69000
rect 110104 68960 110110 68972
rect 143902 68960 143908 68972
rect 143960 68960 143966 69012
rect 155034 68960 155040 69012
rect 155092 69000 155098 69012
rect 155862 69000 155868 69012
rect 155092 68972 155868 69000
rect 155092 68960 155098 68972
rect 155862 68960 155868 68972
rect 155920 69000 155926 69012
rect 197814 69000 197820 69012
rect 155920 68972 197820 69000
rect 155920 68960 155926 68972
rect 197814 68960 197820 68972
rect 197872 68960 197878 69012
rect 100754 68892 100760 68944
rect 100812 68932 100818 68944
rect 101582 68932 101588 68944
rect 100812 68904 101588 68932
rect 100812 68892 100818 68904
rect 101582 68892 101588 68904
rect 101640 68932 101646 68944
rect 135622 68932 135628 68944
rect 101640 68904 135628 68932
rect 101640 68892 101646 68904
rect 135622 68892 135628 68904
rect 135680 68892 135686 68944
rect 163222 68892 163228 68944
rect 163280 68932 163286 68944
rect 163866 68932 163872 68944
rect 163280 68904 163872 68932
rect 163280 68892 163286 68904
rect 163866 68892 163872 68904
rect 163924 68892 163930 68944
rect 164694 68892 164700 68944
rect 164752 68932 164758 68944
rect 165430 68932 165436 68944
rect 164752 68904 165436 68932
rect 164752 68892 164758 68904
rect 165430 68892 165436 68904
rect 165488 68892 165494 68944
rect 165982 68892 165988 68944
rect 166040 68932 166046 68944
rect 166810 68932 166816 68944
rect 166040 68904 166816 68932
rect 166040 68892 166046 68904
rect 166810 68892 166816 68904
rect 166868 68892 166874 68944
rect 167362 68892 167368 68944
rect 167420 68932 167426 68944
rect 168190 68932 168196 68944
rect 167420 68904 168196 68932
rect 167420 68892 167426 68904
rect 168190 68892 168196 68904
rect 168248 68932 168254 68944
rect 202230 68932 202236 68944
rect 168248 68904 202236 68932
rect 168248 68892 168254 68904
rect 202230 68892 202236 68904
rect 202288 68892 202294 68944
rect 108758 68824 108764 68876
rect 108816 68864 108822 68876
rect 142154 68864 142160 68876
rect 108816 68836 142160 68864
rect 108816 68824 108822 68836
rect 142154 68824 142160 68836
rect 142212 68864 142218 68876
rect 142706 68864 142712 68876
rect 142212 68836 142712 68864
rect 142212 68824 142218 68836
rect 142706 68824 142712 68836
rect 142764 68824 142770 68876
rect 167454 68824 167460 68876
rect 167512 68864 167518 68876
rect 168098 68864 168104 68876
rect 167512 68836 168104 68864
rect 167512 68824 167518 68836
rect 168098 68824 168104 68836
rect 168156 68864 168162 68876
rect 202138 68864 202144 68876
rect 168156 68836 202144 68864
rect 168156 68824 168162 68836
rect 202138 68824 202144 68836
rect 202196 68824 202202 68876
rect 108942 68756 108948 68808
rect 109000 68796 109006 68808
rect 142890 68796 142896 68808
rect 109000 68768 142896 68796
rect 109000 68756 109006 68768
rect 142890 68756 142896 68768
rect 142948 68756 142954 68808
rect 166810 68756 166816 68808
rect 166868 68796 166874 68808
rect 200574 68796 200580 68808
rect 166868 68768 200580 68796
rect 166868 68756 166874 68768
rect 200574 68756 200580 68768
rect 200632 68756 200638 68808
rect 112530 68688 112536 68740
rect 112588 68728 112594 68740
rect 144086 68728 144092 68740
rect 112588 68700 144092 68728
rect 112588 68688 112594 68700
rect 144086 68688 144092 68700
rect 144144 68688 144150 68740
rect 168742 68688 168748 68740
rect 168800 68728 168806 68740
rect 169386 68728 169392 68740
rect 168800 68700 169392 68728
rect 168800 68688 168806 68700
rect 169386 68688 169392 68700
rect 169444 68728 169450 68740
rect 203334 68728 203340 68740
rect 169444 68700 203340 68728
rect 169444 68688 169450 68700
rect 203334 68688 203340 68700
rect 203392 68688 203398 68740
rect 106826 68620 106832 68672
rect 106884 68660 106890 68672
rect 138014 68660 138020 68672
rect 106884 68632 138020 68660
rect 106884 68620 106890 68632
rect 138014 68620 138020 68632
rect 138072 68660 138078 68672
rect 138566 68660 138572 68672
rect 138072 68632 138572 68660
rect 138072 68620 138078 68632
rect 138566 68620 138572 68632
rect 138624 68620 138630 68672
rect 175918 68620 175924 68672
rect 175976 68660 175982 68672
rect 199838 68660 199844 68672
rect 175976 68632 199844 68660
rect 175976 68620 175982 68632
rect 199838 68620 199844 68632
rect 199896 68620 199902 68672
rect 102134 68552 102140 68604
rect 102192 68592 102198 68604
rect 103054 68592 103060 68604
rect 102192 68564 103060 68592
rect 102192 68552 102198 68564
rect 103054 68552 103060 68564
rect 103112 68592 103118 68604
rect 134242 68592 134248 68604
rect 103112 68564 134248 68592
rect 103112 68552 103118 68564
rect 134242 68552 134248 68564
rect 134300 68552 134306 68604
rect 163866 68552 163872 68604
rect 163924 68592 163930 68604
rect 198274 68592 198280 68604
rect 163924 68564 198280 68592
rect 163924 68552 163930 68564
rect 198274 68552 198280 68564
rect 198332 68552 198338 68604
rect 114002 68484 114008 68536
rect 114060 68524 114066 68536
rect 143994 68524 144000 68536
rect 114060 68496 144000 68524
rect 114060 68484 114066 68496
rect 143994 68484 144000 68496
rect 144052 68484 144058 68536
rect 160186 68484 160192 68536
rect 160244 68524 160250 68536
rect 194594 68524 194600 68536
rect 160244 68496 194600 68524
rect 160244 68484 160250 68496
rect 194594 68484 194600 68496
rect 194652 68524 194658 68536
rect 195054 68524 195060 68536
rect 194652 68496 195060 68524
rect 194652 68484 194658 68496
rect 195054 68484 195060 68496
rect 195112 68484 195118 68536
rect 102226 68416 102232 68468
rect 102284 68456 102290 68468
rect 132770 68456 132776 68468
rect 102284 68428 132776 68456
rect 102284 68416 102290 68428
rect 132770 68416 132776 68428
rect 132828 68416 132834 68468
rect 165430 68416 165436 68468
rect 165488 68456 165494 68468
rect 175918 68456 175924 68468
rect 165488 68428 175924 68456
rect 165488 68416 165494 68428
rect 175918 68416 175924 68428
rect 175976 68416 175982 68468
rect 176562 68416 176568 68468
rect 176620 68456 176626 68468
rect 210418 68456 210424 68468
rect 176620 68428 210424 68456
rect 176620 68416 176626 68428
rect 210418 68416 210424 68428
rect 210476 68416 210482 68468
rect 116210 68348 116216 68400
rect 116268 68388 116274 68400
rect 141418 68388 141424 68400
rect 116268 68360 141424 68388
rect 116268 68348 116274 68360
rect 141418 68348 141424 68360
rect 141476 68348 141482 68400
rect 164602 68348 164608 68400
rect 164660 68388 164666 68400
rect 189074 68388 189080 68400
rect 164660 68360 189080 68388
rect 164660 68348 164666 68360
rect 189074 68348 189080 68360
rect 189132 68348 189138 68400
rect 48314 68280 48320 68332
rect 48372 68320 48378 68332
rect 100754 68320 100760 68332
rect 48372 68292 100760 68320
rect 48372 68280 48378 68292
rect 100754 68280 100760 68292
rect 100812 68280 100818 68332
rect 110782 68280 110788 68332
rect 110840 68320 110846 68332
rect 120166 68320 120172 68332
rect 110840 68292 120172 68320
rect 110840 68280 110846 68292
rect 120166 68280 120172 68292
rect 120224 68320 120230 68332
rect 141234 68320 141240 68332
rect 120224 68292 141240 68320
rect 120224 68280 120230 68292
rect 141234 68280 141240 68292
rect 141292 68280 141298 68332
rect 160278 68280 160284 68332
rect 160336 68320 160342 68332
rect 161106 68320 161112 68332
rect 160336 68292 161112 68320
rect 160336 68280 160342 68292
rect 161106 68280 161112 68292
rect 161164 68320 161170 68332
rect 184382 68320 184388 68332
rect 161164 68292 184388 68320
rect 161164 68280 161170 68292
rect 184382 68280 184388 68292
rect 184440 68280 184446 68332
rect 195054 68280 195060 68332
rect 195112 68320 195118 68332
rect 358814 68320 358820 68332
rect 195112 68292 358820 68320
rect 195112 68280 195118 68292
rect 358814 68280 358820 68292
rect 358872 68280 358878 68332
rect 175826 68212 175832 68264
rect 175884 68252 175890 68264
rect 176562 68252 176568 68264
rect 175884 68224 176568 68252
rect 175884 68212 175890 68224
rect 176562 68212 176568 68224
rect 176620 68212 176626 68264
rect 177574 68212 177580 68264
rect 177632 68252 177638 68264
rect 200758 68252 200764 68264
rect 177632 68224 200764 68252
rect 177632 68212 177638 68224
rect 200758 68212 200764 68224
rect 200816 68252 200822 68264
rect 201402 68252 201408 68264
rect 200816 68224 201408 68252
rect 200816 68212 200822 68224
rect 201402 68212 201408 68224
rect 201460 68212 201466 68264
rect 189074 67736 189080 67788
rect 189132 67776 189138 67788
rect 422938 67776 422944 67788
rect 189132 67748 422944 67776
rect 189132 67736 189138 67748
rect 422938 67736 422944 67748
rect 422996 67736 423002 67788
rect 188430 67668 188436 67720
rect 188488 67708 188494 67720
rect 507854 67708 507860 67720
rect 188488 67680 507860 67708
rect 188488 67668 188494 67680
rect 507854 67668 507860 67680
rect 507912 67668 507918 67720
rect 141418 67600 141424 67652
rect 141476 67640 141482 67652
rect 142246 67640 142252 67652
rect 141476 67612 142252 67640
rect 141476 67600 141482 67612
rect 142246 67600 142252 67612
rect 142304 67600 142310 67652
rect 144086 67600 144092 67652
rect 144144 67640 144150 67652
rect 144362 67640 144368 67652
rect 144144 67612 144368 67640
rect 144144 67600 144150 67612
rect 144362 67600 144368 67612
rect 144420 67600 144426 67652
rect 201402 67600 201408 67652
rect 201460 67640 201466 67652
rect 536834 67640 536840 67652
rect 201460 67612 536840 67640
rect 201460 67600 201466 67612
rect 536834 67600 536840 67612
rect 536892 67600 536898 67652
rect 99282 67532 99288 67584
rect 99340 67572 99346 67584
rect 132678 67572 132684 67584
rect 99340 67544 132684 67572
rect 99340 67532 99346 67544
rect 132678 67532 132684 67544
rect 132736 67572 132742 67584
rect 133230 67572 133236 67584
rect 132736 67544 133236 67572
rect 132736 67532 132742 67544
rect 133230 67532 133236 67544
rect 133288 67532 133294 67584
rect 150618 67532 150624 67584
rect 150676 67572 150682 67584
rect 151078 67572 151084 67584
rect 150676 67544 151084 67572
rect 150676 67532 150682 67544
rect 151078 67532 151084 67544
rect 151136 67532 151142 67584
rect 172606 67532 172612 67584
rect 172664 67572 172670 67584
rect 212902 67572 212908 67584
rect 172664 67544 212908 67572
rect 172664 67532 172670 67544
rect 212902 67532 212908 67544
rect 212960 67572 212966 67584
rect 213822 67572 213828 67584
rect 212960 67544 213828 67572
rect 212960 67532 212966 67544
rect 213822 67532 213828 67544
rect 213880 67532 213886 67584
rect 108850 67464 108856 67516
rect 108908 67504 108914 67516
rect 135254 67504 135260 67516
rect 108908 67476 135260 67504
rect 108908 67464 108914 67476
rect 135254 67464 135260 67476
rect 135312 67504 135318 67516
rect 142614 67504 142620 67516
rect 135312 67476 142620 67504
rect 135312 67464 135318 67476
rect 142614 67464 142620 67476
rect 142672 67464 142678 67516
rect 172790 67464 172796 67516
rect 172848 67504 172854 67516
rect 173618 67504 173624 67516
rect 172848 67476 173624 67504
rect 172848 67464 172854 67476
rect 173618 67464 173624 67476
rect 173676 67464 173682 67516
rect 174262 67464 174268 67516
rect 174320 67504 174326 67516
rect 174722 67504 174728 67516
rect 174320 67476 174728 67504
rect 174320 67464 174326 67476
rect 174722 67464 174728 67476
rect 174780 67464 174786 67516
rect 175642 67464 175648 67516
rect 175700 67504 175706 67516
rect 215570 67504 215576 67516
rect 175700 67476 215576 67504
rect 175700 67464 175706 67476
rect 215570 67464 215576 67476
rect 215628 67464 215634 67516
rect 120350 67396 120356 67448
rect 120408 67436 120414 67448
rect 151906 67436 151912 67448
rect 120408 67408 151912 67436
rect 120408 67396 120414 67408
rect 151906 67396 151912 67408
rect 151964 67436 151970 67448
rect 152550 67436 152556 67448
rect 151964 67408 152556 67436
rect 151964 67396 151970 67408
rect 152550 67396 152556 67408
rect 152608 67396 152614 67448
rect 172698 67396 172704 67448
rect 172756 67436 172762 67448
rect 173434 67436 173440 67448
rect 172756 67408 173440 67436
rect 172756 67396 172762 67408
rect 173434 67396 173440 67408
rect 173492 67396 173498 67448
rect 174170 67396 174176 67448
rect 174228 67436 174234 67448
rect 174998 67436 175004 67448
rect 174228 67408 175004 67436
rect 174228 67396 174234 67408
rect 174998 67396 175004 67408
rect 175056 67396 175062 67448
rect 175734 67396 175740 67448
rect 175792 67436 175798 67448
rect 176286 67436 176292 67448
rect 175792 67408 176292 67436
rect 175792 67396 175798 67408
rect 176286 67396 176292 67408
rect 176344 67396 176350 67448
rect 208946 67436 208952 67448
rect 176672 67408 208952 67436
rect 117590 67328 117596 67380
rect 117648 67368 117654 67380
rect 149146 67368 149152 67380
rect 117648 67340 149152 67368
rect 117648 67328 117654 67340
rect 149146 67328 149152 67340
rect 149204 67328 149210 67380
rect 174078 67328 174084 67380
rect 174136 67368 174142 67380
rect 174814 67368 174820 67380
rect 174136 67340 174820 67368
rect 174136 67328 174142 67340
rect 174814 67328 174820 67340
rect 174872 67328 174878 67380
rect 175550 67328 175556 67380
rect 175608 67368 175614 67380
rect 176470 67368 176476 67380
rect 175608 67340 176476 67368
rect 175608 67328 175614 67340
rect 176470 67328 176476 67340
rect 176528 67328 176534 67380
rect 104526 67260 104532 67312
rect 104584 67300 104590 67312
rect 136082 67300 136088 67312
rect 104584 67272 136088 67300
rect 104584 67260 104590 67272
rect 136082 67260 136088 67272
rect 136140 67260 136146 67312
rect 174998 67260 175004 67312
rect 175056 67300 175062 67312
rect 176672 67300 176700 67408
rect 208946 67396 208952 67408
rect 209004 67396 209010 67448
rect 177206 67328 177212 67380
rect 177264 67368 177270 67380
rect 207474 67368 207480 67380
rect 177264 67340 207480 67368
rect 177264 67328 177270 67340
rect 207474 67328 207480 67340
rect 207532 67328 207538 67380
rect 208762 67300 208768 67312
rect 175056 67272 176700 67300
rect 176764 67272 208768 67300
rect 175056 67260 175062 67272
rect 107286 67232 107292 67244
rect 103486 67204 107292 67232
rect 80054 66852 80060 66904
rect 80112 66892 80118 66904
rect 103486 66892 103514 67204
rect 107286 67192 107292 67204
rect 107344 67232 107350 67244
rect 138290 67232 138296 67244
rect 107344 67204 138296 67232
rect 107344 67192 107350 67204
rect 138290 67192 138296 67204
rect 138348 67192 138354 67244
rect 174814 67192 174820 67244
rect 174872 67232 174878 67244
rect 176764 67232 176792 67272
rect 208762 67260 208768 67272
rect 208820 67260 208826 67312
rect 174872 67204 176792 67232
rect 174872 67192 174878 67204
rect 177114 67192 177120 67244
rect 177172 67232 177178 67244
rect 207290 67232 207296 67244
rect 177172 67204 207296 67232
rect 177172 67192 177178 67204
rect 207290 67192 207296 67204
rect 207348 67192 207354 67244
rect 108298 67124 108304 67176
rect 108356 67164 108362 67176
rect 138842 67164 138848 67176
rect 108356 67136 138848 67164
rect 108356 67124 108362 67136
rect 138842 67124 138848 67136
rect 138900 67124 138906 67176
rect 150618 67164 150624 67176
rect 147646 67136 150624 67164
rect 122466 67056 122472 67108
rect 122524 67096 122530 67108
rect 147646 67096 147674 67136
rect 150618 67124 150624 67136
rect 150676 67124 150682 67176
rect 176470 67124 176476 67176
rect 176528 67164 176534 67176
rect 210050 67164 210056 67176
rect 176528 67136 210056 67164
rect 176528 67124 176534 67136
rect 210050 67124 210056 67136
rect 210108 67124 210114 67176
rect 122524 67068 147674 67096
rect 122524 67056 122530 67068
rect 149146 67056 149152 67108
rect 149204 67096 149210 67108
rect 149882 67096 149888 67108
rect 149204 67068 149888 67096
rect 149204 67056 149210 67068
rect 149882 67056 149888 67068
rect 149940 67056 149946 67108
rect 154390 67056 154396 67108
rect 154448 67096 154454 67108
rect 274634 67096 274640 67108
rect 154448 67068 274640 67096
rect 154448 67056 154454 67068
rect 274634 67056 274640 67068
rect 274692 67056 274698 67108
rect 162486 66988 162492 67040
rect 162544 67028 162550 67040
rect 189442 67028 189448 67040
rect 162544 67000 189448 67028
rect 162544 66988 162550 67000
rect 189442 66988 189448 67000
rect 189500 67028 189506 67040
rect 317414 67028 317420 67040
rect 189500 67000 317420 67028
rect 189500 66988 189506 67000
rect 317414 66988 317420 67000
rect 317472 66988 317478 67040
rect 176286 66920 176292 66972
rect 176344 66960 176350 66972
rect 209958 66960 209964 66972
rect 176344 66932 209964 66960
rect 176344 66920 176350 66932
rect 209958 66920 209964 66932
rect 210016 66920 210022 66972
rect 213822 66920 213828 66972
rect 213880 66960 213886 66972
rect 529934 66960 529940 66972
rect 213880 66932 529940 66960
rect 213880 66920 213886 66932
rect 529934 66920 529940 66932
rect 529992 66920 529998 66972
rect 80112 66864 103514 66892
rect 80112 66852 80118 66864
rect 147858 66852 147864 66904
rect 147916 66892 147922 66904
rect 203518 66892 203524 66904
rect 147916 66864 203524 66892
rect 147916 66852 147922 66864
rect 203518 66852 203524 66864
rect 203576 66852 203582 66904
rect 215570 66852 215576 66904
rect 215628 66892 215634 66904
rect 545758 66892 545764 66904
rect 215628 66864 545764 66892
rect 215628 66852 215634 66864
rect 545758 66852 545764 66864
rect 545816 66852 545822 66904
rect 153470 66784 153476 66836
rect 153528 66824 153534 66836
rect 154482 66824 154488 66836
rect 153528 66796 154488 66824
rect 153528 66784 153534 66796
rect 154482 66784 154488 66796
rect 154540 66784 154546 66836
rect 174722 66784 174728 66836
rect 174780 66824 174786 66836
rect 207382 66824 207388 66836
rect 174780 66796 207388 66824
rect 174780 66784 174786 66796
rect 207382 66784 207388 66796
rect 207440 66784 207446 66836
rect 173618 66716 173624 66768
rect 173676 66756 173682 66768
rect 177114 66756 177120 66768
rect 173676 66728 177120 66756
rect 173676 66716 173682 66728
rect 177114 66716 177120 66728
rect 177172 66716 177178 66768
rect 173434 66648 173440 66700
rect 173492 66688 173498 66700
rect 177206 66688 177212 66700
rect 173492 66660 177212 66688
rect 173492 66648 173498 66660
rect 177206 66648 177212 66660
rect 177264 66648 177270 66700
rect 143994 66512 144000 66564
rect 144052 66552 144058 66564
rect 147214 66552 147220 66564
rect 144052 66524 147220 66552
rect 144052 66512 144058 66524
rect 147214 66512 147220 66524
rect 147272 66512 147278 66564
rect 141510 66240 141516 66292
rect 141568 66280 141574 66292
rect 142338 66280 142344 66292
rect 141568 66252 142344 66280
rect 141568 66240 141574 66252
rect 142338 66240 142344 66252
rect 142396 66240 142402 66292
rect 100754 66172 100760 66224
rect 100812 66212 100818 66224
rect 101674 66212 101680 66224
rect 100812 66184 101680 66212
rect 100812 66172 100818 66184
rect 101674 66172 101680 66184
rect 101732 66212 101738 66224
rect 134334 66212 134340 66224
rect 101732 66184 134340 66212
rect 101732 66172 101738 66184
rect 134334 66172 134340 66184
rect 134392 66172 134398 66224
rect 161750 66172 161756 66224
rect 161808 66212 161814 66224
rect 162486 66212 162492 66224
rect 161808 66184 162492 66212
rect 161808 66172 161814 66184
rect 162486 66172 162492 66184
rect 162544 66172 162550 66224
rect 164510 66172 164516 66224
rect 164568 66212 164574 66224
rect 165246 66212 165252 66224
rect 164568 66184 165252 66212
rect 164568 66172 164574 66184
rect 165246 66172 165252 66184
rect 165304 66172 165310 66224
rect 168650 66172 168656 66224
rect 168708 66212 168714 66224
rect 169570 66212 169576 66224
rect 168708 66184 169576 66212
rect 168708 66172 168714 66184
rect 169570 66172 169576 66184
rect 169628 66172 169634 66224
rect 210142 66212 210148 66224
rect 169680 66184 210148 66212
rect 100018 66104 100024 66156
rect 100076 66144 100082 66156
rect 134150 66144 134156 66156
rect 100076 66116 134156 66144
rect 100076 66104 100082 66116
rect 134150 66104 134156 66116
rect 134208 66104 134214 66156
rect 142338 66104 142344 66156
rect 142396 66144 142402 66156
rect 142982 66144 142988 66156
rect 142396 66116 142988 66144
rect 142396 66104 142402 66116
rect 142982 66104 142988 66116
rect 143040 66104 143046 66156
rect 162504 66144 162532 66172
rect 169680 66144 169708 66184
rect 210142 66172 210148 66184
rect 210200 66172 210206 66224
rect 162504 66116 169708 66144
rect 170214 66104 170220 66156
rect 170272 66144 170278 66156
rect 209038 66144 209044 66156
rect 170272 66116 209044 66144
rect 170272 66104 170278 66116
rect 209038 66104 209044 66116
rect 209096 66104 209102 66156
rect 100110 66036 100116 66088
rect 100168 66076 100174 66088
rect 134058 66076 134064 66088
rect 100168 66048 134064 66076
rect 100168 66036 100174 66048
rect 134058 66036 134064 66048
rect 134116 66076 134122 66088
rect 134794 66076 134800 66088
rect 134116 66048 134800 66076
rect 134116 66036 134122 66048
rect 134794 66036 134800 66048
rect 134852 66036 134858 66088
rect 161658 66036 161664 66088
rect 161716 66076 161722 66088
rect 162578 66076 162584 66088
rect 161716 66048 162584 66076
rect 161716 66036 161722 66048
rect 162578 66036 162584 66048
rect 162636 66036 162642 66088
rect 165246 66036 165252 66088
rect 165304 66076 165310 66088
rect 205818 66076 205824 66088
rect 165304 66048 205824 66076
rect 165304 66036 165310 66048
rect 205818 66036 205824 66048
rect 205876 66036 205882 66088
rect 102686 65968 102692 66020
rect 102744 66008 102750 66020
rect 135530 66008 135536 66020
rect 102744 65980 135536 66008
rect 102744 65968 102750 65980
rect 135530 65968 135536 65980
rect 135588 65968 135594 66020
rect 165890 65968 165896 66020
rect 165948 66008 165954 66020
rect 200298 66008 200304 66020
rect 165948 65980 200304 66008
rect 165948 65968 165954 65980
rect 200298 65968 200304 65980
rect 200356 66008 200362 66020
rect 201402 66008 201408 66020
rect 200356 65980 201408 66008
rect 200356 65968 200362 65980
rect 201402 65968 201408 65980
rect 201460 65968 201466 66020
rect 99466 65900 99472 65952
rect 99524 65940 99530 65952
rect 100478 65940 100484 65952
rect 99524 65912 100484 65940
rect 99524 65900 99530 65912
rect 100478 65900 100484 65912
rect 100536 65940 100542 65952
rect 133046 65940 133052 65952
rect 100536 65912 133052 65940
rect 100536 65900 100542 65912
rect 133046 65900 133052 65912
rect 133104 65900 133110 65952
rect 154942 65900 154948 65952
rect 155000 65940 155006 65952
rect 189074 65940 189080 65952
rect 155000 65912 189080 65940
rect 155000 65900 155006 65912
rect 189074 65900 189080 65912
rect 189132 65900 189138 65952
rect 119706 65832 119712 65884
rect 119764 65872 119770 65884
rect 150526 65872 150532 65884
rect 119764 65844 150532 65872
rect 119764 65832 119770 65844
rect 150526 65832 150532 65844
rect 150584 65832 150590 65884
rect 162578 65832 162584 65884
rect 162636 65872 162642 65884
rect 170214 65872 170220 65884
rect 162636 65844 170220 65872
rect 162636 65832 162642 65844
rect 170214 65832 170220 65844
rect 170272 65832 170278 65884
rect 185578 65832 185584 65884
rect 185636 65872 185642 65884
rect 214834 65872 214840 65884
rect 185636 65844 214840 65872
rect 185636 65832 185642 65844
rect 214834 65832 214840 65844
rect 214892 65872 214898 65884
rect 214892 65844 219434 65872
rect 214892 65832 214898 65844
rect 108942 65764 108948 65816
rect 109000 65804 109006 65816
rect 140130 65804 140136 65816
rect 109000 65776 140136 65804
rect 109000 65764 109006 65776
rect 140130 65764 140136 65776
rect 140188 65764 140194 65816
rect 177022 65764 177028 65816
rect 177080 65804 177086 65816
rect 203610 65804 203616 65816
rect 177080 65776 203616 65804
rect 177080 65764 177086 65776
rect 203610 65764 203616 65776
rect 203668 65804 203674 65816
rect 204162 65804 204168 65816
rect 203668 65776 204168 65804
rect 203668 65764 203674 65776
rect 204162 65764 204168 65776
rect 204220 65764 204226 65816
rect 124122 65696 124128 65748
rect 124180 65736 124186 65748
rect 161566 65736 161572 65748
rect 124180 65708 161572 65736
rect 124180 65696 124186 65708
rect 161566 65696 161572 65708
rect 161624 65736 161630 65748
rect 162118 65736 162124 65748
rect 161624 65708 162124 65736
rect 161624 65696 161630 65708
rect 162118 65696 162124 65708
rect 162176 65696 162182 65748
rect 169570 65696 169576 65748
rect 169628 65736 169634 65748
rect 186774 65736 186780 65748
rect 169628 65708 186780 65736
rect 169628 65696 169634 65708
rect 186774 65696 186780 65708
rect 186832 65696 186838 65748
rect 219406 65736 219434 65844
rect 238754 65736 238760 65748
rect 219406 65708 238760 65736
rect 238754 65696 238760 65708
rect 238812 65696 238818 65748
rect 149422 65628 149428 65680
rect 149480 65668 149486 65680
rect 223574 65668 223580 65680
rect 149480 65640 223580 65668
rect 149480 65628 149486 65640
rect 223574 65628 223580 65640
rect 223632 65628 223638 65680
rect 35986 65560 35992 65612
rect 36044 65600 36050 65612
rect 100754 65600 100760 65612
rect 36044 65572 100760 65600
rect 36044 65560 36050 65572
rect 100754 65560 100760 65572
rect 100812 65560 100818 65612
rect 189074 65560 189080 65612
rect 189132 65600 189138 65612
rect 295334 65600 295340 65612
rect 189132 65572 295340 65600
rect 189132 65560 189138 65572
rect 295334 65560 295340 65572
rect 295392 65560 295398 65612
rect 8294 65492 8300 65544
rect 8352 65532 8358 65544
rect 99466 65532 99472 65544
rect 8352 65504 99472 65532
rect 8352 65492 8358 65504
rect 99466 65492 99472 65504
rect 99524 65492 99530 65544
rect 112162 65492 112168 65544
rect 112220 65532 112226 65544
rect 131482 65532 131488 65544
rect 112220 65504 131488 65532
rect 112220 65492 112226 65504
rect 131482 65492 131488 65504
rect 131540 65532 131546 65544
rect 141142 65532 141148 65544
rect 131540 65504 141148 65532
rect 131540 65492 131546 65504
rect 141142 65492 141148 65504
rect 141200 65492 141206 65544
rect 201402 65492 201408 65544
rect 201460 65532 201466 65544
rect 432598 65532 432604 65544
rect 201460 65504 432604 65532
rect 201460 65492 201466 65504
rect 432598 65492 432604 65504
rect 432656 65492 432662 65544
rect 150526 65424 150532 65476
rect 150584 65464 150590 65476
rect 151262 65464 151268 65476
rect 150584 65436 151268 65464
rect 150584 65424 150590 65436
rect 151262 65424 151268 65436
rect 151320 65424 151326 65476
rect 142522 65356 142528 65408
rect 142580 65396 142586 65408
rect 142798 65396 142804 65408
rect 142580 65368 142804 65396
rect 142580 65356 142586 65368
rect 142798 65356 142804 65368
rect 142856 65356 142862 65408
rect 204162 64880 204168 64932
rect 204220 64920 204226 64932
rect 570598 64920 570604 64932
rect 204220 64892 570604 64920
rect 204220 64880 204226 64892
rect 570598 64880 570604 64892
rect 570656 64880 570662 64932
rect 104250 64812 104256 64864
rect 104308 64852 104314 64864
rect 137462 64852 137468 64864
rect 104308 64824 137468 64852
rect 104308 64812 104314 64824
rect 137462 64812 137468 64824
rect 137520 64812 137526 64864
rect 165706 64812 165712 64864
rect 165764 64852 165770 64864
rect 200850 64852 200856 64864
rect 165764 64824 200856 64852
rect 165764 64812 165770 64824
rect 200850 64812 200856 64824
rect 200908 64812 200914 64864
rect 104618 64744 104624 64796
rect 104676 64784 104682 64796
rect 137094 64784 137100 64796
rect 104676 64756 137100 64784
rect 104676 64744 104682 64756
rect 137094 64744 137100 64756
rect 137152 64744 137158 64796
rect 153102 64744 153108 64796
rect 153160 64784 153166 64796
rect 186590 64784 186596 64796
rect 153160 64756 186596 64784
rect 153160 64744 153166 64756
rect 186590 64744 186596 64756
rect 186648 64744 186654 64796
rect 165338 64676 165344 64728
rect 165396 64716 165402 64728
rect 199930 64716 199936 64728
rect 165396 64688 199936 64716
rect 165396 64676 165402 64688
rect 199930 64676 199936 64688
rect 199988 64676 199994 64728
rect 166534 64608 166540 64660
rect 166592 64648 166598 64660
rect 200390 64648 200396 64660
rect 166592 64620 200396 64648
rect 166592 64608 166598 64620
rect 200390 64608 200396 64620
rect 200448 64608 200454 64660
rect 158990 64540 158996 64592
rect 159048 64580 159054 64592
rect 193306 64580 193312 64592
rect 159048 64552 193312 64580
rect 159048 64540 159054 64552
rect 193306 64540 193312 64552
rect 193364 64540 193370 64592
rect 168558 64472 168564 64524
rect 168616 64512 168622 64524
rect 202874 64512 202880 64524
rect 168616 64484 202880 64512
rect 168616 64472 168622 64484
rect 202874 64472 202880 64484
rect 202932 64472 202938 64524
rect 171410 64404 171416 64456
rect 171468 64444 171474 64456
rect 187142 64444 187148 64456
rect 171468 64416 187148 64444
rect 171468 64404 171474 64416
rect 187142 64404 187148 64416
rect 187200 64404 187206 64456
rect 186590 64336 186596 64388
rect 186648 64376 186654 64388
rect 256694 64376 256700 64388
rect 186648 64348 256700 64376
rect 186648 64336 186654 64348
rect 256694 64336 256700 64348
rect 256752 64336 256758 64388
rect 149606 64268 149612 64320
rect 149664 64308 149670 64320
rect 220078 64308 220084 64320
rect 149664 64280 220084 64308
rect 149664 64268 149670 64280
rect 220078 64268 220084 64280
rect 220136 64268 220142 64320
rect 193306 64200 193312 64252
rect 193364 64240 193370 64252
rect 345014 64240 345020 64252
rect 193364 64212 345020 64240
rect 193364 64200 193370 64212
rect 345014 64200 345020 64212
rect 345072 64200 345078 64252
rect 62114 64132 62120 64184
rect 62172 64172 62178 64184
rect 104618 64172 104624 64184
rect 62172 64144 104624 64172
rect 62172 64132 62178 64144
rect 104618 64132 104624 64144
rect 104676 64132 104682 64184
rect 146846 64132 146852 64184
rect 146904 64172 146910 64184
rect 183554 64172 183560 64184
rect 146904 64144 183560 64172
rect 146904 64132 146910 64144
rect 183554 64132 183560 64144
rect 183612 64132 183618 64184
rect 202874 64132 202880 64184
rect 202932 64172 202938 64184
rect 472618 64172 472624 64184
rect 202932 64144 472624 64172
rect 202932 64132 202938 64144
rect 472618 64132 472624 64144
rect 472676 64132 472682 64184
rect 165798 63996 165804 64048
rect 165856 64036 165862 64048
rect 166534 64036 166540 64048
rect 165856 64008 166540 64036
rect 165856 63996 165862 64008
rect 166534 63996 166540 64008
rect 166592 63996 166598 64048
rect 164418 63860 164424 63912
rect 164476 63900 164482 63912
rect 165338 63900 165344 63912
rect 164476 63872 165344 63900
rect 164476 63860 164482 63872
rect 165338 63860 165344 63872
rect 165396 63860 165402 63912
rect 146018 63588 146024 63640
rect 146076 63628 146082 63640
rect 149790 63628 149796 63640
rect 146076 63600 149796 63628
rect 146076 63588 146082 63600
rect 149790 63588 149796 63600
rect 149848 63588 149854 63640
rect 165706 63520 165712 63572
rect 165764 63560 165770 63572
rect 166442 63560 166448 63572
rect 165764 63532 166448 63560
rect 165764 63520 165770 63532
rect 166442 63520 166448 63532
rect 166500 63520 166506 63572
rect 187142 63520 187148 63572
rect 187200 63560 187206 63572
rect 511994 63560 512000 63572
rect 187200 63532 512000 63560
rect 187200 63520 187206 63532
rect 511994 63520 512000 63532
rect 512052 63520 512058 63572
rect 164326 63452 164332 63504
rect 164384 63492 164390 63504
rect 199010 63492 199016 63504
rect 164384 63464 199016 63492
rect 164384 63452 164390 63464
rect 199010 63452 199016 63464
rect 199068 63492 199074 63504
rect 199194 63492 199200 63504
rect 199068 63464 199200 63492
rect 199068 63452 199074 63464
rect 199194 63452 199200 63464
rect 199252 63452 199258 63504
rect 143810 63384 143816 63436
rect 143868 63424 143874 63436
rect 148410 63424 148416 63436
rect 143868 63396 148416 63424
rect 143868 63384 143874 63396
rect 148410 63384 148416 63396
rect 148468 63384 148474 63436
rect 154758 63384 154764 63436
rect 154816 63424 154822 63436
rect 189074 63424 189080 63436
rect 154816 63396 189080 63424
rect 154816 63384 154822 63396
rect 189074 63384 189080 63396
rect 189132 63384 189138 63436
rect 151722 62908 151728 62960
rect 151780 62948 151786 62960
rect 245654 62948 245660 62960
rect 151780 62920 245660 62948
rect 151780 62908 151786 62920
rect 245654 62908 245660 62920
rect 245712 62908 245718 62960
rect 189074 62840 189080 62892
rect 189132 62880 189138 62892
rect 189994 62880 190000 62892
rect 189132 62852 190000 62880
rect 189132 62840 189138 62852
rect 189994 62840 190000 62852
rect 190052 62880 190058 62892
rect 292574 62880 292580 62892
rect 190052 62852 292580 62880
rect 190052 62840 190058 62852
rect 292574 62840 292580 62852
rect 292632 62840 292638 62892
rect 199194 62772 199200 62824
rect 199252 62812 199258 62824
rect 412634 62812 412640 62824
rect 199252 62784 412640 62812
rect 199252 62772 199258 62784
rect 412634 62772 412640 62784
rect 412692 62772 412698 62824
rect 102226 62024 102232 62076
rect 102284 62064 102290 62076
rect 103330 62064 103336 62076
rect 102284 62036 103336 62064
rect 102284 62024 102290 62036
rect 103330 62024 103336 62036
rect 103388 62064 103394 62076
rect 136174 62064 136180 62076
rect 103388 62036 136180 62064
rect 103388 62024 103394 62036
rect 136174 62024 136180 62036
rect 136232 62024 136238 62076
rect 167270 62024 167276 62076
rect 167328 62064 167334 62076
rect 202046 62064 202052 62076
rect 167328 62036 202052 62064
rect 167328 62024 167334 62036
rect 202046 62024 202052 62036
rect 202104 62064 202110 62076
rect 202782 62064 202788 62076
rect 202104 62036 202788 62064
rect 202104 62024 202110 62036
rect 202782 62024 202788 62036
rect 202840 62024 202846 62076
rect 102134 61956 102140 62008
rect 102192 61996 102198 62008
rect 102686 61996 102692 62008
rect 102192 61968 102692 61996
rect 102192 61956 102198 61968
rect 102686 61956 102692 61968
rect 102744 61996 102750 62008
rect 134426 61996 134432 62008
rect 102744 61968 134432 61996
rect 102744 61956 102750 61968
rect 134426 61956 134432 61968
rect 134484 61956 134490 62008
rect 156138 61956 156144 62008
rect 156196 61996 156202 62008
rect 190546 61996 190552 62008
rect 156196 61968 190552 61996
rect 156196 61956 156202 61968
rect 190546 61956 190552 61968
rect 190604 61996 190610 62008
rect 191742 61996 191748 62008
rect 190604 61968 191748 61996
rect 190604 61956 190610 61968
rect 191742 61956 191748 61968
rect 191800 61956 191806 62008
rect 163038 61888 163044 61940
rect 163096 61928 163102 61940
rect 197354 61928 197360 61940
rect 163096 61900 197360 61928
rect 163096 61888 163102 61900
rect 197354 61888 197360 61900
rect 197412 61888 197418 61940
rect 175458 61820 175464 61872
rect 175516 61860 175522 61872
rect 199102 61860 199108 61872
rect 175516 61832 199108 61860
rect 175516 61820 175522 61832
rect 199102 61820 199108 61832
rect 199160 61820 199166 61872
rect 148962 61616 148968 61668
rect 149020 61656 149026 61668
rect 197630 61656 197636 61668
rect 149020 61628 197636 61656
rect 149020 61616 149026 61628
rect 197630 61616 197636 61628
rect 197688 61616 197694 61668
rect 191742 61548 191748 61600
rect 191800 61588 191806 61600
rect 313274 61588 313280 61600
rect 191800 61560 313280 61588
rect 191800 61548 191806 61560
rect 313274 61548 313280 61560
rect 313332 61548 313338 61600
rect 154206 61480 154212 61532
rect 154264 61520 154270 61532
rect 277394 61520 277400 61532
rect 154264 61492 277400 61520
rect 154264 61480 154270 61492
rect 277394 61480 277400 61492
rect 277452 61480 277458 61532
rect 197354 61412 197360 61464
rect 197412 61452 197418 61464
rect 398834 61452 398840 61464
rect 197412 61424 398840 61452
rect 197412 61412 197418 61424
rect 398834 61412 398840 61424
rect 398892 61412 398898 61464
rect 43438 61344 43444 61396
rect 43496 61384 43502 61396
rect 102226 61384 102232 61396
rect 43496 61356 102232 61384
rect 43496 61344 43502 61356
rect 102226 61344 102232 61356
rect 102284 61344 102290 61396
rect 202782 61344 202788 61396
rect 202840 61384 202846 61396
rect 459554 61384 459560 61396
rect 202840 61356 459560 61384
rect 202840 61344 202846 61356
rect 459554 61344 459560 61356
rect 459612 61344 459618 61396
rect 199102 60732 199108 60784
rect 199160 60772 199166 60784
rect 563698 60772 563704 60784
rect 199160 60744 563704 60772
rect 199160 60732 199166 60744
rect 563698 60732 563704 60744
rect 563756 60732 563762 60784
rect 98914 60664 98920 60716
rect 98972 60704 98978 60716
rect 132954 60704 132960 60716
rect 98972 60676 132960 60704
rect 98972 60664 98978 60676
rect 132954 60664 132960 60676
rect 133012 60664 133018 60716
rect 154666 60664 154672 60716
rect 154724 60704 154730 60716
rect 214190 60704 214196 60716
rect 154724 60676 214196 60704
rect 154724 60664 154730 60676
rect 214190 60664 214196 60676
rect 214248 60704 214254 60716
rect 214466 60704 214472 60716
rect 214248 60676 214472 60704
rect 214248 60664 214254 60676
rect 214466 60664 214472 60676
rect 214524 60664 214530 60716
rect 102134 60596 102140 60648
rect 102192 60636 102198 60648
rect 103422 60636 103428 60648
rect 102192 60608 103428 60636
rect 102192 60596 102198 60608
rect 103422 60596 103428 60608
rect 103480 60636 103486 60648
rect 135714 60636 135720 60648
rect 103480 60608 135720 60636
rect 103480 60596 103486 60608
rect 135714 60596 135720 60608
rect 135772 60596 135778 60648
rect 158898 60596 158904 60648
rect 158956 60636 158962 60648
rect 193398 60636 193404 60648
rect 158956 60608 193404 60636
rect 158956 60596 158962 60608
rect 193398 60596 193404 60608
rect 193456 60636 193462 60648
rect 194502 60636 194508 60648
rect 193456 60608 194508 60636
rect 193456 60596 193462 60608
rect 194502 60596 194508 60608
rect 194560 60596 194566 60648
rect 111794 60528 111800 60580
rect 111852 60568 111858 60580
rect 112254 60568 112260 60580
rect 111852 60540 112260 60568
rect 111852 60528 111858 60540
rect 112254 60528 112260 60540
rect 112312 60568 112318 60580
rect 139854 60568 139860 60580
rect 112312 60540 139860 60568
rect 112312 60528 112318 60540
rect 139854 60528 139860 60540
rect 139912 60528 139918 60580
rect 166350 60528 166356 60580
rect 166408 60568 166414 60580
rect 196250 60568 196256 60580
rect 166408 60540 196256 60568
rect 166408 60528 166414 60540
rect 196250 60528 196256 60540
rect 196308 60528 196314 60580
rect 214466 60120 214472 60172
rect 214524 60160 214530 60172
rect 299474 60160 299480 60172
rect 214524 60132 299480 60160
rect 214524 60120 214530 60132
rect 299474 60120 299480 60132
rect 299532 60120 299538 60172
rect 44174 60052 44180 60104
rect 44232 60092 44238 60104
rect 102134 60092 102140 60104
rect 44232 60064 102140 60092
rect 44232 60052 44238 60064
rect 102134 60052 102140 60064
rect 102192 60052 102198 60104
rect 194502 60052 194508 60104
rect 194560 60092 194566 60104
rect 351914 60092 351920 60104
rect 194560 60064 351920 60092
rect 194560 60052 194566 60064
rect 351914 60052 351920 60064
rect 351972 60052 351978 60104
rect 21358 59984 21364 60036
rect 21416 60024 21422 60036
rect 98914 60024 98920 60036
rect 21416 59996 98920 60024
rect 21416 59984 21422 59996
rect 98914 59984 98920 59996
rect 98972 59984 98978 60036
rect 196250 59984 196256 60036
rect 196308 60024 196314 60036
rect 196894 60024 196900 60036
rect 196308 59996 196900 60024
rect 196308 59984 196314 59996
rect 196894 59984 196900 59996
rect 196952 60024 196958 60036
rect 402974 60024 402980 60036
rect 196952 59996 402980 60024
rect 196952 59984 196958 59996
rect 402974 59984 402980 59996
rect 403032 59984 403038 60036
rect 3510 59304 3516 59356
rect 3568 59344 3574 59356
rect 40678 59344 40684 59356
rect 3568 59316 40684 59344
rect 3568 59304 3574 59316
rect 40678 59304 40684 59316
rect 40736 59304 40742 59356
rect 109862 59304 109868 59356
rect 109920 59344 109926 59356
rect 110414 59344 110420 59356
rect 109920 59316 110420 59344
rect 109920 59304 109926 59316
rect 110414 59304 110420 59316
rect 110472 59304 110478 59356
rect 135806 59344 135812 59356
rect 110616 59316 135812 59344
rect 104158 59168 104164 59220
rect 104216 59208 104222 59220
rect 110616 59208 110644 59316
rect 135806 59304 135812 59316
rect 135864 59304 135870 59356
rect 161474 59304 161480 59356
rect 161532 59344 161538 59356
rect 196250 59344 196256 59356
rect 161532 59316 196256 59344
rect 161532 59304 161538 59316
rect 196250 59304 196256 59316
rect 196308 59344 196314 59356
rect 196526 59344 196532 59356
rect 196308 59316 196532 59344
rect 196308 59304 196314 59316
rect 196526 59304 196532 59316
rect 196584 59304 196590 59356
rect 137002 59276 137008 59288
rect 104216 59180 110644 59208
rect 113146 59248 137008 59276
rect 104216 59168 104222 59180
rect 105998 59100 106004 59152
rect 106056 59140 106062 59152
rect 106182 59140 106188 59152
rect 106056 59112 106188 59140
rect 106056 59100 106062 59112
rect 106182 59100 106188 59112
rect 106240 59140 106246 59152
rect 113146 59140 113174 59248
rect 137002 59236 137008 59248
rect 137060 59236 137066 59288
rect 157426 59236 157432 59288
rect 157484 59276 157490 59288
rect 192110 59276 192116 59288
rect 157484 59248 192116 59276
rect 157484 59236 157490 59248
rect 192110 59236 192116 59248
rect 192168 59276 192174 59288
rect 193030 59276 193036 59288
rect 192168 59248 193036 59276
rect 192168 59236 192174 59248
rect 193030 59236 193036 59248
rect 193088 59236 193094 59288
rect 106240 59112 113174 59140
rect 106240 59100 106246 59112
rect 148686 58896 148692 58948
rect 148744 58936 148750 58948
rect 198734 58936 198740 58948
rect 148744 58908 198740 58936
rect 148744 58896 148750 58908
rect 198734 58896 198740 58908
rect 198792 58896 198798 58948
rect 151630 58828 151636 58880
rect 151688 58868 151694 58880
rect 249794 58868 249800 58880
rect 151688 58840 249800 58868
rect 151688 58828 151694 58840
rect 249794 58828 249800 58840
rect 249852 58828 249858 58880
rect 154114 58760 154120 58812
rect 154172 58800 154178 58812
rect 281534 58800 281540 58812
rect 154172 58772 281540 58800
rect 154172 58760 154178 58772
rect 281534 58760 281540 58772
rect 281592 58760 281598 58812
rect 193030 58692 193036 58744
rect 193088 58732 193094 58744
rect 327074 58732 327080 58744
rect 193088 58704 327080 58732
rect 193088 58692 193094 58704
rect 327074 58692 327080 58704
rect 327132 58692 327138 58744
rect 69014 58624 69020 58676
rect 69072 58664 69078 58676
rect 105998 58664 106004 58676
rect 69072 58636 106004 58664
rect 69072 58624 69078 58636
rect 105998 58624 106004 58636
rect 106056 58624 106062 58676
rect 196250 58624 196256 58676
rect 196308 58664 196314 58676
rect 380894 58664 380900 58676
rect 196308 58636 380900 58664
rect 196308 58624 196314 58636
rect 380894 58624 380900 58636
rect 380952 58624 380958 58676
rect 158806 57876 158812 57928
rect 158864 57916 158870 57928
rect 193214 57916 193220 57928
rect 158864 57888 193220 57916
rect 158864 57876 158870 57888
rect 193214 57876 193220 57888
rect 193272 57916 193278 57928
rect 194502 57916 194508 57928
rect 193272 57888 194508 57916
rect 193272 57876 193278 57888
rect 194502 57876 194508 57888
rect 194560 57876 194566 57928
rect 170122 57808 170128 57860
rect 170180 57848 170186 57860
rect 196250 57848 196256 57860
rect 170180 57820 196256 57848
rect 170180 57808 170186 57820
rect 196250 57808 196256 57820
rect 196308 57808 196314 57860
rect 194502 57196 194508 57248
rect 194560 57236 194566 57248
rect 349154 57236 349160 57248
rect 194560 57208 349160 57236
rect 194560 57196 194566 57208
rect 349154 57196 349160 57208
rect 349212 57196 349218 57248
rect 196250 56584 196256 56636
rect 196308 56624 196314 56636
rect 484394 56624 484400 56636
rect 196308 56596 484400 56624
rect 196308 56584 196314 56596
rect 484394 56584 484400 56596
rect 484452 56584 484458 56636
rect 113542 56516 113548 56568
rect 113600 56556 113606 56568
rect 138382 56556 138388 56568
rect 113600 56528 138388 56556
rect 113600 56516 113606 56528
rect 138382 56516 138388 56528
rect 138440 56516 138446 56568
rect 167178 56516 167184 56568
rect 167236 56556 167242 56568
rect 201586 56556 201592 56568
rect 167236 56528 201592 56556
rect 167236 56516 167242 56528
rect 201586 56516 201592 56528
rect 201644 56556 201650 56568
rect 202782 56556 202788 56568
rect 201644 56528 202788 56556
rect 201644 56516 201650 56528
rect 202782 56516 202788 56528
rect 202840 56516 202846 56568
rect 145098 55836 145104 55888
rect 145156 55876 145162 55888
rect 170398 55876 170404 55888
rect 145156 55848 170404 55876
rect 145156 55836 145162 55848
rect 170398 55836 170404 55848
rect 170456 55836 170462 55888
rect 202782 55836 202788 55888
rect 202840 55876 202846 55888
rect 450538 55876 450544 55888
rect 202840 55848 450544 55876
rect 202840 55836 202846 55848
rect 450538 55836 450544 55848
rect 450596 55836 450602 55888
rect 138658 55224 138664 55276
rect 138716 55264 138722 55276
rect 142338 55264 142344 55276
rect 138716 55236 142344 55264
rect 138716 55224 138722 55236
rect 142338 55224 142344 55236
rect 142396 55224 142402 55276
rect 156046 55156 156052 55208
rect 156104 55196 156110 55208
rect 190454 55196 190460 55208
rect 156104 55168 190460 55196
rect 156104 55156 156110 55168
rect 190454 55156 190460 55168
rect 190512 55196 190518 55208
rect 191742 55196 191748 55208
rect 190512 55168 191748 55196
rect 190512 55156 190518 55168
rect 191742 55156 191748 55168
rect 191800 55156 191806 55208
rect 176930 55088 176936 55140
rect 176988 55128 176994 55140
rect 203334 55128 203340 55140
rect 176988 55100 203340 55128
rect 176988 55088 176994 55100
rect 203334 55088 203340 55100
rect 203392 55088 203398 55140
rect 167914 55020 167920 55072
rect 167972 55060 167978 55072
rect 189350 55060 189356 55072
rect 167972 55032 189356 55060
rect 167972 55020 167978 55032
rect 189350 55020 189356 55032
rect 189408 55020 189414 55072
rect 151538 54612 151544 54664
rect 151596 54652 151602 54664
rect 239398 54652 239404 54664
rect 151596 54624 239404 54652
rect 151596 54612 151602 54624
rect 239398 54612 239404 54624
rect 239456 54612 239462 54664
rect 191742 54544 191748 54596
rect 191800 54584 191806 54596
rect 315298 54584 315304 54596
rect 191800 54556 315304 54584
rect 191800 54544 191806 54556
rect 315298 54544 315304 54556
rect 315356 54544 315362 54596
rect 189350 54476 189356 54528
rect 189408 54516 189414 54528
rect 382274 54516 382280 54528
rect 189408 54488 382280 54516
rect 189408 54476 189414 54488
rect 382274 54476 382280 54488
rect 382332 54476 382338 54528
rect 203978 53796 203984 53848
rect 204036 53836 204042 53848
rect 571978 53836 571984 53848
rect 204036 53808 571984 53836
rect 204036 53796 204042 53808
rect 571978 53796 571984 53808
rect 572036 53796 572042 53848
rect 162946 53728 162952 53780
rect 163004 53768 163010 53780
rect 198366 53768 198372 53780
rect 163004 53740 198372 53768
rect 163004 53728 163010 53740
rect 198366 53728 198372 53740
rect 198424 53728 198430 53780
rect 172514 53660 172520 53712
rect 172572 53700 172578 53712
rect 207198 53700 207204 53712
rect 172572 53672 207204 53700
rect 172572 53660 172578 53672
rect 207198 53660 207204 53672
rect 207256 53660 207262 53712
rect 165614 53592 165620 53644
rect 165672 53632 165678 53644
rect 198918 53632 198924 53644
rect 165672 53604 198924 53632
rect 165672 53592 165678 53604
rect 198918 53592 198924 53604
rect 198976 53632 198982 53644
rect 199102 53632 199108 53644
rect 198976 53604 199108 53632
rect 198976 53592 198982 53604
rect 199102 53592 199108 53604
rect 199160 53592 199166 53644
rect 198366 53184 198372 53236
rect 198424 53224 198430 53236
rect 391934 53224 391940 53236
rect 198424 53196 391940 53224
rect 198424 53184 198430 53196
rect 391934 53184 391940 53196
rect 391992 53184 391998 53236
rect 199102 53116 199108 53168
rect 199160 53156 199166 53168
rect 437474 53156 437480 53168
rect 199160 53128 437480 53156
rect 199160 53116 199166 53128
rect 437474 53116 437480 53128
rect 437532 53116 437538 53168
rect 145742 53048 145748 53100
rect 145800 53088 145806 53100
rect 163498 53088 163504 53100
rect 145800 53060 163504 53088
rect 145800 53048 145806 53060
rect 163498 53048 163504 53060
rect 163556 53048 163562 53100
rect 207198 53048 207204 53100
rect 207256 53088 207262 53100
rect 516778 53088 516784 53100
rect 207256 53060 516784 53088
rect 207256 53048 207262 53060
rect 516778 53048 516784 53060
rect 516836 53048 516842 53100
rect 158714 52368 158720 52420
rect 158772 52408 158778 52420
rect 193214 52408 193220 52420
rect 158772 52380 193220 52408
rect 158772 52368 158778 52380
rect 193214 52368 193220 52380
rect 193272 52408 193278 52420
rect 194502 52408 194508 52420
rect 193272 52380 194508 52408
rect 193272 52368 193278 52380
rect 194502 52368 194508 52380
rect 194560 52368 194566 52420
rect 162854 52300 162860 52352
rect 162912 52340 162918 52352
rect 197538 52340 197544 52352
rect 162912 52312 197544 52340
rect 162912 52300 162918 52312
rect 197538 52300 197544 52312
rect 197596 52340 197602 52352
rect 198090 52340 198096 52352
rect 197596 52312 198096 52340
rect 197596 52300 197602 52312
rect 198090 52300 198096 52312
rect 198148 52300 198154 52352
rect 168374 52232 168380 52284
rect 168432 52272 168438 52284
rect 201954 52272 201960 52284
rect 168432 52244 201960 52272
rect 168432 52232 168438 52244
rect 201954 52232 201960 52244
rect 202012 52272 202018 52284
rect 202782 52272 202788 52284
rect 202012 52244 202788 52272
rect 202012 52232 202018 52244
rect 202782 52232 202788 52244
rect 202840 52232 202846 52284
rect 143718 51688 143724 51740
rect 143776 51728 143782 51740
rect 157426 51728 157432 51740
rect 143776 51700 157432 51728
rect 143776 51688 143782 51700
rect 157426 51688 157432 51700
rect 157484 51688 157490 51740
rect 198090 51688 198096 51740
rect 198148 51728 198154 51740
rect 400858 51728 400864 51740
rect 198148 51700 400864 51728
rect 198148 51688 198154 51700
rect 400858 51688 400864 51700
rect 400916 51688 400922 51740
rect 194502 51144 194508 51196
rect 194560 51184 194566 51196
rect 356054 51184 356060 51196
rect 194560 51156 356060 51184
rect 194560 51144 194566 51156
rect 356054 51144 356060 51156
rect 356112 51144 356118 51196
rect 202782 51076 202788 51128
rect 202840 51116 202846 51128
rect 464338 51116 464344 51128
rect 202840 51088 464344 51116
rect 202840 51076 202846 51088
rect 464338 51076 464344 51088
rect 464396 51076 464402 51128
rect 176838 51008 176844 51060
rect 176896 51048 176902 51060
rect 207198 51048 207204 51060
rect 176896 51020 207204 51048
rect 176896 51008 176902 51020
rect 207198 51008 207204 51020
rect 207256 51008 207262 51060
rect 150342 50328 150348 50380
rect 150400 50368 150406 50380
rect 225598 50368 225604 50380
rect 150400 50340 225604 50368
rect 150400 50328 150406 50340
rect 225598 50328 225604 50340
rect 225656 50328 225662 50380
rect 207198 49716 207204 49768
rect 207256 49756 207262 49768
rect 569954 49756 569960 49768
rect 207256 49728 569960 49756
rect 207256 49716 207262 49728
rect 569954 49716 569960 49728
rect 570012 49716 570018 49768
rect 166994 49648 167000 49700
rect 167052 49688 167058 49700
rect 201862 49688 201868 49700
rect 167052 49660 201868 49688
rect 167052 49648 167058 49660
rect 201862 49648 201868 49660
rect 201920 49688 201926 49700
rect 202782 49688 202788 49700
rect 201920 49660 202788 49688
rect 201920 49648 201926 49660
rect 202782 49648 202788 49660
rect 202840 49648 202846 49700
rect 147398 49172 147404 49224
rect 147456 49212 147462 49224
rect 186314 49212 186320 49224
rect 147456 49184 186320 49212
rect 147456 49172 147462 49184
rect 186314 49172 186320 49184
rect 186372 49172 186378 49224
rect 150250 49104 150256 49156
rect 150308 49144 150314 49156
rect 222194 49144 222200 49156
rect 150308 49116 222200 49144
rect 150308 49104 150314 49116
rect 222194 49104 222200 49116
rect 222252 49104 222258 49156
rect 147766 49036 147772 49088
rect 147824 49076 147830 49088
rect 201586 49076 201592 49088
rect 147824 49048 201592 49076
rect 147824 49036 147830 49048
rect 201586 49036 201592 49048
rect 201644 49036 201650 49088
rect 202782 49036 202788 49088
rect 202840 49076 202846 49088
rect 448606 49076 448612 49088
rect 202840 49048 448612 49076
rect 202840 49036 202846 49048
rect 448606 49036 448612 49048
rect 448664 49036 448670 49088
rect 133966 48968 133972 49020
rect 134024 49008 134030 49020
rect 142522 49008 142528 49020
rect 134024 48980 142528 49008
rect 134024 48968 134030 48980
rect 142522 48968 142528 48980
rect 142580 48968 142586 49020
rect 145006 48968 145012 49020
rect 145064 49008 145070 49020
rect 168374 49008 168380 49020
rect 145064 48980 168380 49008
rect 145064 48968 145070 48980
rect 168374 48968 168380 48980
rect 168432 48968 168438 49020
rect 172054 48968 172060 49020
rect 172112 49008 172118 49020
rect 502978 49008 502984 49020
rect 172112 48980 502984 49008
rect 172112 48968 172118 48980
rect 502978 48968 502984 48980
rect 503036 48968 503042 49020
rect 144362 48220 144368 48272
rect 144420 48260 144426 48272
rect 147674 48260 147680 48272
rect 144420 48232 147680 48260
rect 144420 48220 144426 48232
rect 147674 48220 147680 48232
rect 147732 48220 147738 48272
rect 147766 47676 147772 47728
rect 147824 47716 147830 47728
rect 208394 47716 208400 47728
rect 147824 47688 208400 47716
rect 147824 47676 147830 47688
rect 208394 47676 208400 47688
rect 208452 47676 208458 47728
rect 150158 47608 150164 47660
rect 150216 47648 150222 47660
rect 215294 47648 215300 47660
rect 150216 47620 215300 47648
rect 150216 47608 150222 47620
rect 215294 47608 215300 47620
rect 215352 47608 215358 47660
rect 169294 47540 169300 47592
rect 169352 47580 169358 47592
rect 468478 47580 468484 47592
rect 169352 47552 468484 47580
rect 169352 47540 169358 47552
rect 468478 47540 468484 47552
rect 468536 47540 468542 47592
rect 154574 46860 154580 46912
rect 154632 46900 154638 46912
rect 216766 46900 216772 46912
rect 154632 46872 216772 46900
rect 154632 46860 154638 46872
rect 216766 46860 216772 46872
rect 216824 46900 216830 46912
rect 217042 46900 217048 46912
rect 216824 46872 217048 46900
rect 216824 46860 216830 46872
rect 217042 46860 217048 46872
rect 217100 46860 217106 46912
rect 176746 46792 176752 46844
rect 176804 46832 176810 46844
rect 207198 46832 207204 46844
rect 176804 46804 207204 46832
rect 176804 46792 176810 46804
rect 207198 46792 207204 46804
rect 207256 46792 207262 46844
rect 145650 46180 145656 46232
rect 145708 46220 145714 46232
rect 166994 46220 167000 46232
rect 145708 46192 167000 46220
rect 145708 46180 145714 46192
rect 166994 46180 167000 46192
rect 167052 46180 167058 46232
rect 216766 46180 216772 46232
rect 216824 46220 216830 46232
rect 292666 46220 292672 46232
rect 216824 46192 292672 46220
rect 216824 46180 216830 46192
rect 292666 46180 292672 46192
rect 292724 46180 292730 46232
rect 207934 45568 207940 45620
rect 207992 45608 207998 45620
rect 560938 45608 560944 45620
rect 207992 45580 560944 45608
rect 207992 45568 207998 45580
rect 560938 45568 560944 45580
rect 560996 45568 561002 45620
rect 152918 44820 152924 44872
rect 152976 44860 152982 44872
rect 267734 44860 267740 44872
rect 152976 44832 267740 44860
rect 152976 44820 152982 44832
rect 267734 44820 267740 44832
rect 267792 44820 267798 44872
rect 177390 44072 177396 44124
rect 177448 44112 177454 44124
rect 211246 44112 211252 44124
rect 177448 44084 211252 44112
rect 177448 44072 177454 44084
rect 211246 44072 211252 44084
rect 211304 44112 211310 44124
rect 212442 44112 212448 44124
rect 211304 44084 212448 44112
rect 211304 44072 211310 44084
rect 212442 44072 212448 44084
rect 212500 44072 212506 44124
rect 151446 43460 151452 43512
rect 151504 43500 151510 43512
rect 233234 43500 233240 43512
rect 151504 43472 233240 43500
rect 151504 43460 151510 43472
rect 233234 43460 233240 43472
rect 233292 43460 233298 43512
rect 212442 43392 212448 43444
rect 212500 43432 212506 43444
rect 578234 43432 578240 43444
rect 212500 43404 578240 43432
rect 212500 43392 212506 43404
rect 578234 43392 578240 43404
rect 578292 43392 578298 43444
rect 149054 42304 149060 42356
rect 149112 42344 149118 42356
rect 218146 42344 218152 42356
rect 149112 42316 218152 42344
rect 149112 42304 149118 42316
rect 218146 42304 218152 42316
rect 218204 42304 218210 42356
rect 155310 42236 155316 42288
rect 155368 42276 155374 42288
rect 285674 42276 285680 42288
rect 155368 42248 285680 42276
rect 155368 42236 155374 42248
rect 285674 42236 285680 42248
rect 285732 42236 285738 42288
rect 165062 42168 165068 42220
rect 165120 42208 165126 42220
rect 426434 42208 426440 42220
rect 165120 42180 426440 42208
rect 165120 42168 165126 42180
rect 426434 42168 426440 42180
rect 426492 42168 426498 42220
rect 170030 42100 170036 42152
rect 170088 42140 170094 42152
rect 495434 42140 495440 42152
rect 170088 42112 495440 42140
rect 170088 42100 170094 42112
rect 495434 42100 495440 42112
rect 495492 42100 495498 42152
rect 70394 42032 70400 42084
rect 70452 42072 70458 42084
rect 136910 42072 136916 42084
rect 70452 42044 136916 42072
rect 70452 42032 70458 42044
rect 136910 42032 136916 42044
rect 136968 42032 136974 42084
rect 172146 42032 172152 42084
rect 172204 42072 172210 42084
rect 503714 42072 503720 42084
rect 172204 42044 503720 42072
rect 172204 42032 172210 42044
rect 503714 42032 503720 42044
rect 503772 42032 503778 42084
rect 148594 41012 148600 41064
rect 148652 41052 148658 41064
rect 204346 41052 204352 41064
rect 148652 41024 204352 41052
rect 148652 41012 148658 41024
rect 204346 41012 204352 41024
rect 204404 41012 204410 41064
rect 156690 40944 156696 40996
rect 156748 40984 156754 40996
rect 309134 40984 309140 40996
rect 156748 40956 309140 40984
rect 156748 40944 156754 40956
rect 309134 40944 309140 40956
rect 309192 40944 309198 40996
rect 158346 40876 158352 40928
rect 158404 40916 158410 40928
rect 332686 40916 332692 40928
rect 158404 40888 332692 40916
rect 158404 40876 158410 40888
rect 332686 40876 332692 40888
rect 332744 40876 332750 40928
rect 169938 40808 169944 40860
rect 169996 40848 170002 40860
rect 491294 40848 491300 40860
rect 169996 40820 491300 40848
rect 169996 40808 170002 40820
rect 491294 40808 491300 40820
rect 491352 40808 491358 40860
rect 171318 40740 171324 40792
rect 171376 40780 171382 40792
rect 498286 40780 498292 40792
rect 171376 40752 498292 40780
rect 171376 40740 171382 40752
rect 498286 40740 498292 40752
rect 498344 40740 498350 40792
rect 74534 40672 74540 40724
rect 74592 40712 74598 40724
rect 138106 40712 138112 40724
rect 74592 40684 138112 40712
rect 74592 40672 74598 40684
rect 138106 40672 138112 40684
rect 138164 40672 138170 40724
rect 174722 40672 174728 40724
rect 174780 40712 174786 40724
rect 549254 40712 549260 40724
rect 174780 40684 549260 40712
rect 174780 40672 174786 40684
rect 549254 40672 549260 40684
rect 549312 40672 549318 40724
rect 138106 39992 138112 40044
rect 138164 40032 138170 40044
rect 142246 40032 142252 40044
rect 138164 40004 142252 40032
rect 138164 39992 138170 40004
rect 142246 39992 142252 40004
rect 142304 39992 142310 40044
rect 150434 39584 150440 39636
rect 150492 39624 150498 39636
rect 235994 39624 236000 39636
rect 150492 39596 236000 39624
rect 150492 39584 150498 39596
rect 235994 39584 236000 39596
rect 236052 39584 236058 39636
rect 158254 39516 158260 39568
rect 158312 39556 158318 39568
rect 324406 39556 324412 39568
rect 158312 39528 324412 39556
rect 158312 39516 158318 39528
rect 324406 39516 324412 39528
rect 324464 39516 324470 39568
rect 169386 39448 169392 39500
rect 169444 39488 169450 39500
rect 463694 39488 463700 39500
rect 169444 39460 463700 39488
rect 169444 39448 169450 39460
rect 463694 39448 463700 39460
rect 463752 39448 463758 39500
rect 167086 39380 167092 39432
rect 167144 39420 167150 39432
rect 462314 39420 462320 39432
rect 167144 39392 462320 39420
rect 167144 39380 167150 39392
rect 462314 39380 462320 39392
rect 462372 39380 462378 39432
rect 77386 39312 77392 39364
rect 77444 39352 77450 39364
rect 138014 39352 138020 39364
rect 77444 39324 138020 39352
rect 77444 39312 77450 39324
rect 138014 39312 138020 39324
rect 138072 39312 138078 39364
rect 173526 39312 173532 39364
rect 173584 39352 173590 39364
rect 516134 39352 516140 39364
rect 173584 39324 516140 39352
rect 173584 39312 173590 39324
rect 516134 39312 516140 39324
rect 516192 39312 516198 39364
rect 145558 38156 145564 38208
rect 145616 38196 145622 38208
rect 168558 38196 168564 38208
rect 145616 38168 168564 38196
rect 145616 38156 145622 38168
rect 168558 38156 168564 38168
rect 168616 38156 168622 38208
rect 153010 38088 153016 38140
rect 153068 38128 153074 38140
rect 251266 38128 251272 38140
rect 153068 38100 251272 38128
rect 153068 38088 153074 38100
rect 251266 38088 251272 38100
rect 251324 38088 251330 38140
rect 169478 38020 169484 38072
rect 169536 38060 169542 38072
rect 470594 38060 470600 38072
rect 169536 38032 470600 38060
rect 169536 38020 169542 38032
rect 470594 38020 470600 38032
rect 470652 38020 470658 38072
rect 168466 37952 168472 38004
rect 168524 37992 168530 38004
rect 476114 37992 476120 38004
rect 168524 37964 476120 37992
rect 168524 37952 168530 37964
rect 476114 37952 476120 37964
rect 476172 37952 476178 38004
rect 13814 37884 13820 37936
rect 13872 37924 13878 37936
rect 132862 37924 132868 37936
rect 13872 37896 132868 37924
rect 13872 37884 13878 37896
rect 132862 37884 132868 37896
rect 132920 37884 132926 37936
rect 174906 37884 174912 37936
rect 174964 37924 174970 37936
rect 534074 37924 534080 37936
rect 174964 37896 534080 37924
rect 174964 37884 174970 37896
rect 534074 37884 534080 37896
rect 534132 37884 534138 37936
rect 154022 36660 154028 36712
rect 154080 36700 154086 36712
rect 267826 36700 267832 36712
rect 154080 36672 267832 36700
rect 154080 36660 154086 36672
rect 267826 36660 267832 36672
rect 267884 36660 267890 36712
rect 170858 36592 170864 36644
rect 170916 36632 170922 36644
rect 481634 36632 481640 36644
rect 170916 36604 481640 36632
rect 170916 36592 170922 36604
rect 481634 36592 481640 36604
rect 481692 36592 481698 36644
rect 95234 36524 95240 36576
rect 95292 36564 95298 36576
rect 139578 36564 139584 36576
rect 95292 36536 139584 36564
rect 95292 36524 95298 36536
rect 139578 36524 139584 36536
rect 139636 36524 139642 36576
rect 173434 36524 173440 36576
rect 173492 36564 173498 36576
rect 527818 36564 527824 36576
rect 173492 36536 527824 36564
rect 173492 36524 173498 36536
rect 527818 36524 527824 36536
rect 527876 36524 527882 36576
rect 158438 35368 158444 35420
rect 158496 35408 158502 35420
rect 321554 35408 321560 35420
rect 158496 35380 321560 35408
rect 158496 35368 158502 35380
rect 321554 35368 321560 35380
rect 321612 35368 321618 35420
rect 166442 35300 166448 35352
rect 166500 35340 166506 35352
rect 440326 35340 440332 35352
rect 166500 35312 440332 35340
rect 166500 35300 166506 35312
rect 440326 35300 440332 35312
rect 440384 35300 440390 35352
rect 174814 35232 174820 35284
rect 174872 35272 174878 35284
rect 538858 35272 538864 35284
rect 174872 35244 538864 35272
rect 174872 35232 174878 35244
rect 538858 35232 538864 35244
rect 538916 35232 538922 35284
rect 23474 35164 23480 35216
rect 23532 35204 23538 35216
rect 134150 35204 134156 35216
rect 23532 35176 134156 35204
rect 23532 35164 23538 35176
rect 134150 35164 134156 35176
rect 134208 35164 134214 35216
rect 176378 35164 176384 35216
rect 176436 35204 176442 35216
rect 558914 35204 558920 35216
rect 176436 35176 558920 35204
rect 176436 35164 176442 35176
rect 558914 35164 558920 35176
rect 558972 35164 558978 35216
rect 160830 33940 160836 33992
rect 160888 33980 160894 33992
rect 357434 33980 357440 33992
rect 160888 33952 357440 33980
rect 160888 33940 160894 33952
rect 357434 33940 357440 33952
rect 357492 33940 357498 33992
rect 162118 33872 162124 33924
rect 162176 33912 162182 33924
rect 378778 33912 378784 33924
rect 162176 33884 378784 33912
rect 162176 33872 162182 33884
rect 378778 33872 378784 33884
rect 378836 33872 378842 33924
rect 169846 33804 169852 33856
rect 169904 33844 169910 33856
rect 488534 33844 488540 33856
rect 169904 33816 488540 33844
rect 169904 33804 169910 33816
rect 488534 33804 488540 33816
rect 488592 33804 488598 33856
rect 31754 33736 31760 33788
rect 31812 33776 31818 33788
rect 134058 33776 134064 33788
rect 31812 33748 134064 33776
rect 31812 33736 31818 33748
rect 134058 33736 134064 33748
rect 134116 33736 134122 33788
rect 144270 33736 144276 33788
rect 144328 33776 144334 33788
rect 160094 33776 160100 33788
rect 144328 33748 160100 33776
rect 144328 33736 144334 33748
rect 160094 33736 160100 33748
rect 160152 33736 160158 33788
rect 177666 33736 177672 33788
rect 177724 33776 177730 33788
rect 576854 33776 576860 33788
rect 177724 33748 576860 33776
rect 177724 33736 177730 33748
rect 576854 33736 576860 33748
rect 576912 33736 576918 33788
rect 3510 33056 3516 33108
rect 3568 33096 3574 33108
rect 97258 33096 97264 33108
rect 3568 33068 97264 33096
rect 3568 33056 3574 33068
rect 97258 33056 97264 33068
rect 97316 33056 97322 33108
rect 148502 32648 148508 32700
rect 148560 32688 148566 32700
rect 205726 32688 205732 32700
rect 148560 32660 205732 32688
rect 148560 32648 148566 32660
rect 205726 32648 205732 32660
rect 205784 32648 205790 32700
rect 152826 32580 152832 32632
rect 152884 32620 152890 32632
rect 264974 32620 264980 32632
rect 152884 32592 264980 32620
rect 152884 32580 152890 32592
rect 264974 32580 264980 32592
rect 265032 32580 265038 32632
rect 159726 32512 159732 32564
rect 159784 32552 159790 32564
rect 346394 32552 346400 32564
rect 159784 32524 346400 32552
rect 159784 32512 159790 32524
rect 346394 32512 346400 32524
rect 346452 32512 346458 32564
rect 163774 32444 163780 32496
rect 163832 32484 163838 32496
rect 404354 32484 404360 32496
rect 163832 32456 404360 32484
rect 163832 32444 163838 32456
rect 404354 32444 404360 32456
rect 404412 32444 404418 32496
rect 170950 32376 170956 32428
rect 171008 32416 171014 32428
rect 492674 32416 492680 32428
rect 171008 32388 492680 32416
rect 171008 32376 171014 32388
rect 492674 32376 492680 32388
rect 492732 32376 492738 32428
rect 155770 31288 155776 31340
rect 155828 31328 155834 31340
rect 299566 31328 299572 31340
rect 155828 31300 299572 31328
rect 155828 31288 155834 31300
rect 299566 31288 299572 31300
rect 299624 31288 299630 31340
rect 160922 31220 160928 31272
rect 160980 31260 160986 31272
rect 360194 31260 360200 31272
rect 160980 31232 360200 31260
rect 160980 31220 160986 31232
rect 360194 31220 360200 31232
rect 360252 31220 360258 31272
rect 163866 31152 163872 31204
rect 163924 31192 163930 31204
rect 407206 31192 407212 31204
rect 163924 31164 407212 31192
rect 163924 31152 163930 31164
rect 407206 31152 407212 31164
rect 407264 31152 407270 31204
rect 184290 31084 184296 31136
rect 184348 31124 184354 31136
rect 561674 31124 561680 31136
rect 184348 31096 561680 31124
rect 184348 31084 184354 31096
rect 561674 31084 561680 31096
rect 561732 31084 561738 31136
rect 42794 31016 42800 31068
rect 42852 31056 42858 31068
rect 135530 31056 135536 31068
rect 42852 31028 135536 31056
rect 42852 31016 42858 31028
rect 135530 31016 135536 31028
rect 135588 31016 135594 31068
rect 176286 31016 176292 31068
rect 176344 31056 176350 31068
rect 564526 31056 564532 31068
rect 176344 31028 564532 31056
rect 176344 31016 176350 31028
rect 564526 31016 564532 31028
rect 564584 31016 564590 31068
rect 150066 29928 150072 29980
rect 150124 29968 150130 29980
rect 229094 29968 229100 29980
rect 150124 29940 229100 29968
rect 150124 29928 150130 29940
rect 229094 29928 229100 29940
rect 229152 29928 229158 29980
rect 156966 29860 156972 29912
rect 157024 29900 157030 29912
rect 303614 29900 303620 29912
rect 157024 29872 303620 29900
rect 157024 29860 157030 29872
rect 303614 29860 303620 29872
rect 303672 29860 303678 29912
rect 165154 29792 165160 29844
rect 165212 29832 165218 29844
rect 409874 29832 409880 29844
rect 165212 29804 409880 29832
rect 165212 29792 165218 29804
rect 409874 29792 409880 29804
rect 409932 29792 409938 29844
rect 169570 29724 169576 29776
rect 169628 29764 169634 29776
rect 474734 29764 474740 29776
rect 169628 29736 474740 29764
rect 169628 29724 169634 29736
rect 474734 29724 474740 29736
rect 474792 29724 474798 29776
rect 171226 29656 171232 29708
rect 171284 29696 171290 29708
rect 502334 29696 502340 29708
rect 171284 29668 502340 29696
rect 171284 29656 171290 29668
rect 502334 29656 502340 29668
rect 502392 29656 502398 29708
rect 177758 29588 177764 29640
rect 177816 29628 177822 29640
rect 574094 29628 574100 29640
rect 177816 29600 574100 29628
rect 177816 29588 177822 29600
rect 574094 29588 574100 29600
rect 574152 29588 574158 29640
rect 151354 28500 151360 28552
rect 151412 28540 151418 28552
rect 242986 28540 242992 28552
rect 151412 28512 242992 28540
rect 151412 28500 151418 28512
rect 242986 28500 242992 28512
rect 243044 28500 243050 28552
rect 159818 28432 159824 28484
rect 159876 28472 159882 28484
rect 339494 28472 339500 28484
rect 159876 28444 339500 28472
rect 159876 28432 159882 28444
rect 339494 28432 339500 28444
rect 339552 28432 339558 28484
rect 161014 28364 161020 28416
rect 161072 28404 161078 28416
rect 360838 28404 360844 28416
rect 161072 28376 360844 28404
rect 161072 28364 161078 28376
rect 360838 28364 360844 28376
rect 360896 28364 360902 28416
rect 166626 28296 166632 28348
rect 166684 28336 166690 28348
rect 438854 28336 438860 28348
rect 166684 28308 438860 28336
rect 166684 28296 166690 28308
rect 438854 28296 438860 28308
rect 438912 28296 438918 28348
rect 172422 28228 172428 28280
rect 172480 28268 172486 28280
rect 506566 28268 506572 28280
rect 172480 28240 506572 28268
rect 172480 28228 172486 28240
rect 506566 28228 506572 28240
rect 506624 28228 506630 28280
rect 154390 27072 154396 27124
rect 154448 27112 154454 27124
rect 275278 27112 275284 27124
rect 154448 27084 275284 27112
rect 154448 27072 154454 27084
rect 275278 27072 275284 27084
rect 275336 27072 275342 27124
rect 162302 27004 162308 27056
rect 162360 27044 162366 27056
rect 374086 27044 374092 27056
rect 162360 27016 374092 27044
rect 162360 27004 162366 27016
rect 374086 27004 374092 27016
rect 374144 27004 374150 27056
rect 171134 26936 171140 26988
rect 171192 26976 171198 26988
rect 509234 26976 509240 26988
rect 171192 26948 509240 26976
rect 171192 26936 171198 26948
rect 509234 26936 509240 26948
rect 509292 26936 509298 26988
rect 172238 26868 172244 26920
rect 172296 26908 172302 26920
rect 510614 26908 510620 26920
rect 172296 26880 510620 26908
rect 172296 26868 172302 26880
rect 510614 26868 510620 26880
rect 510672 26868 510678 26920
rect 153286 25712 153292 25764
rect 153344 25752 153350 25764
rect 278774 25752 278780 25764
rect 153344 25724 278780 25752
rect 153344 25712 153350 25724
rect 278774 25712 278780 25724
rect 278832 25712 278838 25764
rect 144178 25644 144184 25696
rect 144236 25684 144242 25696
rect 144914 25684 144920 25696
rect 144236 25656 144920 25684
rect 144236 25644 144242 25656
rect 144914 25644 144920 25656
rect 144972 25644 144978 25696
rect 162394 25644 162400 25696
rect 162452 25684 162458 25696
rect 378134 25684 378140 25696
rect 162452 25656 378140 25684
rect 162452 25644 162458 25656
rect 378134 25644 378140 25656
rect 378192 25644 378198 25696
rect 172330 25576 172336 25628
rect 172388 25616 172394 25628
rect 513374 25616 513380 25628
rect 172388 25588 513380 25616
rect 172388 25576 172394 25588
rect 513374 25576 513380 25588
rect 513432 25576 513438 25628
rect 146018 25508 146024 25560
rect 146076 25548 146082 25560
rect 171778 25548 171784 25560
rect 146076 25520 171784 25548
rect 146076 25508 146082 25520
rect 171778 25508 171784 25520
rect 171836 25508 171842 25560
rect 173618 25508 173624 25560
rect 173676 25548 173682 25560
rect 531406 25548 531412 25560
rect 173676 25520 531412 25548
rect 173676 25508 173682 25520
rect 531406 25508 531412 25520
rect 531464 25508 531470 25560
rect 153194 24352 153200 24404
rect 153252 24392 153258 24404
rect 282914 24392 282920 24404
rect 153252 24364 282920 24392
rect 153252 24352 153258 24364
rect 282914 24352 282920 24364
rect 282972 24352 282978 24404
rect 163958 24284 163964 24336
rect 164016 24324 164022 24336
rect 396074 24324 396080 24336
rect 164016 24296 396080 24324
rect 164016 24284 164022 24296
rect 396074 24284 396080 24296
rect 396132 24284 396138 24336
rect 165246 24216 165252 24268
rect 165304 24256 165310 24268
rect 425054 24256 425060 24268
rect 165304 24228 425060 24256
rect 165304 24216 165310 24228
rect 425054 24216 425060 24228
rect 425112 24216 425118 24268
rect 173802 24148 173808 24200
rect 173860 24188 173866 24200
rect 520274 24188 520280 24200
rect 173860 24160 520280 24188
rect 173860 24148 173866 24160
rect 520274 24148 520280 24160
rect 520332 24148 520338 24200
rect 174998 24080 175004 24132
rect 175056 24120 175062 24132
rect 546494 24120 546500 24132
rect 175056 24092 546500 24120
rect 175056 24080 175062 24092
rect 546494 24080 546500 24092
rect 546552 24080 546558 24132
rect 157058 22924 157064 22976
rect 157116 22964 157122 22976
rect 310514 22964 310520 22976
rect 157116 22936 310520 22964
rect 157116 22924 157122 22936
rect 310514 22924 310520 22936
rect 310572 22924 310578 22976
rect 164050 22856 164056 22908
rect 164108 22896 164114 22908
rect 398926 22896 398932 22908
rect 164108 22868 398932 22896
rect 164108 22856 164114 22868
rect 398926 22856 398932 22868
rect 398984 22856 398990 22908
rect 173710 22788 173716 22840
rect 173768 22828 173774 22840
rect 527174 22828 527180 22840
rect 173768 22800 527180 22828
rect 173768 22788 173774 22800
rect 527174 22788 527180 22800
rect 527232 22788 527238 22840
rect 176470 22720 176476 22772
rect 176528 22760 176534 22772
rect 552658 22760 552664 22772
rect 176528 22732 552664 22760
rect 176528 22720 176534 22732
rect 552658 22720 552664 22732
rect 552716 22720 552722 22772
rect 166534 21360 166540 21412
rect 166592 21400 166598 21412
rect 431954 21400 431960 21412
rect 166592 21372 431960 21400
rect 166592 21360 166598 21372
rect 431954 21360 431960 21372
rect 432012 21360 432018 21412
rect 574738 20612 574744 20664
rect 574796 20652 574802 20664
rect 580166 20652 580172 20664
rect 574796 20624 580172 20652
rect 574796 20612 574802 20624
rect 580166 20612 580172 20624
rect 580224 20612 580230 20664
rect 153838 20136 153844 20188
rect 153896 20176 153902 20188
rect 280154 20176 280160 20188
rect 153896 20148 280160 20176
rect 153896 20136 153902 20148
rect 280154 20136 280160 20148
rect 280212 20136 280218 20188
rect 155862 20068 155868 20120
rect 155920 20108 155926 20120
rect 287054 20108 287060 20120
rect 155920 20080 287060 20108
rect 155920 20068 155926 20080
rect 287054 20068 287060 20080
rect 287112 20068 287118 20120
rect 155218 20000 155224 20052
rect 155276 20040 155282 20052
rect 291194 20040 291200 20052
rect 155276 20012 291200 20040
rect 155276 20000 155282 20012
rect 291194 20000 291200 20012
rect 291252 20000 291258 20052
rect 144822 19932 144828 19984
rect 144880 19972 144886 19984
rect 154574 19972 154580 19984
rect 144880 19944 154580 19972
rect 144880 19932 144886 19944
rect 154574 19932 154580 19944
rect 154632 19932 154638 19984
rect 161106 19932 161112 19984
rect 161164 19972 161170 19984
rect 357526 19972 357532 19984
rect 161164 19944 357532 19972
rect 161164 19932 161170 19944
rect 357526 19932 357532 19944
rect 357584 19932 357590 19984
rect 152734 18776 152740 18828
rect 152792 18816 152798 18828
rect 266354 18816 266360 18828
rect 152792 18788 266360 18816
rect 152792 18776 152798 18788
rect 266354 18776 266360 18788
rect 266412 18776 266418 18828
rect 157334 18708 157340 18760
rect 157392 18748 157398 18760
rect 329834 18748 329840 18760
rect 157392 18720 329840 18748
rect 157392 18708 157398 18720
rect 329834 18708 329840 18720
rect 329892 18708 329898 18760
rect 176562 18640 176568 18692
rect 176620 18680 176626 18692
rect 567194 18680 567200 18692
rect 176620 18652 567200 18680
rect 176620 18640 176626 18652
rect 567194 18640 567200 18652
rect 567252 18640 567258 18692
rect 177850 18572 177856 18624
rect 177908 18612 177914 18624
rect 571334 18612 571340 18624
rect 177908 18584 571340 18612
rect 177908 18572 177914 18584
rect 571334 18572 571340 18584
rect 571392 18572 571398 18624
rect 149974 17416 149980 17468
rect 150032 17456 150038 17468
rect 219434 17456 219440 17468
rect 150032 17428 219440 17456
rect 150032 17416 150038 17428
rect 219434 17416 219440 17428
rect 219492 17416 219498 17468
rect 168098 17348 168104 17400
rect 168156 17388 168162 17400
rect 445754 17388 445760 17400
rect 168156 17360 445760 17388
rect 168156 17348 168162 17360
rect 445754 17348 445760 17360
rect 445812 17348 445818 17400
rect 169202 17280 169208 17332
rect 169260 17320 169266 17332
rect 477494 17320 477500 17332
rect 169260 17292 477500 17320
rect 169260 17280 169266 17292
rect 477494 17280 477500 17292
rect 477552 17280 477558 17332
rect 177942 17212 177948 17264
rect 178000 17252 178006 17264
rect 518894 17252 518900 17264
rect 178000 17224 518900 17252
rect 178000 17212 178006 17224
rect 518894 17212 518900 17224
rect 518952 17212 518958 17264
rect 151262 16056 151268 16108
rect 151320 16096 151326 16108
rect 248414 16096 248420 16108
rect 151320 16068 248420 16096
rect 151320 16056 151326 16068
rect 248414 16056 248420 16068
rect 248472 16056 248478 16108
rect 161198 15988 161204 16040
rect 161256 16028 161262 16040
rect 364610 16028 364616 16040
rect 161256 16000 364616 16028
rect 161256 15988 161262 16000
rect 364610 15988 364616 16000
rect 364668 15988 364674 16040
rect 165430 15920 165436 15972
rect 165488 15960 165494 15972
rect 420914 15960 420920 15972
rect 165488 15932 420920 15960
rect 165488 15920 165494 15932
rect 420914 15920 420920 15932
rect 420972 15920 420978 15972
rect 87506 15852 87512 15904
rect 87564 15892 87570 15904
rect 138198 15892 138204 15904
rect 87564 15864 138204 15892
rect 87564 15852 87570 15864
rect 138198 15852 138204 15864
rect 138256 15852 138262 15904
rect 166718 15852 166724 15904
rect 166776 15892 166782 15904
rect 442166 15892 442172 15904
rect 166776 15864 442172 15892
rect 166776 15852 166782 15864
rect 442166 15852 442172 15864
rect 442224 15852 442230 15904
rect 153930 14696 153936 14748
rect 153988 14736 153994 14748
rect 272426 14736 272432 14748
rect 153988 14708 272432 14736
rect 153988 14696 153994 14708
rect 272426 14696 272432 14708
rect 272484 14696 272490 14748
rect 155954 14628 155960 14680
rect 156012 14668 156018 14680
rect 314654 14668 314660 14680
rect 156012 14640 314660 14668
rect 156012 14628 156018 14640
rect 314654 14628 314660 14640
rect 314712 14628 314718 14680
rect 162762 14560 162768 14612
rect 162820 14600 162826 14612
rect 385954 14600 385960 14612
rect 162820 14572 385960 14600
rect 162820 14560 162826 14572
rect 385954 14560 385960 14572
rect 386012 14560 386018 14612
rect 165338 14492 165344 14544
rect 165396 14532 165402 14544
rect 411898 14532 411904 14544
rect 165396 14504 411904 14532
rect 165396 14492 165402 14504
rect 411898 14492 411904 14504
rect 411956 14492 411962 14544
rect 169754 14424 169760 14476
rect 169812 14464 169818 14476
rect 486418 14464 486424 14476
rect 169812 14436 486424 14464
rect 169812 14424 169818 14436
rect 486418 14424 486424 14436
rect 486476 14424 486482 14476
rect 152642 13336 152648 13388
rect 152700 13376 152706 13388
rect 258258 13376 258264 13388
rect 152700 13348 258264 13376
rect 152700 13336 152706 13348
rect 258258 13336 258264 13348
rect 258316 13336 258322 13388
rect 157150 13268 157156 13320
rect 157208 13308 157214 13320
rect 307938 13308 307944 13320
rect 157208 13280 307944 13308
rect 157208 13268 157214 13280
rect 307938 13268 307944 13280
rect 307996 13268 308002 13320
rect 162670 13200 162676 13252
rect 162728 13240 162734 13252
rect 382366 13240 382372 13252
rect 162728 13212 382372 13240
rect 162728 13200 162734 13212
rect 382366 13200 382372 13212
rect 382424 13200 382430 13252
rect 162486 13132 162492 13184
rect 162544 13172 162550 13184
rect 390646 13172 390652 13184
rect 162544 13144 390652 13172
rect 162544 13132 162550 13144
rect 390646 13132 390652 13144
rect 390704 13132 390710 13184
rect 171042 13064 171048 13116
rect 171100 13104 171106 13116
rect 482186 13104 482192 13116
rect 171100 13076 482192 13104
rect 171100 13064 171106 13076
rect 482186 13064 482192 13076
rect 482244 13064 482250 13116
rect 151170 11976 151176 12028
rect 151228 12016 151234 12028
rect 245194 12016 245200 12028
rect 151228 11988 245200 12016
rect 151228 11976 151234 11988
rect 245194 11976 245200 11988
rect 245252 11976 245258 12028
rect 158530 11908 158536 11960
rect 158588 11948 158594 11960
rect 328730 11948 328736 11960
rect 158588 11920 328736 11948
rect 158588 11908 158594 11920
rect 328730 11908 328736 11920
rect 328788 11908 328794 11960
rect 164142 11840 164148 11892
rect 164200 11880 164206 11892
rect 376018 11880 376024 11892
rect 164200 11852 376024 11880
rect 164200 11840 164206 11852
rect 376018 11840 376024 11852
rect 376076 11840 376082 11892
rect 164234 11772 164240 11824
rect 164292 11812 164298 11824
rect 417418 11812 417424 11824
rect 164292 11784 417424 11812
rect 164292 11772 164298 11784
rect 417418 11772 417424 11784
rect 417476 11772 417482 11824
rect 143534 11704 143540 11756
rect 143592 11744 143598 11756
rect 144730 11744 144736 11756
rect 143592 11716 144736 11744
rect 143592 11704 143598 11716
rect 144730 11704 144736 11716
rect 144788 11704 144794 11756
rect 175090 11704 175096 11756
rect 175148 11744 175154 11756
rect 545482 11744 545488 11756
rect 175148 11716 545488 11744
rect 175148 11704 175154 11716
rect 545482 11704 545488 11716
rect 545540 11704 545546 11756
rect 184934 11636 184940 11688
rect 184992 11676 184998 11688
rect 186130 11676 186136 11688
rect 184992 11648 186136 11676
rect 184992 11636 184998 11648
rect 186130 11636 186136 11648
rect 186188 11636 186194 11688
rect 234614 11636 234620 11688
rect 234672 11676 234678 11688
rect 235810 11676 235816 11688
rect 234672 11648 235816 11676
rect 234672 11636 234678 11648
rect 235810 11636 235816 11648
rect 235868 11636 235874 11688
rect 151078 10548 151084 10600
rect 151136 10588 151142 10600
rect 241698 10588 241704 10600
rect 151136 10560 241704 10588
rect 151136 10548 151142 10560
rect 241698 10548 241704 10560
rect 241756 10548 241762 10600
rect 158622 10480 158628 10532
rect 158680 10520 158686 10532
rect 336274 10520 336280 10532
rect 158680 10492 336280 10520
rect 158680 10480 158686 10492
rect 336274 10480 336280 10492
rect 336332 10480 336338 10532
rect 162578 10412 162584 10464
rect 162636 10452 162642 10464
rect 386690 10452 386696 10464
rect 162636 10424 386696 10452
rect 162636 10412 162642 10424
rect 386690 10412 386696 10424
rect 386748 10412 386754 10464
rect 166810 10344 166816 10396
rect 166868 10384 166874 10396
rect 432046 10384 432052 10396
rect 166868 10356 432052 10384
rect 166868 10344 166874 10356
rect 432046 10344 432052 10356
rect 432104 10344 432110 10396
rect 175182 10276 175188 10328
rect 175240 10316 175246 10328
rect 548426 10316 548432 10328
rect 175240 10288 548432 10316
rect 175240 10276 175246 10288
rect 548426 10276 548432 10288
rect 548484 10276 548490 10328
rect 157242 9052 157248 9104
rect 157300 9092 157306 9104
rect 316218 9092 316224 9104
rect 157300 9064 316224 9092
rect 157300 9052 157306 9064
rect 316218 9052 316224 9064
rect 316276 9052 316282 9104
rect 165522 8984 165528 9036
rect 165580 9024 165586 9036
rect 414290 9024 414296 9036
rect 165580 8996 414296 9024
rect 165580 8984 165586 8996
rect 414290 8984 414296 8996
rect 414348 8984 414354 9036
rect 52546 8916 52552 8968
rect 52604 8956 52610 8968
rect 135346 8956 135352 8968
rect 52604 8928 135352 8956
rect 52604 8916 52610 8928
rect 135346 8916 135352 8928
rect 135404 8916 135410 8968
rect 175366 8916 175372 8968
rect 175424 8956 175430 8968
rect 556154 8956 556160 8968
rect 175424 8928 556160 8956
rect 175424 8916 175430 8928
rect 556154 8916 556160 8928
rect 556212 8916 556218 8968
rect 142798 8236 142804 8288
rect 142856 8276 142862 8288
rect 143534 8276 143540 8288
rect 142856 8248 143540 8276
rect 142856 8236 142862 8248
rect 143534 8236 143540 8248
rect 143592 8236 143598 8288
rect 149882 7828 149888 7880
rect 149940 7868 149946 7880
rect 227530 7868 227536 7880
rect 149940 7840 227536 7868
rect 149940 7828 149946 7840
rect 227530 7828 227536 7840
rect 227588 7828 227594 7880
rect 159910 7760 159916 7812
rect 159968 7800 159974 7812
rect 343358 7800 343364 7812
rect 159968 7772 343364 7800
rect 159968 7760 159974 7772
rect 343358 7760 343364 7772
rect 343416 7760 343422 7812
rect 161290 7692 161296 7744
rect 161348 7732 161354 7744
rect 365806 7732 365812 7744
rect 161348 7704 365812 7732
rect 161348 7692 161354 7704
rect 365806 7692 365812 7704
rect 365864 7692 365870 7744
rect 166902 7624 166908 7676
rect 166960 7664 166966 7676
rect 435542 7664 435548 7676
rect 166960 7636 435548 7664
rect 166960 7624 166966 7636
rect 435542 7624 435548 7636
rect 435600 7624 435606 7676
rect 25314 7556 25320 7608
rect 25372 7596 25378 7608
rect 133874 7596 133880 7608
rect 25372 7568 133880 7596
rect 25372 7556 25378 7568
rect 133874 7556 133880 7568
rect 133932 7556 133938 7608
rect 173986 7556 173992 7608
rect 174044 7596 174050 7608
rect 538398 7596 538404 7608
rect 174044 7568 538404 7596
rect 174044 7556 174050 7568
rect 538398 7556 538404 7568
rect 538456 7556 538462 7608
rect 152550 6536 152556 6588
rect 152608 6576 152614 6588
rect 259546 6576 259552 6588
rect 152608 6548 259552 6576
rect 152608 6536 152614 6548
rect 259546 6536 259552 6548
rect 259604 6536 259610 6588
rect 160002 6468 160008 6520
rect 160060 6508 160066 6520
rect 350442 6508 350448 6520
rect 160060 6480 350448 6508
rect 160060 6468 160066 6480
rect 350442 6468 350448 6480
rect 350500 6468 350506 6520
rect 179138 6400 179144 6452
rect 179196 6440 179202 6452
rect 443822 6440 443828 6452
rect 179196 6412 443828 6440
rect 179196 6400 179202 6412
rect 443822 6400 443828 6412
rect 443880 6400 443886 6452
rect 180610 6332 180616 6384
rect 180668 6372 180674 6384
rect 450906 6372 450912 6384
rect 180668 6344 450912 6372
rect 180668 6332 180674 6344
rect 450906 6332 450912 6344
rect 450964 6332 450970 6384
rect 168190 6264 168196 6316
rect 168248 6304 168254 6316
rect 453298 6304 453304 6316
rect 168248 6276 453304 6304
rect 168248 6264 168254 6276
rect 453298 6264 453304 6276
rect 453356 6264 453362 6316
rect 176194 6196 176200 6248
rect 176252 6236 176258 6248
rect 563238 6236 563244 6248
rect 176252 6208 563244 6236
rect 176252 6196 176258 6208
rect 563238 6196 563244 6208
rect 563296 6196 563302 6248
rect 103330 6128 103336 6180
rect 103388 6168 103394 6180
rect 139762 6168 139768 6180
rect 103388 6140 139768 6168
rect 103388 6128 103394 6140
rect 139762 6128 139768 6140
rect 139820 6128 139826 6180
rect 182082 6128 182088 6180
rect 182140 6168 182146 6180
rect 583386 6168 583392 6180
rect 182140 6140 583392 6168
rect 182140 6128 182146 6140
rect 583386 6128 583392 6140
rect 583444 6128 583450 6180
rect 154482 4972 154488 5024
rect 154540 5012 154546 5024
rect 273622 5012 273628 5024
rect 154540 4984 273628 5012
rect 154540 4972 154546 4984
rect 273622 4972 273628 4984
rect 273680 4972 273686 5024
rect 161382 4904 161388 4956
rect 161440 4944 161446 4956
rect 371694 4944 371700 4956
rect 161440 4916 371700 4944
rect 161440 4904 161446 4916
rect 371694 4904 371700 4916
rect 371752 4904 371758 4956
rect 168282 4836 168288 4888
rect 168340 4876 168346 4888
rect 456886 4876 456892 4888
rect 168340 4848 456892 4876
rect 168340 4836 168346 4848
rect 456886 4836 456892 4848
rect 456944 4836 456950 4888
rect 6454 4768 6460 4820
rect 6512 4808 6518 4820
rect 132678 4808 132684 4820
rect 6512 4780 132684 4808
rect 6512 4768 6518 4780
rect 132678 4768 132684 4780
rect 132736 4768 132742 4820
rect 173894 4768 173900 4820
rect 173952 4808 173958 4820
rect 541986 4808 541992 4820
rect 173952 4780 541992 4808
rect 173952 4768 173958 4780
rect 541986 4768 541992 4780
rect 542044 4768 542050 4820
rect 231044 4168 231256 4196
rect 566 4088 572 4140
rect 624 4128 630 4140
rect 7558 4128 7564 4140
rect 624 4100 7564 4128
rect 624 4088 630 4100
rect 7558 4088 7564 4100
rect 7616 4088 7622 4140
rect 73798 4088 73804 4140
rect 73856 4128 73862 4140
rect 75178 4128 75184 4140
rect 73856 4100 75184 4128
rect 73856 4088 73862 4100
rect 75178 4088 75184 4100
rect 75236 4088 75242 4140
rect 112806 4088 112812 4140
rect 112864 4128 112870 4140
rect 113818 4128 113824 4140
rect 112864 4100 113824 4128
rect 112864 4088 112870 4100
rect 113818 4088 113824 4100
rect 113876 4088 113882 4140
rect 141234 4088 141240 4140
rect 141292 4128 141298 4140
rect 142338 4128 142344 4140
rect 141292 4100 142344 4128
rect 141292 4088 141298 4100
rect 142338 4088 142344 4100
rect 142396 4088 142402 4140
rect 149698 4088 149704 4140
rect 149756 4128 149762 4140
rect 153010 4128 153016 4140
rect 149756 4100 153016 4128
rect 149756 4088 149762 4100
rect 153010 4088 153016 4100
rect 153068 4088 153074 4140
rect 189810 4088 189816 4140
rect 189868 4128 189874 4140
rect 203886 4128 203892 4140
rect 189868 4100 203892 4128
rect 189868 4088 189874 4100
rect 203886 4088 203892 4100
rect 203944 4088 203950 4140
rect 211798 4088 211804 4140
rect 211856 4128 211862 4140
rect 217318 4128 217324 4140
rect 211856 4100 217324 4128
rect 211856 4088 211862 4100
rect 217318 4088 217324 4100
rect 217376 4088 217382 4140
rect 229738 4088 229744 4140
rect 229796 4128 229802 4140
rect 230934 4128 230940 4140
rect 229796 4100 230940 4128
rect 229796 4088 229802 4100
rect 230934 4088 230940 4100
rect 230992 4088 230998 4140
rect 181438 4020 181444 4072
rect 181496 4060 181502 4072
rect 190822 4060 190828 4072
rect 181496 4032 190828 4060
rect 181496 4020 181502 4032
rect 190822 4020 190828 4032
rect 190880 4020 190886 4072
rect 193858 4020 193864 4072
rect 193916 4060 193922 4072
rect 195606 4060 195612 4072
rect 193916 4032 195612 4060
rect 193916 4020 193922 4032
rect 195606 4020 195612 4032
rect 195664 4020 195670 4072
rect 195698 4020 195704 4072
rect 195756 4060 195762 4072
rect 216490 4060 216496 4072
rect 195756 4032 216496 4060
rect 195756 4020 195762 4032
rect 216490 4020 216496 4032
rect 216548 4020 216554 4072
rect 216674 4020 216680 4072
rect 216732 4060 216738 4072
rect 231044 4060 231072 4168
rect 231228 4128 231256 4168
rect 247586 4128 247592 4140
rect 231228 4100 247592 4128
rect 247586 4088 247592 4100
rect 247644 4088 247650 4140
rect 247678 4088 247684 4140
rect 247736 4128 247742 4140
rect 254670 4128 254676 4140
rect 247736 4100 254676 4128
rect 247736 4088 247742 4100
rect 254670 4088 254676 4100
rect 254728 4088 254734 4140
rect 315298 4088 315304 4140
rect 315356 4128 315362 4140
rect 317322 4128 317328 4140
rect 315356 4100 317328 4128
rect 315356 4088 315362 4100
rect 317322 4088 317328 4100
rect 317380 4088 317386 4140
rect 323578 4088 323584 4140
rect 323636 4128 323642 4140
rect 326798 4128 326804 4140
rect 323636 4100 326804 4128
rect 323636 4088 323642 4100
rect 326798 4088 326804 4100
rect 326856 4088 326862 4140
rect 450538 4088 450544 4140
rect 450596 4128 450602 4140
rect 452102 4128 452108 4140
rect 450596 4100 452108 4128
rect 450596 4088 450602 4100
rect 452102 4088 452108 4100
rect 452160 4088 452166 4140
rect 486510 4088 486516 4140
rect 486568 4128 486574 4140
rect 489914 4128 489920 4140
rect 486568 4100 489920 4128
rect 486568 4088 486574 4100
rect 489914 4088 489920 4100
rect 489972 4088 489978 4140
rect 527910 4088 527916 4140
rect 527968 4128 527974 4140
rect 529014 4128 529020 4140
rect 527968 4100 529020 4128
rect 527968 4088 527974 4100
rect 529014 4088 529020 4100
rect 529072 4088 529078 4140
rect 216732 4032 231072 4060
rect 216732 4020 216738 4032
rect 251174 4020 251180 4072
rect 251232 4060 251238 4072
rect 252370 4060 252376 4072
rect 251232 4032 252376 4060
rect 251232 4020 251238 4032
rect 252370 4020 252376 4032
rect 252428 4020 252434 4072
rect 181530 3952 181536 4004
rect 181588 3992 181594 4004
rect 212166 3992 212172 4004
rect 181588 3964 212172 3992
rect 181588 3952 181594 3964
rect 212166 3952 212172 3964
rect 212224 3952 212230 4004
rect 217318 3952 217324 4004
rect 217376 3992 217382 4004
rect 231026 3992 231032 4004
rect 217376 3964 231032 3992
rect 217376 3952 217382 3964
rect 231026 3952 231032 3964
rect 231084 3952 231090 4004
rect 231118 3952 231124 4004
rect 231176 3992 231182 4004
rect 298462 3992 298468 4004
rect 231176 3964 298468 3992
rect 231176 3952 231182 3964
rect 298462 3952 298468 3964
rect 298520 3952 298526 4004
rect 299566 3952 299572 4004
rect 299624 3992 299630 4004
rect 300762 3992 300768 4004
rect 299624 3964 300768 3992
rect 299624 3952 299630 3964
rect 300762 3952 300768 3964
rect 300820 3952 300826 4004
rect 311158 3952 311164 4004
rect 311216 3992 311222 4004
rect 312630 3992 312636 4004
rect 311216 3964 312636 3992
rect 311216 3952 311222 3964
rect 312630 3952 312636 3964
rect 312688 3952 312694 4004
rect 360838 3952 360844 4004
rect 360896 3992 360902 4004
rect 362310 3992 362316 4004
rect 360896 3964 362316 3992
rect 360896 3952 360902 3964
rect 362310 3952 362316 3964
rect 362368 3952 362374 4004
rect 127066 3924 127072 3936
rect 122806 3896 127072 3924
rect 122282 3680 122288 3732
rect 122340 3720 122346 3732
rect 122806 3720 122834 3896
rect 127066 3884 127072 3896
rect 127124 3884 127130 3936
rect 152458 3884 152464 3936
rect 152516 3924 152522 3936
rect 161382 3924 161388 3936
rect 152516 3896 161388 3924
rect 152516 3884 152522 3896
rect 161382 3884 161388 3896
rect 161440 3884 161446 3936
rect 178678 3884 178684 3936
rect 178736 3924 178742 3936
rect 401318 3924 401324 3936
rect 178736 3896 401324 3924
rect 178736 3884 178742 3896
rect 401318 3884 401324 3896
rect 401376 3884 401382 3936
rect 131298 3856 131304 3868
rect 122340 3692 122834 3720
rect 123220 3828 131304 3856
rect 122340 3680 122346 3692
rect 65518 3612 65524 3664
rect 65576 3652 65582 3664
rect 65576 3624 74534 3652
rect 65576 3612 65582 3624
rect 17034 3544 17040 3596
rect 17092 3584 17098 3596
rect 18598 3584 18604 3596
rect 17092 3556 18604 3584
rect 17092 3544 17098 3556
rect 18598 3544 18604 3556
rect 18656 3544 18662 3596
rect 19426 3544 19432 3596
rect 19484 3584 19490 3596
rect 21358 3584 21364 3596
rect 19484 3556 21364 3584
rect 19484 3544 19490 3556
rect 21358 3544 21364 3556
rect 21416 3544 21422 3596
rect 27614 3544 27620 3596
rect 27672 3584 27678 3596
rect 28534 3584 28540 3596
rect 27672 3556 28540 3584
rect 27672 3544 27678 3556
rect 28534 3544 28540 3556
rect 28592 3544 28598 3596
rect 51350 3544 51356 3596
rect 51408 3584 51414 3596
rect 54478 3584 54484 3596
rect 51408 3556 54484 3584
rect 51408 3544 51414 3556
rect 54478 3544 54484 3556
rect 54536 3544 54542 3596
rect 56042 3544 56048 3596
rect 56100 3584 56106 3596
rect 57238 3584 57244 3596
rect 56100 3556 57244 3584
rect 56100 3544 56106 3556
rect 57238 3544 57244 3556
rect 57296 3544 57302 3596
rect 60734 3544 60740 3596
rect 60792 3584 60798 3596
rect 61654 3584 61660 3596
rect 60792 3556 61660 3584
rect 60792 3544 60798 3556
rect 61654 3544 61660 3556
rect 61712 3544 61718 3596
rect 69106 3544 69112 3596
rect 69164 3584 69170 3596
rect 71038 3584 71044 3596
rect 69164 3556 71044 3584
rect 69164 3544 69170 3556
rect 71038 3544 71044 3556
rect 71096 3544 71102 3596
rect 74506 3584 74534 3624
rect 83274 3612 83280 3664
rect 83332 3652 83338 3664
rect 123220 3652 123248 3828
rect 131298 3816 131304 3828
rect 131356 3816 131362 3868
rect 132954 3816 132960 3868
rect 133012 3856 133018 3868
rect 140038 3856 140044 3868
rect 133012 3828 140044 3856
rect 133012 3816 133018 3828
rect 140038 3816 140044 3828
rect 140096 3816 140102 3868
rect 146938 3816 146944 3868
rect 146996 3856 147002 3868
rect 149606 3856 149612 3868
rect 146996 3828 149612 3856
rect 146996 3816 147002 3828
rect 149606 3816 149612 3828
rect 149664 3816 149670 3868
rect 149790 3816 149796 3868
rect 149848 3856 149854 3868
rect 163682 3856 163688 3868
rect 149848 3828 163688 3856
rect 149848 3816 149854 3828
rect 163682 3816 163688 3828
rect 163740 3816 163746 3868
rect 170398 3816 170404 3868
rect 170456 3856 170462 3868
rect 173158 3856 173164 3868
rect 170456 3828 173164 3856
rect 170456 3816 170462 3828
rect 173158 3816 173164 3828
rect 173216 3816 173222 3868
rect 178770 3816 178776 3868
rect 178828 3856 178834 3868
rect 408402 3856 408408 3868
rect 178828 3828 408408 3856
rect 178828 3816 178834 3828
rect 408402 3816 408408 3828
rect 408460 3816 408466 3868
rect 129826 3788 129832 3800
rect 83332 3624 123248 3652
rect 123312 3760 129832 3788
rect 83332 3612 83338 3624
rect 123312 3584 123340 3760
rect 129826 3748 129832 3760
rect 129884 3748 129890 3800
rect 131022 3748 131028 3800
rect 131080 3788 131086 3800
rect 150618 3788 150624 3800
rect 131080 3760 150624 3788
rect 131080 3748 131086 3760
rect 150618 3748 150624 3760
rect 150676 3748 150682 3800
rect 160094 3748 160100 3800
rect 160152 3788 160158 3800
rect 161290 3788 161296 3800
rect 160152 3760 161296 3788
rect 160152 3748 160158 3760
rect 161290 3748 161296 3760
rect 161348 3748 161354 3800
rect 161382 3748 161388 3800
rect 161440 3788 161446 3800
rect 171962 3788 171968 3800
rect 161440 3760 171968 3788
rect 161440 3748 161446 3760
rect 171962 3748 171968 3760
rect 172020 3748 172026 3800
rect 179322 3748 179328 3800
rect 179380 3788 179386 3800
rect 429654 3788 429660 3800
rect 179380 3760 429660 3788
rect 179380 3748 179386 3760
rect 429654 3748 429660 3760
rect 429712 3748 429718 3800
rect 74506 3556 123340 3584
rect 123404 3692 129964 3720
rect 15930 3476 15936 3528
rect 15988 3516 15994 3528
rect 123404 3516 123432 3692
rect 129936 3652 129964 3692
rect 130838 3680 130844 3732
rect 130896 3720 130902 3732
rect 162486 3720 162492 3732
rect 130896 3692 162492 3720
rect 130896 3680 130902 3692
rect 162486 3680 162492 3692
rect 162544 3680 162550 3732
rect 170766 3720 170772 3732
rect 163332 3692 170772 3720
rect 131390 3652 131396 3664
rect 129936 3624 131396 3652
rect 131390 3612 131396 3624
rect 131448 3612 131454 3664
rect 137646 3612 137652 3664
rect 137704 3652 137710 3664
rect 138658 3652 138664 3664
rect 137704 3624 138664 3652
rect 137704 3612 137710 3624
rect 138658 3612 138664 3624
rect 138716 3612 138722 3664
rect 147030 3612 147036 3664
rect 147088 3652 147094 3664
rect 149514 3652 149520 3664
rect 147088 3624 149520 3652
rect 147088 3612 147094 3624
rect 149514 3612 149520 3624
rect 149572 3612 149578 3664
rect 149606 3612 149612 3664
rect 149664 3652 149670 3664
rect 163332 3652 163360 3692
rect 170766 3680 170772 3692
rect 170824 3680 170830 3732
rect 179230 3680 179236 3732
rect 179288 3720 179294 3732
rect 436738 3720 436744 3732
rect 179288 3692 436744 3720
rect 179288 3680 179294 3692
rect 436738 3680 436744 3692
rect 436796 3680 436802 3732
rect 442258 3680 442264 3732
rect 442316 3720 442322 3732
rect 497090 3720 497096 3732
rect 442316 3692 497096 3720
rect 442316 3680 442322 3692
rect 497090 3680 497096 3692
rect 497148 3680 497154 3732
rect 166074 3652 166080 3664
rect 149664 3624 163360 3652
rect 163424 3624 166080 3652
rect 149664 3612 149670 3624
rect 125870 3544 125876 3596
rect 125928 3584 125934 3596
rect 129918 3584 129924 3596
rect 125928 3556 129924 3584
rect 125928 3544 125934 3556
rect 129918 3544 129924 3556
rect 129976 3544 129982 3596
rect 130930 3544 130936 3596
rect 130988 3584 130994 3596
rect 163424 3584 163452 3624
rect 166074 3612 166080 3624
rect 166132 3612 166138 3664
rect 179046 3612 179052 3664
rect 179104 3652 179110 3664
rect 447410 3652 447416 3664
rect 179104 3624 447416 3652
rect 179104 3612 179110 3624
rect 447410 3612 447416 3624
rect 447468 3612 447474 3664
rect 130988 3556 163452 3584
rect 130988 3544 130994 3556
rect 163498 3544 163504 3596
rect 163556 3584 163562 3596
rect 164878 3584 164884 3596
rect 163556 3556 164884 3584
rect 163556 3544 163562 3556
rect 164878 3544 164884 3556
rect 164936 3544 164942 3596
rect 168374 3544 168380 3596
rect 168432 3584 168438 3596
rect 169570 3584 169576 3596
rect 168432 3556 169576 3584
rect 168432 3544 168438 3556
rect 169570 3544 169576 3556
rect 169628 3544 169634 3596
rect 186222 3544 186228 3596
rect 186280 3584 186286 3596
rect 468294 3584 468300 3596
rect 186280 3556 468300 3584
rect 186280 3544 186286 3556
rect 468294 3544 468300 3556
rect 468352 3544 468358 3596
rect 468478 3544 468484 3596
rect 468536 3584 468542 3596
rect 469858 3584 469864 3596
rect 468536 3556 469864 3584
rect 468536 3544 468542 3556
rect 469858 3544 469864 3556
rect 469916 3544 469922 3596
rect 470566 3556 478184 3584
rect 15988 3488 123432 3516
rect 15988 3476 15994 3488
rect 123478 3476 123484 3528
rect 123536 3516 123542 3528
rect 124858 3516 124864 3528
rect 123536 3488 124864 3516
rect 123536 3476 123542 3488
rect 124858 3476 124864 3488
rect 124916 3476 124922 3528
rect 128170 3476 128176 3528
rect 128228 3516 128234 3528
rect 128998 3516 129004 3528
rect 128228 3488 129004 3516
rect 128228 3476 128234 3488
rect 128998 3476 129004 3488
rect 129056 3476 129062 3528
rect 140038 3476 140044 3528
rect 140096 3516 140102 3528
rect 141510 3516 141516 3528
rect 140096 3488 141516 3516
rect 140096 3476 140102 3488
rect 141510 3476 141516 3488
rect 141568 3476 141574 3528
rect 147214 3476 147220 3528
rect 147272 3516 147278 3528
rect 175458 3516 175464 3528
rect 147272 3488 175464 3516
rect 147272 3476 147278 3488
rect 175458 3476 175464 3488
rect 175516 3476 175522 3528
rect 180702 3476 180708 3528
rect 180760 3516 180766 3528
rect 470566 3516 470594 3556
rect 180760 3488 470594 3516
rect 180760 3476 180766 3488
rect 472618 3476 472624 3528
rect 472676 3516 472682 3528
rect 473446 3516 473452 3528
rect 472676 3488 473452 3516
rect 472676 3476 472682 3488
rect 473446 3476 473452 3488
rect 473504 3476 473510 3528
rect 478156 3516 478184 3556
rect 478230 3544 478236 3596
rect 478288 3584 478294 3596
rect 498194 3584 498200 3596
rect 478288 3556 498200 3584
rect 478288 3544 478294 3556
rect 498194 3544 498200 3556
rect 498252 3544 498258 3596
rect 516778 3544 516784 3596
rect 516836 3584 516842 3596
rect 518342 3584 518348 3596
rect 516836 3556 518348 3584
rect 516836 3544 516842 3556
rect 518342 3544 518348 3556
rect 518400 3544 518406 3596
rect 479334 3516 479340 3528
rect 478156 3488 479340 3516
rect 479334 3476 479340 3488
rect 479392 3476 479398 3528
rect 482278 3476 482284 3528
rect 482336 3516 482342 3528
rect 507670 3516 507676 3528
rect 482336 3488 507676 3516
rect 482336 3476 482342 3488
rect 507670 3476 507676 3488
rect 507728 3476 507734 3528
rect 526438 3476 526444 3528
rect 526496 3516 526502 3528
rect 533706 3516 533712 3528
rect 526496 3488 533712 3516
rect 526496 3476 526502 3488
rect 533706 3476 533712 3488
rect 533764 3476 533770 3528
rect 538858 3476 538864 3528
rect 538916 3516 538922 3528
rect 539594 3516 539600 3528
rect 538916 3488 539600 3516
rect 538916 3476 538922 3488
rect 539594 3476 539600 3488
rect 539652 3476 539658 3528
rect 540238 3476 540244 3528
rect 540296 3516 540302 3528
rect 547874 3516 547880 3528
rect 540296 3488 547880 3516
rect 540296 3476 540302 3488
rect 547874 3476 547880 3488
rect 547932 3476 547938 3528
rect 552750 3476 552756 3528
rect 552808 3516 552814 3528
rect 560846 3516 560852 3528
rect 552808 3488 560852 3516
rect 552808 3476 552814 3488
rect 560846 3476 560852 3488
rect 560904 3476 560910 3528
rect 563698 3476 563704 3528
rect 563756 3516 563762 3528
rect 565630 3516 565636 3528
rect 563756 3488 565636 3516
rect 563756 3476 563762 3488
rect 565630 3476 565636 3488
rect 565688 3476 565694 3528
rect 567838 3476 567844 3528
rect 567896 3516 567902 3528
rect 569126 3516 569132 3528
rect 567896 3488 569132 3516
rect 567896 3476 567902 3488
rect 569126 3476 569132 3488
rect 569184 3476 569190 3528
rect 1670 3408 1676 3460
rect 1728 3448 1734 3460
rect 8938 3448 8944 3460
rect 1728 3420 8944 3448
rect 1728 3408 1734 3420
rect 8938 3408 8944 3420
rect 8996 3408 9002 3460
rect 11146 3408 11152 3460
rect 11204 3448 11210 3460
rect 11204 3420 122834 3448
rect 11204 3408 11210 3420
rect 91554 3340 91560 3392
rect 91612 3380 91618 3392
rect 93118 3380 93124 3392
rect 91612 3352 93124 3380
rect 91612 3340 91618 3352
rect 93118 3340 93124 3352
rect 93176 3340 93182 3392
rect 101030 3340 101036 3392
rect 101088 3380 101094 3392
rect 102870 3380 102876 3392
rect 101088 3352 102876 3380
rect 101088 3340 101094 3352
rect 102870 3340 102876 3352
rect 102928 3340 102934 3392
rect 105722 3340 105728 3392
rect 105780 3380 105786 3392
rect 106918 3380 106924 3392
rect 105780 3352 106924 3380
rect 105780 3340 105786 3352
rect 106918 3340 106924 3352
rect 106976 3340 106982 3392
rect 111610 3340 111616 3392
rect 111668 3380 111674 3392
rect 112438 3380 112444 3392
rect 111668 3352 112444 3380
rect 111668 3340 111674 3352
rect 112438 3340 112444 3352
rect 112496 3340 112502 3392
rect 120074 3340 120080 3392
rect 120132 3380 120138 3392
rect 120718 3380 120724 3392
rect 120132 3352 120724 3380
rect 120132 3340 120138 3352
rect 120718 3340 120724 3352
rect 120776 3340 120782 3392
rect 122806 3380 122834 3420
rect 148318 3408 148324 3460
rect 148376 3448 148382 3460
rect 176654 3448 176660 3460
rect 148376 3420 176660 3448
rect 148376 3408 148382 3420
rect 176654 3408 176660 3420
rect 176712 3408 176718 3460
rect 180518 3408 180524 3460
rect 180576 3448 180582 3460
rect 487614 3448 487620 3460
rect 180576 3420 487620 3448
rect 180576 3408 180582 3420
rect 487614 3408 487620 3420
rect 487672 3408 487678 3460
rect 498838 3408 498844 3460
rect 498896 3448 498902 3460
rect 540790 3448 540796 3460
rect 498896 3420 540796 3448
rect 498896 3408 498902 3420
rect 540790 3408 540796 3420
rect 540848 3408 540854 3460
rect 545758 3408 545764 3460
rect 545816 3448 545822 3460
rect 554958 3448 554964 3460
rect 545816 3420 554964 3448
rect 545816 3408 545822 3420
rect 554958 3408 554964 3420
rect 555016 3408 555022 3460
rect 560938 3408 560944 3460
rect 560996 3448 561002 3460
rect 573910 3448 573916 3460
rect 560996 3420 573916 3448
rect 560996 3408 561002 3420
rect 573910 3408 573916 3420
rect 573968 3408 573974 3460
rect 131114 3380 131120 3392
rect 122806 3352 131120 3380
rect 131114 3340 131120 3352
rect 131172 3340 131178 3392
rect 147306 3340 147312 3392
rect 147364 3380 147370 3392
rect 151814 3380 151820 3392
rect 147364 3352 151820 3380
rect 147364 3340 147370 3352
rect 151814 3340 151820 3352
rect 151872 3340 151878 3392
rect 182818 3340 182824 3392
rect 182876 3380 182882 3392
rect 193214 3380 193220 3392
rect 182876 3352 193220 3380
rect 182876 3340 182882 3352
rect 193214 3340 193220 3352
rect 193272 3340 193278 3392
rect 210418 3340 210424 3392
rect 210476 3380 210482 3392
rect 218054 3380 218060 3392
rect 210476 3352 218060 3380
rect 210476 3340 210482 3352
rect 218054 3340 218060 3352
rect 218112 3340 218118 3392
rect 225598 3340 225604 3392
rect 225656 3380 225662 3392
rect 226334 3380 226340 3392
rect 225656 3352 226340 3380
rect 225656 3340 225662 3352
rect 226334 3340 226340 3352
rect 226392 3340 226398 3392
rect 239398 3340 239404 3392
rect 239456 3380 239462 3392
rect 240502 3380 240508 3392
rect 239456 3352 240508 3380
rect 239456 3340 239462 3352
rect 240502 3340 240508 3352
rect 240560 3340 240566 3392
rect 242158 3340 242164 3392
rect 242216 3380 242222 3392
rect 242894 3380 242900 3392
rect 242216 3352 242900 3380
rect 242216 3340 242222 3352
rect 242894 3340 242900 3352
rect 242952 3340 242958 3392
rect 259454 3340 259460 3392
rect 259512 3380 259518 3392
rect 260650 3380 260656 3392
rect 259512 3352 260656 3380
rect 259512 3340 259518 3352
rect 260650 3340 260656 3352
rect 260708 3340 260714 3392
rect 261478 3340 261484 3392
rect 261536 3380 261542 3392
rect 262950 3380 262956 3392
rect 261536 3352 262956 3380
rect 261536 3340 261542 3352
rect 262950 3340 262956 3352
rect 263008 3340 263014 3392
rect 275278 3340 275284 3392
rect 275336 3380 275342 3392
rect 276014 3380 276020 3392
rect 275336 3352 276020 3380
rect 275336 3340 275342 3352
rect 276014 3340 276020 3352
rect 276072 3340 276078 3392
rect 307018 3340 307024 3392
rect 307076 3380 307082 3392
rect 309042 3380 309048 3392
rect 307076 3352 309048 3380
rect 307076 3340 307082 3352
rect 309042 3340 309048 3352
rect 309100 3340 309106 3392
rect 324406 3340 324412 3392
rect 324464 3380 324470 3392
rect 325602 3380 325608 3392
rect 324464 3352 325608 3380
rect 324464 3340 324470 3352
rect 325602 3340 325608 3352
rect 325660 3340 325666 3392
rect 332594 3340 332600 3392
rect 332652 3380 332658 3392
rect 333882 3380 333888 3392
rect 332652 3352 333888 3380
rect 332652 3340 332658 3352
rect 333882 3340 333888 3352
rect 333940 3340 333946 3392
rect 340874 3340 340880 3392
rect 340932 3380 340938 3392
rect 342162 3380 342168 3392
rect 340932 3352 342168 3380
rect 340932 3340 340938 3352
rect 342162 3340 342168 3352
rect 342220 3340 342226 3392
rect 342898 3340 342904 3392
rect 342956 3380 342962 3392
rect 344554 3380 344560 3392
rect 342956 3352 344560 3380
rect 342956 3340 342962 3352
rect 344554 3340 344560 3352
rect 344612 3340 344618 3392
rect 357526 3340 357532 3392
rect 357584 3380 357590 3392
rect 358722 3380 358728 3392
rect 357584 3352 358728 3380
rect 357584 3340 357590 3352
rect 358722 3340 358728 3352
rect 358780 3340 358786 3392
rect 364978 3340 364984 3392
rect 365036 3380 365042 3392
rect 367002 3380 367008 3392
rect 365036 3352 367008 3380
rect 365036 3340 365042 3352
rect 367002 3340 367008 3352
rect 367060 3340 367066 3392
rect 374086 3340 374092 3392
rect 374144 3380 374150 3392
rect 375282 3380 375288 3392
rect 374144 3352 375288 3380
rect 374144 3340 374150 3352
rect 375282 3340 375288 3352
rect 375340 3340 375346 3392
rect 378778 3340 378784 3392
rect 378836 3380 378842 3392
rect 379974 3380 379980 3392
rect 378836 3352 379980 3380
rect 378836 3340 378842 3352
rect 379974 3340 379980 3352
rect 380032 3340 380038 3392
rect 382274 3340 382280 3392
rect 382332 3380 382338 3392
rect 383562 3380 383568 3392
rect 382332 3352 383568 3380
rect 382332 3340 382338 3352
rect 383562 3340 383568 3352
rect 383620 3340 383626 3392
rect 398926 3340 398932 3392
rect 398984 3380 398990 3392
rect 400122 3380 400128 3392
rect 398984 3352 400128 3380
rect 398984 3340 398990 3352
rect 400122 3340 400128 3352
rect 400180 3340 400186 3392
rect 400858 3340 400864 3392
rect 400916 3380 400922 3392
rect 402514 3380 402520 3392
rect 400916 3352 402520 3380
rect 400916 3340 400922 3352
rect 402514 3340 402520 3352
rect 402572 3340 402578 3392
rect 414658 3340 414664 3392
rect 414716 3380 414722 3392
rect 416682 3380 416688 3392
rect 414716 3352 416688 3380
rect 414716 3340 414722 3352
rect 416682 3340 416688 3352
rect 416740 3340 416746 3392
rect 418798 3340 418804 3392
rect 418856 3380 418862 3392
rect 420178 3380 420184 3392
rect 418856 3352 420184 3380
rect 418856 3340 418862 3352
rect 420178 3340 420184 3352
rect 420236 3340 420242 3392
rect 422938 3340 422944 3392
rect 422996 3380 423002 3392
rect 424962 3380 424968 3392
rect 422996 3352 424968 3380
rect 422996 3340 423002 3352
rect 424962 3340 424968 3352
rect 425020 3340 425026 3392
rect 432598 3340 432604 3392
rect 432656 3380 432662 3392
rect 434438 3380 434444 3392
rect 432656 3352 434444 3380
rect 432656 3340 432662 3352
rect 434438 3340 434444 3352
rect 434496 3340 434502 3392
rect 440234 3340 440240 3392
rect 440292 3380 440298 3392
rect 441522 3380 441528 3392
rect 440292 3352 441528 3380
rect 440292 3340 440298 3352
rect 441522 3340 441528 3352
rect 441580 3340 441586 3392
rect 448606 3340 448612 3392
rect 448664 3380 448670 3392
rect 449802 3380 449808 3392
rect 448664 3352 449808 3380
rect 448664 3340 448670 3352
rect 449802 3340 449808 3352
rect 449860 3340 449866 3392
rect 456794 3340 456800 3392
rect 456852 3380 456858 3392
rect 458082 3380 458088 3392
rect 456852 3352 458088 3380
rect 456852 3340 456858 3352
rect 458082 3340 458088 3352
rect 458140 3340 458146 3392
rect 571978 3340 571984 3392
rect 572036 3380 572042 3392
rect 576302 3380 576308 3392
rect 572036 3352 576308 3380
rect 572036 3340 572042 3352
rect 576302 3340 576308 3352
rect 576360 3340 576366 3392
rect 126974 3272 126980 3324
rect 127032 3312 127038 3324
rect 128446 3312 128452 3324
rect 127032 3284 128452 3312
rect 127032 3272 127038 3284
rect 128446 3272 128452 3284
rect 128504 3272 128510 3324
rect 193122 3272 193128 3324
rect 193180 3312 193186 3324
rect 195698 3312 195704 3324
rect 193180 3284 195704 3312
rect 193180 3272 193186 3284
rect 195698 3272 195704 3284
rect 195756 3272 195762 3324
rect 207750 3272 207756 3324
rect 207808 3312 207814 3324
rect 210970 3312 210976 3324
rect 207808 3284 210976 3312
rect 207808 3272 207814 3284
rect 210970 3272 210976 3284
rect 211028 3272 211034 3324
rect 431954 3272 431960 3324
rect 432012 3312 432018 3324
rect 433242 3312 433248 3324
rect 432012 3284 433248 3312
rect 432012 3272 432018 3284
rect 433242 3272 433248 3284
rect 433300 3272 433306 3324
rect 184198 3204 184204 3256
rect 184256 3244 184262 3256
rect 189718 3244 189724 3256
rect 184256 3216 189724 3244
rect 184256 3204 184262 3216
rect 189718 3204 189724 3216
rect 189776 3204 189782 3256
rect 520918 3204 520924 3256
rect 520976 3244 520982 3256
rect 524230 3244 524236 3256
rect 520976 3216 524236 3244
rect 520976 3204 520982 3216
rect 524230 3204 524236 3216
rect 524288 3204 524294 3256
rect 33594 3136 33600 3188
rect 33652 3176 33658 3188
rect 35158 3176 35164 3188
rect 33652 3148 35164 3176
rect 33652 3136 33658 3148
rect 35158 3136 35164 3148
rect 35216 3136 35222 3188
rect 38378 3136 38384 3188
rect 38436 3176 38442 3188
rect 39298 3176 39304 3188
rect 38436 3148 39304 3176
rect 38436 3136 38442 3148
rect 39298 3136 39304 3148
rect 39356 3136 39362 3188
rect 41874 3136 41880 3188
rect 41932 3176 41938 3188
rect 43438 3176 43444 3188
rect 41932 3148 43444 3176
rect 41932 3136 41938 3148
rect 43438 3136 43444 3148
rect 43496 3136 43502 3188
rect 136450 3136 136456 3188
rect 136508 3176 136514 3188
rect 141418 3176 141424 3188
rect 136508 3148 141424 3176
rect 136508 3136 136514 3148
rect 141418 3136 141424 3148
rect 141476 3136 141482 3188
rect 548518 3136 548524 3188
rect 548576 3176 548582 3188
rect 551462 3176 551468 3188
rect 548576 3148 551468 3176
rect 548576 3136 548582 3148
rect 551462 3136 551468 3148
rect 551520 3136 551526 3188
rect 12342 3068 12348 3120
rect 12400 3108 12406 3120
rect 17218 3108 17224 3120
rect 12400 3080 17224 3108
rect 12400 3068 12406 3080
rect 17218 3068 17224 3080
rect 17276 3068 17282 3120
rect 30098 3068 30104 3120
rect 30156 3108 30162 3120
rect 32398 3108 32404 3120
rect 30156 3080 32404 3108
rect 30156 3068 30162 3080
rect 32398 3068 32404 3080
rect 32456 3068 32462 3120
rect 124674 3068 124680 3120
rect 124732 3108 124738 3120
rect 131482 3108 131488 3120
rect 124732 3080 131488 3108
rect 124732 3068 124738 3080
rect 131482 3068 131488 3080
rect 131540 3068 131546 3120
rect 171870 3068 171876 3120
rect 171928 3108 171934 3120
rect 174262 3108 174268 3120
rect 171928 3080 174268 3108
rect 171928 3068 171934 3080
rect 174262 3068 174268 3080
rect 174320 3068 174326 3120
rect 382918 3068 382924 3120
rect 382976 3108 382982 3120
rect 384758 3108 384764 3120
rect 382976 3080 384764 3108
rect 382976 3068 382982 3080
rect 384758 3068 384764 3080
rect 384816 3068 384822 3120
rect 570598 3068 570604 3120
rect 570656 3108 570662 3120
rect 572714 3108 572720 3120
rect 570656 3080 572720 3108
rect 570656 3068 570662 3080
rect 572714 3068 572720 3080
rect 572772 3068 572778 3120
rect 20622 3000 20628 3052
rect 20680 3040 20686 3052
rect 22738 3040 22744 3052
rect 20680 3012 22744 3040
rect 20680 3000 20686 3012
rect 22738 3000 22744 3012
rect 22796 3000 22802 3052
rect 23014 3000 23020 3052
rect 23072 3040 23078 3052
rect 25498 3040 25504 3052
rect 23072 3012 25504 3040
rect 23072 3000 23078 3012
rect 25498 3000 25504 3012
rect 25556 3000 25562 3052
rect 118786 3000 118792 3052
rect 118844 3040 118850 3052
rect 121454 3040 121460 3052
rect 118844 3012 121460 3040
rect 118844 3000 118850 3012
rect 121454 3000 121460 3012
rect 121512 3000 121518 3052
rect 148410 3000 148416 3052
rect 148468 3040 148474 3052
rect 154206 3040 154212 3052
rect 148468 3012 154212 3040
rect 148468 3000 148474 3012
rect 154206 3000 154212 3012
rect 154264 3000 154270 3052
rect 464338 3000 464344 3052
rect 464396 3040 464402 3052
rect 466270 3040 466276 3052
rect 464396 3012 466276 3040
rect 464396 3000 464402 3012
rect 466270 3000 466276 3012
rect 466328 3000 466334 3052
rect 503070 3000 503076 3052
rect 503128 3040 503134 3052
rect 505370 3040 505376 3052
rect 503128 3012 505376 3040
rect 503128 3000 503134 3012
rect 505370 3000 505376 3012
rect 505428 3000 505434 3052
rect 514018 3000 514024 3052
rect 514076 3040 514082 3052
rect 515950 3040 515956 3052
rect 514076 3012 515956 3040
rect 514076 3000 514082 3012
rect 515950 3000 515956 3012
rect 516008 3000 516014 3052
rect 203518 2932 203524 2984
rect 203576 2972 203582 2984
rect 207382 2972 207388 2984
rect 203576 2944 207388 2972
rect 203576 2932 203582 2944
rect 207382 2932 207388 2944
rect 207440 2932 207446 2984
rect 220078 2932 220084 2984
rect 220136 2972 220142 2984
rect 225138 2972 225144 2984
rect 220136 2944 225144 2972
rect 220136 2932 220142 2944
rect 225138 2932 225144 2944
rect 225196 2932 225202 2984
rect 509878 2932 509884 2984
rect 509936 2972 509942 2984
rect 514754 2972 514760 2984
rect 509936 2944 514760 2972
rect 509936 2932 509942 2944
rect 514754 2932 514760 2944
rect 514812 2932 514818 2984
rect 171778 2864 171784 2916
rect 171836 2904 171842 2916
rect 177850 2904 177856 2916
rect 171836 2876 177856 2904
rect 171836 2864 171842 2876
rect 177850 2864 177856 2876
rect 177908 2864 177914 2916
rect 260098 2864 260104 2916
rect 260156 2904 260162 2916
rect 261754 2904 261760 2916
rect 260156 2876 261760 2904
rect 260156 2864 260162 2876
rect 261754 2864 261760 2876
rect 261812 2864 261818 2916
rect 390554 1776 390560 1828
rect 390612 1816 390618 1828
rect 391842 1816 391848 1828
rect 390612 1788 391848 1816
rect 390612 1776 390618 1788
rect 391842 1776 391848 1788
rect 391900 1776 391906 1828
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 137836 700816 137888 700868
rect 157984 700816 158036 700868
rect 155960 700748 156012 700800
rect 202788 700748 202840 700800
rect 89168 700680 89220 700732
rect 160744 700680 160796 700732
rect 154580 700612 154632 700664
rect 267648 700612 267700 700664
rect 24308 700544 24360 700596
rect 162216 700544 162268 700596
rect 8116 700476 8168 700528
rect 162124 700476 162176 700528
rect 153844 700408 153896 700460
rect 332508 700408 332560 700460
rect 152464 700340 152516 700392
rect 413652 700340 413704 700392
rect 148324 700272 148376 700324
rect 543464 700272 543516 700324
rect 543004 700204 543056 700256
rect 559656 700272 559708 700324
rect 105452 699660 105504 699712
rect 106924 699660 106976 699712
rect 396724 699660 396776 699712
rect 397460 699660 397512 699712
rect 428464 699660 428516 699712
rect 429844 699660 429896 699712
rect 146944 696940 146996 696992
rect 580172 696940 580224 696992
rect 3424 683204 3476 683256
rect 161480 683204 161532 683256
rect 147036 683136 147088 683188
rect 580172 683136 580224 683188
rect 3516 670692 3568 670744
rect 163504 670692 163556 670744
rect 185584 670692 185636 670744
rect 580172 670692 580224 670744
rect 149060 660288 149112 660340
rect 462320 660288 462372 660340
rect 3424 656888 3476 656940
rect 163596 656888 163648 656940
rect 184204 643084 184256 643136
rect 580172 643084 580224 643136
rect 3424 632068 3476 632120
rect 164240 632068 164292 632120
rect 203524 630640 203576 630692
rect 580172 630640 580224 630692
rect 3148 618264 3200 618316
rect 164884 618264 164936 618316
rect 143540 616836 143592 616888
rect 580172 616836 580224 616888
rect 3240 605820 3292 605872
rect 164976 605820 165028 605872
rect 142160 590656 142212 590708
rect 579804 590656 579856 590708
rect 3332 579640 3384 579692
rect 165620 579640 165672 579692
rect 144184 576852 144236 576904
rect 580172 576852 580224 576904
rect 3424 565836 3476 565888
rect 167644 565836 167696 565888
rect 142804 563048 142856 563100
rect 579804 563048 579856 563100
rect 3424 553392 3476 553444
rect 166264 553392 166316 553444
rect 178684 536800 178736 536852
rect 580172 536800 580224 536852
rect 3424 527144 3476 527196
rect 167000 527144 167052 527196
rect 142896 524424 142948 524476
rect 580172 524424 580224 524476
rect 3424 514768 3476 514820
rect 8944 514768 8996 514820
rect 181444 510620 181496 510672
rect 580172 510620 580224 510672
rect 3056 500964 3108 501016
rect 167276 500964 167328 501016
rect 139400 484372 139452 484424
rect 580172 484372 580224 484424
rect 139676 470568 139728 470620
rect 579988 470568 580040 470620
rect 3516 462340 3568 462392
rect 170404 462340 170456 462392
rect 180064 456764 180116 456816
rect 580172 456764 580224 456816
rect 3148 448536 3200 448588
rect 170496 448536 170548 448588
rect 158628 447788 158680 447840
rect 169760 447788 169812 447840
rect 138664 430584 138716 430636
rect 580172 430584 580224 430636
rect 3516 422288 3568 422340
rect 169760 422288 169812 422340
rect 138756 418140 138808 418192
rect 580172 418140 580224 418192
rect 2872 409844 2924 409896
rect 171784 409844 171836 409896
rect 199384 404336 199436 404388
rect 580172 404336 580224 404388
rect 3516 397468 3568 397520
rect 171876 397468 171928 397520
rect 182824 378156 182876 378208
rect 580172 378156 580224 378208
rect 2780 371288 2832 371340
rect 4804 371288 4856 371340
rect 3148 357416 3200 357468
rect 10324 357416 10376 357468
rect 135260 351908 135312 351960
rect 580172 351908 580224 351960
rect 3516 345176 3568 345228
rect 7564 345176 7616 345228
rect 134524 324300 134576 324352
rect 580172 324300 580224 324352
rect 3332 318792 3384 318844
rect 173900 318792 173952 318844
rect 135904 311856 135956 311908
rect 579988 311856 580040 311908
rect 3516 304988 3568 305040
rect 175924 304988 175976 305040
rect 134616 298120 134668 298172
rect 580172 298120 580224 298172
rect 3516 292544 3568 292596
rect 174544 292544 174596 292596
rect 10324 289076 10376 289128
rect 173164 289076 173216 289128
rect 145564 287648 145616 287700
rect 203524 287648 203576 287700
rect 137284 286288 137336 286340
rect 182824 286288 182876 286340
rect 150440 284928 150492 284980
rect 396724 284928 396776 284980
rect 147680 283568 147732 283620
rect 527180 283568 527232 283620
rect 145656 282140 145708 282192
rect 184204 282140 184256 282192
rect 140780 280780 140832 280832
rect 178684 280780 178736 280832
rect 40040 279420 40092 279472
rect 160100 279420 160152 279472
rect 189080 277992 189132 278044
rect 234620 277992 234672 278044
rect 156052 277380 156104 277432
rect 189080 277380 189132 277432
rect 204720 276632 204772 276684
rect 299480 276632 299532 276684
rect 153292 276020 153344 276072
rect 204444 276020 204496 276072
rect 204720 276020 204772 276072
rect 8944 273980 8996 274032
rect 169024 273980 169076 274032
rect 151084 273912 151136 273964
rect 428464 273912 428516 273964
rect 133144 271872 133196 271924
rect 580172 271872 580224 271924
rect 7564 271192 7616 271244
rect 172520 271192 172572 271244
rect 149152 271124 149204 271176
rect 494060 271124 494112 271176
rect 71780 269832 71832 269884
rect 158812 269832 158864 269884
rect 147772 269764 147824 269816
rect 543004 269764 543056 269816
rect 146208 268404 146260 268456
rect 185584 268404 185636 268456
rect 4804 268336 4856 268388
rect 172704 268336 172756 268388
rect 137836 266976 137888 267028
rect 199384 266976 199436 267028
rect 3056 266364 3108 266416
rect 175924 266364 175976 266416
rect 164884 265820 164936 265872
rect 165160 265820 165212 265872
rect 141424 265684 141476 265736
rect 181444 265684 181496 265736
rect 3424 265616 3476 265668
rect 169116 265616 169168 265668
rect 174544 265548 174596 265600
rect 195980 265480 196032 265532
rect 166264 265412 166316 265464
rect 192116 265412 192168 265464
rect 171784 265344 171836 265396
rect 197636 265344 197688 265396
rect 173440 265276 173492 265328
rect 199200 265276 199252 265328
rect 170404 265208 170456 265260
rect 170680 265208 170732 265260
rect 199108 265208 199160 265260
rect 113088 265140 113140 265192
rect 138756 265140 138808 265192
rect 162216 265140 162268 265192
rect 195244 265140 195296 265192
rect 116584 265072 116636 265124
rect 143632 265072 143684 265124
rect 144184 265072 144236 265124
rect 170220 265072 170272 265124
rect 170496 265072 170548 265124
rect 203248 265072 203300 265124
rect 112812 265004 112864 265056
rect 145564 265004 145616 265056
rect 160836 265004 160888 265056
rect 194876 265004 194928 265056
rect 119620 264936 119672 264988
rect 152188 264936 152240 264988
rect 152464 264936 152516 264988
rect 165160 264936 165212 264988
rect 203156 264936 203208 264988
rect 106924 264188 106976 264240
rect 118700 264188 118752 264240
rect 139400 264188 139452 264240
rect 180064 264188 180116 264240
rect 121000 263916 121052 263968
rect 134248 263916 134300 263968
rect 134616 263916 134668 263968
rect 119528 263848 119580 263900
rect 137836 263848 137888 263900
rect 120908 263780 120960 263832
rect 139400 263780 139452 263832
rect 117964 263712 118016 263764
rect 137192 263712 137244 263764
rect 172704 263712 172756 263764
rect 190644 263712 190696 263764
rect 119712 263644 119764 263696
rect 141148 263644 141200 263696
rect 141424 263644 141476 263696
rect 157892 263644 157944 263696
rect 158628 263644 158680 263696
rect 188252 263644 188304 263696
rect 118700 263576 118752 263628
rect 119988 263576 120040 263628
rect 159088 263576 159140 263628
rect 175740 263576 175792 263628
rect 197728 263576 197780 263628
rect 137468 263508 137520 263560
rect 580264 263508 580316 263560
rect 190000 263440 190052 263492
rect 282920 263440 282972 263492
rect 171692 263372 171744 263424
rect 171876 263372 171928 263424
rect 163412 263236 163464 263288
rect 163596 263236 163648 263288
rect 116860 263100 116912 263152
rect 129280 263100 129332 263152
rect 171692 263100 171744 263152
rect 196624 263100 196676 263152
rect 3424 263032 3476 263084
rect 178408 263032 178460 263084
rect 180156 263032 180208 263084
rect 194968 263032 195020 263084
rect 117044 262964 117096 263016
rect 125968 262964 126020 263016
rect 132316 262964 132368 263016
rect 580356 262964 580408 263016
rect 116676 262896 116728 262948
rect 127532 262896 127584 262948
rect 115388 262828 115440 262880
rect 131764 262828 131816 262880
rect 580448 262896 580500 262948
rect 115480 262760 115532 262812
rect 134524 262760 134576 262812
rect 134800 262760 134852 262812
rect 153200 262760 153252 262812
rect 158720 262760 158772 262812
rect 164976 262760 165028 262812
rect 193588 262760 193640 262812
rect 118332 262692 118384 262744
rect 122840 262692 122892 262744
rect 127532 262692 127584 262744
rect 133144 262692 133196 262744
rect 163412 262692 163464 262744
rect 192484 262692 192536 262744
rect 118240 262624 118292 262676
rect 127624 262624 127676 262676
rect 157984 262624 158036 262676
rect 192208 262624 192260 262676
rect 114008 262556 114060 262608
rect 129832 262556 129884 262608
rect 155868 262556 155920 262608
rect 189264 262556 189316 262608
rect 190000 262556 190052 262608
rect 119804 262488 119856 262540
rect 153292 262488 153344 262540
rect 153844 262488 153896 262540
rect 157156 262488 157208 262540
rect 192392 262488 192444 262540
rect 218060 262828 218112 262880
rect 3516 262420 3568 262472
rect 176752 262420 176804 262472
rect 179236 262420 179288 262472
rect 192668 262420 192720 262472
rect 122840 262352 122892 262404
rect 131120 262352 131172 262404
rect 182916 262352 182968 262404
rect 190460 262352 190512 262404
rect 181260 262284 181312 262336
rect 190552 262284 190604 262336
rect 116492 262216 116544 262268
rect 122748 262216 122800 262268
rect 184572 262216 184624 262268
rect 189172 262216 189224 262268
rect 158720 261604 158772 261656
rect 193680 261604 193732 261656
rect 129832 261536 129884 261588
rect 189816 261536 189868 261588
rect 176752 261468 176804 261520
rect 199292 261468 199344 261520
rect 131120 261400 131172 261452
rect 471244 261400 471296 261452
rect 181812 261332 181864 261384
rect 193496 261332 193548 261384
rect 177304 261264 177356 261316
rect 193772 261264 193824 261316
rect 178408 261196 178460 261248
rect 197912 261196 197964 261248
rect 112904 261128 112956 261180
rect 128728 261128 128780 261180
rect 176200 261128 176252 261180
rect 195060 261128 195112 261180
rect 116768 261060 116820 261112
rect 133236 261060 133288 261112
rect 184020 261060 184072 261112
rect 196440 261060 196492 261112
rect 111064 260992 111116 261044
rect 127072 260992 127124 261044
rect 180524 260992 180576 261044
rect 198004 260992 198056 261044
rect 4804 260924 4856 260976
rect 176200 260924 176252 260976
rect 184756 260924 184808 260976
rect 197084 260924 197136 260976
rect 112628 260856 112680 260908
rect 130384 260856 130436 260908
rect 181996 260856 182048 260908
rect 197820 260856 197872 260908
rect 119896 260788 119948 260840
rect 124312 260788 124364 260840
rect 119252 260720 119304 260772
rect 122840 260720 122892 260772
rect 122748 260652 122800 260704
rect 123208 260652 123260 260704
rect 180800 260516 180852 260568
rect 189540 260516 189592 260568
rect 173900 260448 173952 260500
rect 185584 260448 185636 260500
rect 133236 260380 133288 260432
rect 485044 260380 485096 260432
rect 7564 260312 7616 260364
rect 177304 260312 177356 260364
rect 114192 260244 114244 260296
rect 126520 260244 126572 260296
rect 118148 260176 118200 260228
rect 164240 260244 164292 260296
rect 175832 260244 175884 260296
rect 135260 260176 135312 260228
rect 136226 260176 136278 260228
rect 139492 260176 139544 260228
rect 140090 260176 140142 260228
rect 143540 260176 143592 260228
rect 144506 260176 144558 260228
rect 155960 260176 156012 260228
rect 156650 260176 156702 260228
rect 167276 260176 167328 260228
rect 168242 260176 168294 260228
rect 169760 260176 169812 260228
rect 171002 260176 171054 260228
rect 172520 260176 172572 260228
rect 173210 260176 173262 260228
rect 175924 260176 175976 260228
rect 192300 260312 192352 260364
rect 185584 260244 185636 260296
rect 193864 260244 193916 260296
rect 113732 260108 113784 260160
rect 139676 260108 139728 260160
rect 140642 260108 140694 260160
rect 167000 260108 167052 260160
rect 167690 260108 167742 260160
rect 180800 260108 180852 260160
rect 118056 260040 118108 260092
rect 135076 260040 135128 260092
rect 169346 260040 169398 260092
rect 191012 260176 191064 260228
rect 112444 259972 112496 260024
rect 132040 259972 132092 260024
rect 189724 260108 189776 260160
rect 120632 259904 120684 259956
rect 142160 259904 142212 259956
rect 143080 259904 143132 259956
rect 168380 259904 168432 259956
rect 119344 259836 119396 259888
rect 143540 259836 143592 259888
rect 166172 259836 166224 259888
rect 183284 259904 183336 259956
rect 175832 259836 175884 259888
rect 189632 260040 189684 260092
rect 183468 259972 183520 260024
rect 190920 260040 190972 260092
rect 183468 259836 183520 259888
rect 192576 259904 192628 259956
rect 117872 259768 117924 259820
rect 150440 259768 150492 259820
rect 151360 259768 151412 259820
rect 171140 259768 171192 259820
rect 201868 259768 201920 259820
rect 115020 259700 115072 259752
rect 149060 259700 149112 259752
rect 149704 259700 149756 259752
rect 156972 259700 157024 259752
rect 185768 259700 185820 259752
rect 113824 259632 113876 259684
rect 123760 259632 123812 259684
rect 134340 259632 134392 259684
rect 187700 259632 187752 259684
rect 117780 259564 117832 259616
rect 178040 259564 178092 259616
rect 196716 259564 196768 259616
rect 114100 259496 114152 259548
rect 124864 259496 124916 259548
rect 173348 259496 173400 259548
rect 201960 259496 202012 259548
rect 115204 259428 115256 259480
rect 128360 259428 128412 259480
rect 185768 259428 185820 259480
rect 190736 259428 190788 259480
rect 187700 259360 187752 259412
rect 580172 259360 580224 259412
rect 485044 245556 485096 245608
rect 580172 245556 580224 245608
rect 2780 241204 2832 241256
rect 4804 241204 4856 241256
rect 3516 215092 3568 215144
rect 7564 215092 7616 215144
rect 471244 206932 471296 206984
rect 579804 206932 579856 206984
rect 126244 200676 126296 200728
rect 132224 200676 132276 200728
rect 107292 200540 107344 200592
rect 129004 200608 129056 200660
rect 128544 200540 128596 200592
rect 131948 200540 132000 200592
rect 104808 200472 104860 200524
rect 131580 200472 131632 200524
rect 132224 200540 132276 200592
rect 121368 200336 121420 200388
rect 132224 200404 132276 200456
rect 132040 200336 132092 200388
rect 130292 200268 130344 200320
rect 110236 200200 110288 200252
rect 127624 200200 127676 200252
rect 132224 200200 132276 200252
rect 130476 200132 130528 200184
rect 132040 200132 132092 200184
rect 131488 200064 131540 200116
rect 130384 199996 130436 200048
rect 131856 199996 131908 200048
rect 132224 199928 132276 199980
rect 119896 199860 119948 199912
rect 125140 199860 125192 199912
rect 128360 199860 128412 199912
rect 132638 199860 132690 199912
rect 132914 199860 132966 199912
rect 133742 199860 133794 199912
rect 127532 199792 127584 199844
rect 129004 199724 129056 199776
rect 132960 199724 133012 199776
rect 111708 199656 111760 199708
rect 130476 199656 130528 199708
rect 130568 199656 130620 199708
rect 132316 199656 132368 199708
rect 109868 199588 109920 199640
rect 130384 199588 130436 199640
rect 114468 199520 114520 199572
rect 132316 199520 132368 199572
rect 114376 199452 114428 199504
rect 132224 199452 132276 199504
rect 133926 199860 133978 199912
rect 134018 199860 134070 199912
rect 134202 199860 134254 199912
rect 134294 199860 134346 199912
rect 134478 199860 134530 199912
rect 134570 199860 134622 199912
rect 134662 199860 134714 199912
rect 134846 199860 134898 199912
rect 134938 199860 134990 199912
rect 135122 199860 135174 199912
rect 135306 199860 135358 199912
rect 135490 199860 135542 199912
rect 133788 199588 133840 199640
rect 134248 199656 134300 199708
rect 134064 199588 134116 199640
rect 134156 199588 134208 199640
rect 133972 199452 134024 199504
rect 132868 199384 132920 199436
rect 132960 199384 133012 199436
rect 133880 199384 133932 199436
rect 134524 199588 134576 199640
rect 134892 199724 134944 199776
rect 134800 199656 134852 199708
rect 135168 199588 135220 199640
rect 134340 199520 134392 199572
rect 135260 199520 135312 199572
rect 135352 199520 135404 199572
rect 135444 199520 135496 199572
rect 135674 199860 135726 199912
rect 136042 199860 136094 199912
rect 136226 199860 136278 199912
rect 136318 199860 136370 199912
rect 136686 199860 136738 199912
rect 137054 199860 137106 199912
rect 137238 199860 137290 199912
rect 137330 199860 137382 199912
rect 135720 199520 135772 199572
rect 137284 199724 137336 199776
rect 137100 199656 137152 199708
rect 137606 199860 137658 199912
rect 137698 199860 137750 199912
rect 137790 199860 137842 199912
rect 137882 199860 137934 199912
rect 138066 199860 138118 199912
rect 138158 199860 138210 199912
rect 138250 199860 138302 199912
rect 138434 199860 138486 199912
rect 137652 199724 137704 199776
rect 137744 199724 137796 199776
rect 138112 199724 138164 199776
rect 138204 199724 138256 199776
rect 137836 199656 137888 199708
rect 136272 199588 136324 199640
rect 136732 199588 136784 199640
rect 137468 199588 137520 199640
rect 137560 199588 137612 199640
rect 136640 199520 136692 199572
rect 138388 199724 138440 199776
rect 138618 199860 138670 199912
rect 138986 199860 139038 199912
rect 139354 199860 139406 199912
rect 139446 199860 139498 199912
rect 139630 199860 139682 199912
rect 139722 199860 139774 199912
rect 138572 199656 138624 199708
rect 138940 199588 138992 199640
rect 139492 199656 139544 199708
rect 139814 199792 139866 199844
rect 139998 199792 140050 199844
rect 139860 199656 139912 199708
rect 139952 199656 140004 199708
rect 140274 199860 140326 199912
rect 140458 199860 140510 199912
rect 140550 199860 140602 199912
rect 140826 199860 140878 199912
rect 141010 199860 141062 199912
rect 141102 199860 141154 199912
rect 141286 199860 141338 199912
rect 141378 199860 141430 199912
rect 141746 199860 141798 199912
rect 141838 199860 141890 199912
rect 140182 199656 140234 199708
rect 134432 199384 134484 199436
rect 134616 199384 134668 199436
rect 135996 199452 136048 199504
rect 138020 199452 138072 199504
rect 139768 199520 139820 199572
rect 140136 199520 140188 199572
rect 138756 199452 138808 199504
rect 139032 199452 139084 199504
rect 139124 199452 139176 199504
rect 140596 199588 140648 199640
rect 140412 199520 140464 199572
rect 140872 199724 140924 199776
rect 141148 199724 141200 199776
rect 140780 199588 140832 199640
rect 141240 199520 141292 199572
rect 141470 199724 141522 199776
rect 141516 199588 141568 199640
rect 141332 199452 141384 199504
rect 141424 199452 141476 199504
rect 141792 199452 141844 199504
rect 142022 199860 142074 199912
rect 142390 199860 142442 199912
rect 143218 199860 143270 199912
rect 142942 199792 142994 199844
rect 142022 199656 142074 199708
rect 142988 199520 143040 199572
rect 143264 199520 143316 199572
rect 143770 199792 143822 199844
rect 143862 199792 143914 199844
rect 143954 199792 144006 199844
rect 144138 199792 144190 199844
rect 143586 199656 143638 199708
rect 143908 199656 143960 199708
rect 144092 199656 144144 199708
rect 144506 199860 144558 199912
rect 144598 199860 144650 199912
rect 144690 199860 144742 199912
rect 144782 199860 144834 199912
rect 144552 199656 144604 199708
rect 144644 199656 144696 199708
rect 144736 199656 144788 199708
rect 144966 199860 145018 199912
rect 145058 199860 145110 199912
rect 145012 199724 145064 199776
rect 145702 199860 145754 199912
rect 145334 199724 145386 199776
rect 144368 199588 144420 199640
rect 144828 199588 144880 199640
rect 143540 199520 143592 199572
rect 143632 199520 143684 199572
rect 145288 199520 145340 199572
rect 145886 199860 145938 199912
rect 146070 199860 146122 199912
rect 146162 199860 146214 199912
rect 146254 199860 146306 199912
rect 143816 199452 143868 199504
rect 137008 199384 137060 199436
rect 137192 199384 137244 199436
rect 144276 199384 144328 199436
rect 145656 199384 145708 199436
rect 146208 199724 146260 199776
rect 146024 199588 146076 199640
rect 146438 199860 146490 199912
rect 146806 199860 146858 199912
rect 146990 199860 147042 199912
rect 147542 199860 147594 199912
rect 146484 199724 146536 199776
rect 146300 199452 146352 199504
rect 146116 199384 146168 199436
rect 146760 199588 146812 199640
rect 147818 199792 147870 199844
rect 148462 199792 148514 199844
rect 148646 199792 148698 199844
rect 147496 199724 147548 199776
rect 147588 199656 147640 199708
rect 148370 199656 148422 199708
rect 147312 199588 147364 199640
rect 148600 199656 148652 199708
rect 149106 199860 149158 199912
rect 149198 199860 149250 199912
rect 149474 199860 149526 199912
rect 149842 199860 149894 199912
rect 149152 199656 149204 199708
rect 149658 199792 149710 199844
rect 149612 199588 149664 199640
rect 149428 199520 149480 199572
rect 149060 199452 149112 199504
rect 148324 199384 148376 199436
rect 150026 199860 150078 199912
rect 150210 199860 150262 199912
rect 150486 199860 150538 199912
rect 150578 199860 150630 199912
rect 150670 199860 150722 199912
rect 150946 199860 150998 199912
rect 151038 199860 151090 199912
rect 151222 199860 151274 199912
rect 151314 199860 151366 199912
rect 151406 199860 151458 199912
rect 151682 199860 151734 199912
rect 150302 199792 150354 199844
rect 150440 199724 150492 199776
rect 150532 199724 150584 199776
rect 150854 199792 150906 199844
rect 150256 199656 150308 199708
rect 150716 199656 150768 199708
rect 150808 199656 150860 199708
rect 150164 199588 150216 199640
rect 150072 199520 150124 199572
rect 151084 199588 151136 199640
rect 151176 199588 151228 199640
rect 151452 199724 151504 199776
rect 151636 199588 151688 199640
rect 151268 199520 151320 199572
rect 151866 199860 151918 199912
rect 152050 199860 152102 199912
rect 152142 199860 152194 199912
rect 152234 199860 152286 199912
rect 151912 199656 151964 199708
rect 152418 199792 152470 199844
rect 152096 199656 152148 199708
rect 152188 199656 152240 199708
rect 152372 199588 152424 199640
rect 152694 199860 152746 199912
rect 152786 199860 152838 199912
rect 152970 199860 153022 199912
rect 153062 199860 153114 199912
rect 153154 199860 153206 199912
rect 153338 199860 153390 199912
rect 153430 199860 153482 199912
rect 153614 199860 153666 199912
rect 153706 199860 153758 199912
rect 152740 199724 152792 199776
rect 153016 199724 153068 199776
rect 153108 199724 153160 199776
rect 153200 199724 153252 199776
rect 153384 199724 153436 199776
rect 153568 199724 153620 199776
rect 153476 199656 153528 199708
rect 152924 199588 152976 199640
rect 153660 199588 153712 199640
rect 153982 199860 154034 199912
rect 154074 199860 154126 199912
rect 154166 199860 154218 199912
rect 154258 199860 154310 199912
rect 154442 199860 154494 199912
rect 154028 199656 154080 199708
rect 154212 199588 154264 199640
rect 154120 199520 154172 199572
rect 154626 199792 154678 199844
rect 154718 199792 154770 199844
rect 155086 199860 155138 199912
rect 154534 199588 154586 199640
rect 154396 199520 154448 199572
rect 154948 199520 155000 199572
rect 154672 199452 154724 199504
rect 154856 199452 154908 199504
rect 155362 199792 155414 199844
rect 156558 199860 156610 199912
rect 155638 199792 155690 199844
rect 155822 199792 155874 199844
rect 156006 199792 156058 199844
rect 156190 199792 156242 199844
rect 156282 199792 156334 199844
rect 155684 199656 155736 199708
rect 155868 199656 155920 199708
rect 156052 199656 156104 199708
rect 156236 199656 156288 199708
rect 156926 199724 156978 199776
rect 157478 199860 157530 199912
rect 157294 199792 157346 199844
rect 157386 199792 157438 199844
rect 157432 199656 157484 199708
rect 155592 199588 155644 199640
rect 156512 199588 156564 199640
rect 156880 199588 156932 199640
rect 157156 199588 157208 199640
rect 157340 199588 157392 199640
rect 155316 199520 155368 199572
rect 157662 199860 157714 199912
rect 158122 199860 158174 199912
rect 158490 199860 158542 199912
rect 158674 199860 158726 199912
rect 157708 199656 157760 199708
rect 157938 199724 157990 199776
rect 157892 199520 157944 199572
rect 157248 199452 157300 199504
rect 157524 199452 157576 199504
rect 157616 199452 157668 199504
rect 158122 199724 158174 199776
rect 158582 199792 158634 199844
rect 159042 199792 159094 199844
rect 158444 199588 158496 199640
rect 158536 199588 158588 199640
rect 159226 199860 159278 199912
rect 159318 199860 159370 199912
rect 159410 199860 159462 199912
rect 159594 199860 159646 199912
rect 159686 199860 159738 199912
rect 160146 199860 160198 199912
rect 159272 199724 159324 199776
rect 159088 199588 159140 199640
rect 159364 199656 159416 199708
rect 159640 199656 159692 199708
rect 160054 199792 160106 199844
rect 159548 199588 159600 199640
rect 159732 199588 159784 199640
rect 158076 199520 158128 199572
rect 159456 199520 159508 199572
rect 160192 199520 160244 199572
rect 160606 199860 160658 199912
rect 160698 199860 160750 199912
rect 160560 199656 160612 199708
rect 160882 199792 160934 199844
rect 160974 199792 161026 199844
rect 160744 199588 160796 199640
rect 160652 199520 160704 199572
rect 160928 199656 160980 199708
rect 161158 199860 161210 199912
rect 161250 199860 161302 199912
rect 161434 199860 161486 199912
rect 161526 199860 161578 199912
rect 161710 199860 161762 199912
rect 161802 199860 161854 199912
rect 161894 199860 161946 199912
rect 162170 199860 162222 199912
rect 162354 199860 162406 199912
rect 162446 199860 162498 199912
rect 162538 199860 162590 199912
rect 162630 199860 162682 199912
rect 161204 199724 161256 199776
rect 161480 199724 161532 199776
rect 161664 199724 161716 199776
rect 161756 199724 161808 199776
rect 162308 199724 162360 199776
rect 162400 199724 162452 199776
rect 161388 199656 161440 199708
rect 161848 199656 161900 199708
rect 162124 199656 162176 199708
rect 162584 199656 162636 199708
rect 161480 199588 161532 199640
rect 161572 199588 161624 199640
rect 161204 199520 161256 199572
rect 162400 199452 162452 199504
rect 162998 199860 163050 199912
rect 156236 199384 156288 199436
rect 160192 199384 160244 199436
rect 161388 199384 161440 199436
rect 118608 199316 118660 199368
rect 118424 199248 118476 199300
rect 135076 199248 135128 199300
rect 145104 199316 145156 199368
rect 145196 199316 145248 199368
rect 148416 199316 148468 199368
rect 150624 199316 150676 199368
rect 135720 199248 135772 199300
rect 146208 199248 146260 199300
rect 149520 199248 149572 199300
rect 117228 199180 117280 199232
rect 145380 199180 145432 199232
rect 115756 199112 115808 199164
rect 145932 199112 145984 199164
rect 157800 199248 157852 199300
rect 158720 199248 158772 199300
rect 159548 199316 159600 199368
rect 162032 199316 162084 199368
rect 162492 199316 162544 199368
rect 163274 199860 163326 199912
rect 163366 199860 163418 199912
rect 163274 199724 163326 199776
rect 163274 199588 163326 199640
rect 163412 199588 163464 199640
rect 163228 199452 163280 199504
rect 163320 199384 163372 199436
rect 163918 199860 163970 199912
rect 163826 199792 163878 199844
rect 164286 199860 164338 199912
rect 163872 199656 163924 199708
rect 164332 199724 164384 199776
rect 164562 199860 164614 199912
rect 164240 199588 164292 199640
rect 164424 199588 164476 199640
rect 163688 199520 163740 199572
rect 163964 199520 164016 199572
rect 164608 199520 164660 199572
rect 164838 199792 164890 199844
rect 164930 199792 164982 199844
rect 165022 199792 165074 199844
rect 165298 199792 165350 199844
rect 165160 199588 165212 199640
rect 165666 199724 165718 199776
rect 165620 199588 165672 199640
rect 165712 199520 165764 199572
rect 163596 199384 163648 199436
rect 164516 199452 164568 199504
rect 164792 199452 164844 199504
rect 164976 199452 165028 199504
rect 165344 199452 165396 199504
rect 166402 199860 166454 199912
rect 166494 199860 166546 199912
rect 166586 199860 166638 199912
rect 166678 199860 166730 199912
rect 166770 199860 166822 199912
rect 166356 199724 166408 199776
rect 166540 199724 166592 199776
rect 166448 199656 166500 199708
rect 166632 199656 166684 199708
rect 167046 199860 167098 199912
rect 167506 199860 167558 199912
rect 167598 199860 167650 199912
rect 166908 199588 166960 199640
rect 166724 199520 166776 199572
rect 167322 199792 167374 199844
rect 167276 199588 167328 199640
rect 167368 199520 167420 199572
rect 166264 199452 166316 199504
rect 167552 199656 167604 199708
rect 167782 199656 167834 199708
rect 167736 199520 167788 199572
rect 168150 199860 168202 199912
rect 168242 199860 168294 199912
rect 168196 199656 168248 199708
rect 168104 199588 168156 199640
rect 168518 199724 168570 199776
rect 168426 199656 168478 199708
rect 168794 199860 168846 199912
rect 168886 199860 168938 199912
rect 169070 199792 169122 199844
rect 168932 199724 168984 199776
rect 168840 199656 168892 199708
rect 169024 199656 169076 199708
rect 177764 200676 177816 200728
rect 178868 200676 178920 200728
rect 179972 200676 180024 200728
rect 178684 200608 178736 200660
rect 189080 200744 189132 200796
rect 180248 200676 180300 200728
rect 177856 200540 177908 200592
rect 178776 200540 178828 200592
rect 199016 200404 199068 200456
rect 177764 200336 177816 200388
rect 193312 200336 193364 200388
rect 187700 200268 187752 200320
rect 186688 200200 186740 200252
rect 169254 199792 169306 199844
rect 169438 199792 169490 199844
rect 169530 199792 169582 199844
rect 168564 199588 168616 199640
rect 168656 199588 168708 199640
rect 169116 199588 169168 199640
rect 168288 199520 168340 199572
rect 168380 199520 168432 199572
rect 168472 199452 168524 199504
rect 169116 199452 169168 199504
rect 169392 199588 169444 199640
rect 169484 199588 169536 199640
rect 169576 199520 169628 199572
rect 170174 199792 170226 199844
rect 170220 199656 170272 199708
rect 170450 199792 170502 199844
rect 170404 199520 170456 199572
rect 171002 199860 171054 199912
rect 171094 199860 171146 199912
rect 170818 199792 170870 199844
rect 170726 199724 170778 199776
rect 171048 199656 171100 199708
rect 171462 199860 171514 199912
rect 171554 199860 171606 199912
rect 171140 199588 171192 199640
rect 171232 199588 171284 199640
rect 170772 199520 170824 199572
rect 169944 199452 169996 199504
rect 170496 199452 170548 199504
rect 171738 199792 171790 199844
rect 172014 199860 172066 199912
rect 172382 199860 172434 199912
rect 213920 200132 213972 200184
rect 172382 199724 172434 199776
rect 171692 199588 171744 199640
rect 171876 199588 171928 199640
rect 172152 199588 172204 199640
rect 172244 199588 172296 199640
rect 172060 199520 172112 199572
rect 172336 199520 172388 199572
rect 171508 199452 171560 199504
rect 172428 199452 172480 199504
rect 172842 199860 172894 199912
rect 173026 199792 173078 199844
rect 178040 199996 178092 200048
rect 173210 199724 173262 199776
rect 173762 199860 173814 199912
rect 173854 199860 173906 199912
rect 173946 199860 173998 199912
rect 173808 199724 173860 199776
rect 173900 199724 173952 199776
rect 174130 199860 174182 199912
rect 181996 199928 182048 199980
rect 174498 199860 174550 199912
rect 174774 199860 174826 199912
rect 174866 199860 174918 199912
rect 174958 199860 175010 199912
rect 174452 199724 174504 199776
rect 174682 199792 174734 199844
rect 174544 199656 174596 199708
rect 173808 199520 173860 199572
rect 172704 199452 172756 199504
rect 172980 199452 173032 199504
rect 174268 199588 174320 199640
rect 173992 199520 174044 199572
rect 174544 199520 174596 199572
rect 174912 199656 174964 199708
rect 175326 199860 175378 199912
rect 175510 199860 175562 199912
rect 175418 199792 175470 199844
rect 175372 199588 175424 199640
rect 175970 199860 176022 199912
rect 176062 199860 176114 199912
rect 176798 199860 176850 199912
rect 176890 199860 176942 199912
rect 178868 199860 178920 199912
rect 176016 199724 176068 199776
rect 177672 199792 177724 199844
rect 180156 199792 180208 199844
rect 176844 199724 176896 199776
rect 180340 199724 180392 199776
rect 187884 199724 187936 199776
rect 175924 199588 175976 199640
rect 176752 199588 176804 199640
rect 177672 199588 177724 199640
rect 214012 199656 214064 199708
rect 177948 199588 178000 199640
rect 215852 199588 215904 199640
rect 174176 199452 174228 199504
rect 174268 199452 174320 199504
rect 174728 199452 174780 199504
rect 174820 199452 174872 199504
rect 175188 199452 175240 199504
rect 175648 199452 175700 199504
rect 163964 199384 164016 199436
rect 169208 199384 169260 199436
rect 169760 199384 169812 199436
rect 175924 199452 175976 199504
rect 180156 199452 180208 199504
rect 182916 199452 182968 199504
rect 190460 199452 190512 199504
rect 181076 199384 181128 199436
rect 190552 199384 190604 199436
rect 157248 199180 157300 199232
rect 161664 199180 161716 199232
rect 215576 199316 215628 199368
rect 163688 199248 163740 199300
rect 193220 199248 193272 199300
rect 108580 199044 108632 199096
rect 131580 199044 131632 199096
rect 115848 198976 115900 199028
rect 131764 198976 131816 199028
rect 132040 198976 132092 199028
rect 133512 199044 133564 199096
rect 135076 199044 135128 199096
rect 135720 199044 135772 199096
rect 135904 199044 135956 199096
rect 144828 199044 144880 199096
rect 154580 199044 154632 199096
rect 156420 199044 156472 199096
rect 156696 199044 156748 199096
rect 130016 198908 130068 198960
rect 132132 198908 132184 198960
rect 138296 198976 138348 199028
rect 147680 198976 147732 199028
rect 150716 198976 150768 199028
rect 157800 198976 157852 199028
rect 161664 199044 161716 199096
rect 190000 199180 190052 199232
rect 163964 199112 164016 199164
rect 189264 199112 189316 199164
rect 132868 198908 132920 198960
rect 135904 198908 135956 198960
rect 137008 198908 137060 198960
rect 139400 198908 139452 198960
rect 141424 198908 141476 198960
rect 121276 198840 121328 198892
rect 142160 198840 142212 198892
rect 142620 198908 142672 198960
rect 142988 198908 143040 198960
rect 143908 198908 143960 198960
rect 146300 198908 146352 198960
rect 152280 198908 152332 198960
rect 143172 198840 143224 198892
rect 160192 198908 160244 198960
rect 163228 198908 163280 198960
rect 190552 199044 190604 199096
rect 165344 198976 165396 199028
rect 168472 198976 168524 199028
rect 168656 198976 168708 199028
rect 200304 198976 200356 199028
rect 168288 198908 168340 198960
rect 171232 198908 171284 198960
rect 172060 198908 172112 198960
rect 172704 198908 172756 198960
rect 174268 198908 174320 198960
rect 178868 198908 178920 198960
rect 186596 198908 186648 198960
rect 126336 198772 126388 198824
rect 147864 198772 147916 198824
rect 154764 198772 154816 198824
rect 163964 198772 164016 198824
rect 168472 198772 168524 198824
rect 182824 198772 182876 198824
rect 126428 198704 126480 198756
rect 149060 198704 149112 198756
rect 157340 198704 157392 198756
rect 180064 198704 180116 198756
rect 184296 198704 184348 198756
rect 189172 198704 189224 198756
rect 129280 198636 129332 198688
rect 144092 198636 144144 198688
rect 154856 198636 154908 198688
rect 162492 198636 162544 198688
rect 164516 198636 164568 198688
rect 170680 198636 170732 198688
rect 170864 198636 170916 198688
rect 177856 198636 177908 198688
rect 129004 198568 129056 198620
rect 149336 198568 149388 198620
rect 157708 198568 157760 198620
rect 167092 198568 167144 198620
rect 170220 198568 170272 198620
rect 172612 198568 172664 198620
rect 211344 198568 211396 198620
rect 126520 198500 126572 198552
rect 147772 198500 147824 198552
rect 165528 198500 165580 198552
rect 172980 198500 173032 198552
rect 211528 198500 211580 198552
rect 122380 198432 122432 198484
rect 147128 198432 147180 198484
rect 159548 198432 159600 198484
rect 166264 198432 166316 198484
rect 168840 198432 168892 198484
rect 170864 198432 170916 198484
rect 170956 198432 171008 198484
rect 208860 198432 208912 198484
rect 125048 198364 125100 198416
rect 149428 198364 149480 198416
rect 159732 198364 159784 198416
rect 172060 198364 172112 198416
rect 173808 198364 173860 198416
rect 212724 198364 212776 198416
rect 122288 198296 122340 198348
rect 146852 198296 146904 198348
rect 105728 198228 105780 198280
rect 127532 198228 127584 198280
rect 107016 198160 107068 198212
rect 135996 198160 136048 198212
rect 141056 198160 141108 198212
rect 141516 198160 141568 198212
rect 151728 198160 151780 198212
rect 165712 198296 165764 198348
rect 167092 198296 167144 198348
rect 168104 198296 168156 198348
rect 171140 198296 171192 198348
rect 172612 198296 172664 198348
rect 173624 198296 173676 198348
rect 212908 198296 212960 198348
rect 163044 198228 163096 198280
rect 168840 198228 168892 198280
rect 170496 198228 170548 198280
rect 170956 198228 171008 198280
rect 172520 198228 172572 198280
rect 212632 198228 212684 198280
rect 159824 198160 159876 198212
rect 171140 198160 171192 198212
rect 174912 198160 174964 198212
rect 215484 198160 215536 198212
rect 108948 198092 109000 198144
rect 143356 198092 143408 198144
rect 148416 198092 148468 198144
rect 156236 198092 156288 198144
rect 163412 198092 163464 198144
rect 168104 198092 168156 198144
rect 170036 198092 170088 198144
rect 211804 198092 211856 198144
rect 103152 198024 103204 198076
rect 134064 198024 134116 198076
rect 149336 198024 149388 198076
rect 149888 198024 149940 198076
rect 155776 198024 155828 198076
rect 140780 197956 140832 198008
rect 145288 197956 145340 198008
rect 146208 197956 146260 198008
rect 159456 197956 159508 198008
rect 171508 198024 171560 198076
rect 171876 198024 171928 198076
rect 170496 197956 170548 198008
rect 176660 198024 176712 198076
rect 181168 198024 181220 198076
rect 181444 198024 181496 198076
rect 214380 198024 214432 198076
rect 124864 197888 124916 197940
rect 108396 197820 108448 197872
rect 142528 197820 142580 197872
rect 149612 197888 149664 197940
rect 149888 197888 149940 197940
rect 161572 197888 161624 197940
rect 211436 197956 211488 198008
rect 174176 197888 174228 197940
rect 187056 197888 187108 197940
rect 144644 197820 144696 197872
rect 149244 197820 149296 197872
rect 171048 197820 171100 197872
rect 124956 197752 125008 197804
rect 144460 197752 144512 197804
rect 149980 197752 150032 197804
rect 151084 197752 151136 197804
rect 160284 197752 160336 197804
rect 169760 197752 169812 197804
rect 171140 197752 171192 197804
rect 172152 197752 172204 197804
rect 160744 197684 160796 197736
rect 173808 197684 173860 197736
rect 176384 197684 176436 197736
rect 177672 197684 177724 197736
rect 129188 197616 129240 197668
rect 143632 197616 143684 197668
rect 157432 197616 157484 197668
rect 171876 197616 171928 197668
rect 181444 197820 181496 197872
rect 149796 197548 149848 197600
rect 150072 197548 150124 197600
rect 156052 197548 156104 197600
rect 149796 197412 149848 197464
rect 153936 197412 153988 197464
rect 133512 197344 133564 197396
rect 141332 197344 141384 197396
rect 156052 197344 156104 197396
rect 156604 197344 156656 197396
rect 167184 197548 167236 197600
rect 169760 197480 169812 197532
rect 175188 197480 175240 197532
rect 167828 197412 167880 197464
rect 168380 197412 168432 197464
rect 173900 197412 173952 197464
rect 174084 197412 174136 197464
rect 175372 197412 175424 197464
rect 176108 197412 176160 197464
rect 188344 197548 188396 197600
rect 177120 197344 177172 197396
rect 182456 197344 182508 197396
rect 105636 197276 105688 197328
rect 130292 197276 130344 197328
rect 131856 197276 131908 197328
rect 139492 197276 139544 197328
rect 139584 197276 139636 197328
rect 139952 197276 140004 197328
rect 141240 197276 141292 197328
rect 141884 197276 141936 197328
rect 166356 197276 166408 197328
rect 179420 197276 179472 197328
rect 121092 197208 121144 197260
rect 145840 197208 145892 197260
rect 157248 197208 157300 197260
rect 158996 197208 159048 197260
rect 160836 197208 160888 197260
rect 180432 197208 180484 197260
rect 108304 197140 108356 197192
rect 137376 197140 137428 197192
rect 137468 197140 137520 197192
rect 138112 197140 138164 197192
rect 139768 197140 139820 197192
rect 140044 197140 140096 197192
rect 141884 197140 141936 197192
rect 142344 197140 142396 197192
rect 160008 197140 160060 197192
rect 160652 197140 160704 197192
rect 162768 197140 162820 197192
rect 167920 197140 167972 197192
rect 168104 197140 168156 197192
rect 197360 197140 197412 197192
rect 119068 197072 119120 197124
rect 151820 197072 151872 197124
rect 164700 197072 164752 197124
rect 199660 197072 199712 197124
rect 112996 197004 113048 197056
rect 142068 197004 142120 197056
rect 171232 197004 171284 197056
rect 201684 197004 201736 197056
rect 111524 196936 111576 196988
rect 143264 196936 143316 196988
rect 154672 196936 154724 196988
rect 155408 196936 155460 196988
rect 159088 196936 159140 196988
rect 159916 196936 159968 196988
rect 164424 196936 164476 196988
rect 197544 196936 197596 196988
rect 112720 196868 112772 196920
rect 132868 196868 132920 196920
rect 137284 196868 137336 196920
rect 138388 196868 138440 196920
rect 139676 196868 139728 196920
rect 140504 196868 140556 196920
rect 143448 196868 143500 196920
rect 143816 196868 143868 196920
rect 155316 196868 155368 196920
rect 189172 196868 189224 196920
rect 114284 196800 114336 196852
rect 146116 196800 146168 196852
rect 160376 196800 160428 196852
rect 160560 196800 160612 196852
rect 161940 196800 161992 196852
rect 196348 196800 196400 196852
rect 111156 196732 111208 196784
rect 133144 196732 133196 196784
rect 139860 196732 139912 196784
rect 140320 196732 140372 196784
rect 164332 196732 164384 196784
rect 165344 196732 165396 196784
rect 172796 196732 172848 196784
rect 173348 196732 173400 196784
rect 175556 196732 175608 196784
rect 176476 196732 176528 196784
rect 177120 196732 177172 196784
rect 177396 196732 177448 196784
rect 181168 196732 181220 196784
rect 215300 196732 215352 196784
rect 105544 196664 105596 196716
rect 136640 196664 136692 196716
rect 138572 196664 138624 196716
rect 138848 196664 138900 196716
rect 139952 196664 140004 196716
rect 140412 196664 140464 196716
rect 141424 196664 141476 196716
rect 143724 196664 143776 196716
rect 148692 196664 148744 196716
rect 155500 196664 155552 196716
rect 157524 196664 157576 196716
rect 157708 196664 157760 196716
rect 160284 196664 160336 196716
rect 160928 196664 160980 196716
rect 161388 196664 161440 196716
rect 162768 196664 162820 196716
rect 164516 196664 164568 196716
rect 165620 196664 165672 196716
rect 165712 196664 165764 196716
rect 166724 196664 166776 196716
rect 167000 196664 167052 196716
rect 168196 196664 168248 196716
rect 168472 196664 168524 196716
rect 169300 196664 169352 196716
rect 169576 196664 169628 196716
rect 169852 196664 169904 196716
rect 172888 196664 172940 196716
rect 173532 196664 173584 196716
rect 177028 196664 177080 196716
rect 177580 196664 177632 196716
rect 181996 196664 182048 196716
rect 215668 196664 215720 196716
rect 97908 196596 97960 196648
rect 140872 196596 140924 196648
rect 141792 196596 141844 196648
rect 142988 196596 143040 196648
rect 143172 196596 143224 196648
rect 147220 196596 147272 196648
rect 151360 196596 151412 196648
rect 151820 196596 151872 196648
rect 152372 196596 152424 196648
rect 152648 196596 152700 196648
rect 152924 196596 152976 196648
rect 154764 196596 154816 196648
rect 155684 196596 155736 196648
rect 165988 196596 166040 196648
rect 166908 196596 166960 196648
rect 167644 196596 167696 196648
rect 170036 196596 170088 196648
rect 170128 196596 170180 196648
rect 216680 196596 216732 196648
rect 133512 196528 133564 196580
rect 149336 196528 149388 196580
rect 150256 196528 150308 196580
rect 154948 196528 155000 196580
rect 156604 196528 156656 196580
rect 176660 196528 176712 196580
rect 177212 196528 177264 196580
rect 177304 196528 177356 196580
rect 178224 196528 178276 196580
rect 126704 196460 126756 196512
rect 146576 196460 146628 196512
rect 164884 196460 164936 196512
rect 165436 196460 165488 196512
rect 169852 196460 169904 196512
rect 170220 196460 170272 196512
rect 175832 196460 175884 196512
rect 182272 196460 182324 196512
rect 129924 196392 129976 196444
rect 140596 196392 140648 196444
rect 162952 196392 163004 196444
rect 163228 196392 163280 196444
rect 169024 196392 169076 196444
rect 126612 196324 126664 196376
rect 148324 196324 148376 196376
rect 161940 196324 161992 196376
rect 162676 196324 162728 196376
rect 132868 196256 132920 196308
rect 144552 196256 144604 196308
rect 144920 196256 144972 196308
rect 145840 196256 145892 196308
rect 151912 196256 151964 196308
rect 153016 196256 153068 196308
rect 157984 196256 158036 196308
rect 159548 196256 159600 196308
rect 131028 196188 131080 196240
rect 134708 196188 134760 196240
rect 143908 196188 143960 196240
rect 144092 196188 144144 196240
rect 157800 196188 157852 196240
rect 158444 196188 158496 196240
rect 133144 196120 133196 196172
rect 144000 196120 144052 196172
rect 144920 196120 144972 196172
rect 146484 196120 146536 196172
rect 161756 196120 161808 196172
rect 168564 196120 168616 196172
rect 169392 196324 169444 196376
rect 183008 196324 183060 196376
rect 176936 196256 176988 196308
rect 177488 196256 177540 196308
rect 171048 196188 171100 196240
rect 178960 196188 179012 196240
rect 176844 196120 176896 196172
rect 177764 196120 177816 196172
rect 141608 196052 141660 196104
rect 143908 196052 143960 196104
rect 138480 195984 138532 196036
rect 138664 195984 138716 196036
rect 145472 195984 145524 196036
rect 146024 195984 146076 196036
rect 120724 195916 120776 195968
rect 145196 195916 145248 195968
rect 145380 195916 145432 195968
rect 146576 195916 146628 195968
rect 153476 195916 153528 195968
rect 153660 195916 153712 195968
rect 156236 195916 156288 195968
rect 157984 195916 158036 195968
rect 161664 195916 161716 195968
rect 169392 195916 169444 195968
rect 183100 195916 183152 195968
rect 123484 195848 123536 195900
rect 149152 195848 149204 195900
rect 157432 195848 157484 195900
rect 158076 195848 158128 195900
rect 158996 195848 159048 195900
rect 159272 195848 159324 195900
rect 161296 195848 161348 195900
rect 176200 195848 176252 195900
rect 119896 195780 119948 195832
rect 148968 195780 149020 195832
rect 153476 195780 153528 195832
rect 154304 195780 154356 195832
rect 156236 195780 156288 195832
rect 156512 195780 156564 195832
rect 175188 195780 175240 195832
rect 194600 195780 194652 195832
rect 118516 195712 118568 195764
rect 148140 195712 148192 195764
rect 150992 195712 151044 195764
rect 151636 195712 151688 195764
rect 173808 195712 173860 195764
rect 194692 195712 194744 195764
rect 117136 195644 117188 195696
rect 147864 195644 147916 195696
rect 172060 195644 172112 195696
rect 111340 195576 111392 195628
rect 128452 195576 128504 195628
rect 162492 195576 162544 195628
rect 173532 195576 173584 195628
rect 193404 195644 193456 195696
rect 182456 195576 182508 195628
rect 203616 195576 203668 195628
rect 115664 195508 115716 195560
rect 147312 195508 147364 195560
rect 158812 195508 158864 195560
rect 173716 195508 173768 195560
rect 179972 195508 180024 195560
rect 203708 195508 203760 195560
rect 104440 195440 104492 195492
rect 137652 195440 137704 195492
rect 138296 195440 138348 195492
rect 139032 195440 139084 195492
rect 154580 195440 154632 195492
rect 155040 195440 155092 195492
rect 157064 195440 157116 195492
rect 190460 195440 190512 195492
rect 104532 195372 104584 195424
rect 123392 195372 123444 195424
rect 123576 195372 123628 195424
rect 142804 195372 142856 195424
rect 109960 195304 110012 195356
rect 108856 195236 108908 195288
rect 143356 195236 143408 195288
rect 123576 195168 123628 195220
rect 128176 195168 128228 195220
rect 132132 195100 132184 195152
rect 149980 195372 150032 195424
rect 154488 195372 154540 195424
rect 187792 195372 187844 195424
rect 158720 195304 158772 195356
rect 192024 195304 192076 195356
rect 159364 195236 159416 195288
rect 218152 195236 218204 195288
rect 163136 195168 163188 195220
rect 164056 195168 164108 195220
rect 168932 195168 168984 195220
rect 183192 195168 183244 195220
rect 123392 195032 123444 195084
rect 137928 195032 137980 195084
rect 128452 194964 128504 195016
rect 163044 195100 163096 195152
rect 163780 195100 163832 195152
rect 165988 195100 166040 195152
rect 166448 195100 166500 195152
rect 173992 195100 174044 195152
rect 174728 195100 174780 195152
rect 176568 195100 176620 195152
rect 177212 195100 177264 195152
rect 155132 195032 155184 195084
rect 155684 195032 155736 195084
rect 175648 195032 175700 195084
rect 176384 195032 176436 195084
rect 148600 194964 148652 195016
rect 142896 194896 142948 194948
rect 155960 194896 156012 194948
rect 156788 194896 156840 194948
rect 165252 194896 165304 194948
rect 167184 194828 167236 194880
rect 167828 194828 167880 194880
rect 173716 194828 173768 194880
rect 176108 194828 176160 194880
rect 177580 194828 177632 194880
rect 132040 194760 132092 194812
rect 139216 194760 139268 194812
rect 176200 194760 176252 194812
rect 180340 194760 180392 194812
rect 183836 194692 183888 194744
rect 186504 194692 186556 194744
rect 174084 194556 174136 194608
rect 175004 194556 175056 194608
rect 130568 194488 130620 194540
rect 144920 194488 144972 194540
rect 130384 194420 130436 194472
rect 146760 194420 146812 194472
rect 130936 194352 130988 194404
rect 147588 194352 147640 194404
rect 156144 194352 156196 194404
rect 181444 194352 181496 194404
rect 127808 194284 127860 194336
rect 144644 194284 144696 194336
rect 153384 194284 153436 194336
rect 181536 194284 181588 194336
rect 127992 194216 128044 194268
rect 148048 194216 148100 194268
rect 176292 194216 176344 194268
rect 209964 194216 210016 194268
rect 122196 194148 122248 194200
rect 143540 194148 143592 194200
rect 173808 194148 173860 194200
rect 207296 194148 207348 194200
rect 108488 194080 108540 194132
rect 140780 194080 140832 194132
rect 170864 194080 170916 194132
rect 203064 194080 203116 194132
rect 108672 194012 108724 194064
rect 139124 194012 139176 194064
rect 174360 194012 174412 194064
rect 208768 194012 208820 194064
rect 113916 193944 113968 193996
rect 145564 193944 145616 193996
rect 153292 193944 153344 193996
rect 154028 193944 154080 193996
rect 173440 193944 173492 193996
rect 207572 193944 207624 193996
rect 111432 193876 111484 193928
rect 145656 193876 145708 193928
rect 173624 193876 173676 193928
rect 207664 193876 207716 193928
rect 111248 193808 111300 193860
rect 145012 193808 145064 193860
rect 166816 193808 166868 193860
rect 213092 193808 213144 193860
rect 130752 193740 130804 193792
rect 147496 193740 147548 193792
rect 130568 193672 130620 193724
rect 144092 193672 144144 193724
rect 174268 193672 174320 193724
rect 174820 193672 174872 193724
rect 130844 193604 130896 193656
rect 145104 193604 145156 193656
rect 141700 193536 141752 193588
rect 143632 193536 143684 193588
rect 149704 193536 149756 193588
rect 150440 193536 150492 193588
rect 150624 193128 150676 193180
rect 151544 193128 151596 193180
rect 189816 193128 189868 193180
rect 580172 193128 580224 193180
rect 107108 193060 107160 193112
rect 130016 193060 130068 193112
rect 162124 193060 162176 193112
rect 162676 193060 162728 193112
rect 174452 193060 174504 193112
rect 175096 193060 175148 193112
rect 179420 193060 179472 193112
rect 198924 193060 198976 193112
rect 105820 192992 105872 193044
rect 129924 192992 129976 193044
rect 138480 192992 138532 193044
rect 139308 192992 139360 193044
rect 171600 192992 171652 193044
rect 204720 192992 204772 193044
rect 122472 192924 122524 192976
rect 147220 192924 147272 192976
rect 157524 192924 157576 192976
rect 158352 192924 158404 192976
rect 178040 192924 178092 192976
rect 205916 192924 205968 192976
rect 100484 192856 100536 192908
rect 128544 192856 128596 192908
rect 170772 192856 170824 192908
rect 204536 192856 204588 192908
rect 110328 192788 110380 192840
rect 144368 192788 144420 192840
rect 173164 192788 173216 192840
rect 206008 192788 206060 192840
rect 110144 192720 110196 192772
rect 144184 192720 144236 192772
rect 150532 192720 150584 192772
rect 185676 192720 185728 192772
rect 123944 192652 123996 192704
rect 161848 192652 161900 192704
rect 170220 192652 170272 192704
rect 204904 192652 204956 192704
rect 108764 192584 108816 192636
rect 143080 192584 143132 192636
rect 156880 192584 156932 192636
rect 210332 192584 210384 192636
rect 104348 192516 104400 192568
rect 138020 192516 138072 192568
rect 155868 192516 155920 192568
rect 209780 192516 209832 192568
rect 110052 192448 110104 192500
rect 143540 192448 143592 192500
rect 155224 192448 155276 192500
rect 211160 192448 211212 192500
rect 161848 192380 161900 192432
rect 162400 192380 162452 192432
rect 168380 192108 168432 192160
rect 169668 192108 169720 192160
rect 158628 192040 158680 192092
rect 160652 192040 160704 192092
rect 171324 192040 171376 192092
rect 205732 192040 205784 192092
rect 170680 191972 170732 192024
rect 204352 191972 204404 192024
rect 171968 191904 172020 191956
rect 206100 191904 206152 191956
rect 170956 191836 171008 191888
rect 204812 191836 204864 191888
rect 171324 191768 171376 191820
rect 172244 191768 172296 191820
rect 132592 191700 132644 191752
rect 133420 191700 133472 191752
rect 130292 191632 130344 191684
rect 132500 191632 132552 191684
rect 131028 191564 131080 191616
rect 135260 191564 135312 191616
rect 166264 191564 166316 191616
rect 185860 191564 185912 191616
rect 132224 191496 132276 191548
rect 139584 191496 139636 191548
rect 164148 191496 164200 191548
rect 184204 191496 184256 191548
rect 122564 191428 122616 191480
rect 141240 191428 141292 191480
rect 162676 191428 162728 191480
rect 185768 191428 185820 191480
rect 123852 191360 123904 191412
rect 154580 191360 154632 191412
rect 163596 191360 163648 191412
rect 164148 191360 164200 191412
rect 167644 191360 167696 191412
rect 201500 191360 201552 191412
rect 103336 191292 103388 191344
rect 131028 191292 131080 191344
rect 167460 191292 167512 191344
rect 201776 191292 201828 191344
rect 99196 191224 99248 191276
rect 130292 191224 130344 191276
rect 100392 191156 100444 191208
rect 133972 191224 134024 191276
rect 168656 191224 168708 191276
rect 202972 191224 203024 191276
rect 134064 191156 134116 191208
rect 134524 191156 134576 191208
rect 135720 191156 135772 191208
rect 136272 191156 136324 191208
rect 137100 191156 137152 191208
rect 137560 191156 137612 191208
rect 161204 191156 161256 191208
rect 216772 191156 216824 191208
rect 103060 191088 103112 191140
rect 143448 191088 143500 191140
rect 152188 191088 152240 191140
rect 218336 191088 218388 191140
rect 134156 191020 134208 191072
rect 135168 191020 135220 191072
rect 135536 191020 135588 191072
rect 136456 191020 136508 191072
rect 149888 190952 149940 191004
rect 150164 190952 150216 191004
rect 121828 190408 121880 190460
rect 149980 190408 150032 190460
rect 177212 190408 177264 190460
rect 210424 190408 210476 190460
rect 107384 190340 107436 190392
rect 138664 190340 138716 190392
rect 177304 190340 177356 190392
rect 211712 190340 211764 190392
rect 106188 190272 106240 190324
rect 130292 190272 130344 190324
rect 130660 190272 130712 190324
rect 130936 190272 130988 190324
rect 175556 190272 175608 190324
rect 210056 190272 210108 190324
rect 104256 190204 104308 190256
rect 136364 190204 136416 190256
rect 172888 190204 172940 190256
rect 207480 190204 207532 190256
rect 100576 190136 100628 190188
rect 132316 190136 132368 190188
rect 160560 190136 160612 190188
rect 195152 190136 195204 190188
rect 103428 190068 103480 190120
rect 135628 190068 135680 190120
rect 174268 190068 174320 190120
rect 208952 190068 209004 190120
rect 111616 190000 111668 190052
rect 144736 190000 144788 190052
rect 164700 190000 164752 190052
rect 205824 190000 205876 190052
rect 104624 189932 104676 189984
rect 102876 189864 102928 189916
rect 130108 189864 130160 189916
rect 130292 189932 130344 189984
rect 137744 189932 137796 189984
rect 163504 189932 163556 189984
rect 214288 189932 214340 189984
rect 137284 189864 137336 189916
rect 159180 189864 159232 189916
rect 216956 189864 217008 189916
rect 102968 189796 103020 189848
rect 136916 189796 136968 189848
rect 155408 189796 155460 189848
rect 218244 189796 218296 189848
rect 101588 189728 101640 189780
rect 136088 189728 136140 189780
rect 154396 189728 154448 189780
rect 218428 189728 218480 189780
rect 130108 189660 130160 189712
rect 137468 189660 137520 189712
rect 174452 189660 174504 189712
rect 207388 189660 207440 189712
rect 156328 189592 156380 189644
rect 187424 189592 187476 189644
rect 160468 189524 160520 189576
rect 185584 189524 185636 189576
rect 3424 188980 3476 189032
rect 117780 188980 117832 189032
rect 166080 187552 166132 187604
rect 200396 187552 200448 187604
rect 161848 187484 161900 187536
rect 209044 187484 209096 187536
rect 160008 187416 160060 187468
rect 207020 187416 207072 187468
rect 159088 187348 159140 187400
rect 207112 187348 207164 187400
rect 161940 187280 161992 187332
rect 210148 187280 210200 187332
rect 101496 187212 101548 187264
rect 134984 187212 135036 187264
rect 154764 187212 154816 187264
rect 214196 187212 214248 187264
rect 99104 187144 99156 187196
rect 133604 187144 133656 187196
rect 152832 187144 152884 187196
rect 214104 187144 214156 187196
rect 99288 187076 99340 187128
rect 132776 187076 132828 187128
rect 149336 187076 149388 187128
rect 211620 187076 211672 187128
rect 99012 187008 99064 187060
rect 133236 187008 133288 187060
rect 151084 187008 151136 187060
rect 215760 187008 215812 187060
rect 100208 186940 100260 186992
rect 134340 186940 134392 186992
rect 150808 186940 150860 186992
rect 218520 186940 218572 186992
rect 188528 178032 188580 178084
rect 580172 178032 580224 178084
rect 189816 165588 189868 165640
rect 580172 165588 580224 165640
rect 168748 158380 168800 158432
rect 189724 158380 189776 158432
rect 172888 158312 172940 158364
rect 201960 158312 202012 158364
rect 170036 158244 170088 158296
rect 203248 158244 203300 158296
rect 166080 158176 166132 158228
rect 203156 158176 203208 158228
rect 159732 158108 159784 158160
rect 214472 158108 214524 158160
rect 152096 158040 152148 158092
rect 213184 158040 213236 158092
rect 152188 157972 152240 158024
rect 217140 157972 217192 158024
rect 171508 155864 171560 155916
rect 201868 155864 201920 155916
rect 170220 155796 170272 155848
rect 191012 155796 191064 155848
rect 167276 155728 167328 155780
rect 201868 155728 201920 155780
rect 167552 155660 167604 155712
rect 202236 155660 202288 155712
rect 165988 155592 166040 155644
rect 200764 155592 200816 155644
rect 165896 155524 165948 155576
rect 200672 155524 200724 155576
rect 167368 155456 167420 155508
rect 202144 155456 202196 155508
rect 177028 155388 177080 155440
rect 211896 155388 211948 155440
rect 168564 155320 168616 155372
rect 203432 155320 203484 155372
rect 168656 155252 168708 155304
rect 203524 155252 203576 155304
rect 168288 155184 168340 155236
rect 202328 155184 202380 155236
rect 174268 155116 174320 155168
rect 193864 155116 193916 155168
rect 183560 154504 183612 154556
rect 184296 154504 184348 154556
rect 112444 154368 112496 154420
rect 132684 154368 132736 154420
rect 116584 154300 116636 154352
rect 143540 154300 143592 154352
rect 113732 154232 113784 154284
rect 141240 154232 141292 154284
rect 115112 154164 115164 154216
rect 146392 154164 146444 154216
rect 101220 154096 101272 154148
rect 134156 154096 134208 154148
rect 98920 154028 98972 154080
rect 133328 154028 133380 154080
rect 100024 153960 100076 154012
rect 134340 153960 134392 154012
rect 100116 153892 100168 153944
rect 134432 153892 134484 153944
rect 99932 153824 99984 153876
rect 134064 153824 134116 153876
rect 97264 153212 97316 153264
rect 183560 153212 183612 153264
rect 160376 153144 160428 153196
rect 184664 153144 184716 153196
rect 161664 153076 161716 153128
rect 185952 153076 186004 153128
rect 161756 153008 161808 153060
rect 186136 153008 186188 153060
rect 158904 152940 158956 152992
rect 184572 152940 184624 152992
rect 158996 152872 159048 152924
rect 185492 152872 185544 152924
rect 157800 152804 157852 152856
rect 184388 152804 184440 152856
rect 157708 152736 157760 152788
rect 184480 152736 184532 152788
rect 178960 152668 179012 152720
rect 210516 152668 210568 152720
rect 176844 152600 176896 152652
rect 210608 152600 210660 152652
rect 166908 152532 166960 152584
rect 200580 152532 200632 152584
rect 176936 152464 176988 152516
rect 211988 152464 212040 152516
rect 165712 152396 165764 152448
rect 186228 152396 186280 152448
rect 165252 152328 165304 152380
rect 184296 152328 184348 152380
rect 188436 151784 188488 151836
rect 579988 151784 580040 151836
rect 115112 151648 115164 151700
rect 141148 151648 141200 151700
rect 113548 151580 113600 151632
rect 142988 151580 143040 151632
rect 168472 151580 168524 151632
rect 186780 151580 186832 151632
rect 111984 151512 112036 151564
rect 142436 151512 142488 151564
rect 157616 151512 157668 151564
rect 188712 151512 188764 151564
rect 106832 151444 106884 151496
rect 138204 151444 138256 151496
rect 156236 151444 156288 151496
rect 187240 151444 187292 151496
rect 109592 151376 109644 151428
rect 140964 151376 141016 151428
rect 162768 151376 162820 151428
rect 198464 151376 198516 151428
rect 104164 151308 104216 151360
rect 137192 151308 137244 151360
rect 163320 151308 163372 151360
rect 204996 151308 205048 151360
rect 99840 151240 99892 151292
rect 132592 151240 132644 151292
rect 163412 151240 163464 151292
rect 207848 151240 207900 151292
rect 106740 151172 106792 151224
rect 139676 151172 139728 151224
rect 154764 151172 154816 151224
rect 204444 151172 204496 151224
rect 102600 151104 102652 151156
rect 135536 151104 135588 151156
rect 150624 151104 150676 151156
rect 209136 151104 209188 151156
rect 104072 151036 104124 151088
rect 138296 151036 138348 151088
rect 154672 151036 154724 151088
rect 217232 151036 217284 151088
rect 124772 150424 124824 150476
rect 125140 150424 125192 150476
rect 580448 150424 580500 150476
rect 176752 150356 176804 150408
rect 207756 150356 207808 150408
rect 182088 150016 182140 150068
rect 198004 150016 198056 150068
rect 172796 149948 172848 150000
rect 203800 149948 203852 150000
rect 175372 149880 175424 149932
rect 206468 149880 206520 149932
rect 112168 149812 112220 149864
rect 141792 149812 141844 149864
rect 174084 149812 174136 149864
rect 206284 149812 206336 149864
rect 102692 149744 102744 149796
rect 135812 149744 135864 149796
rect 173992 149744 174044 149796
rect 206376 149744 206428 149796
rect 101312 149676 101364 149728
rect 135904 149676 135956 149728
rect 172704 149676 172756 149728
rect 205088 149676 205140 149728
rect 3148 149132 3200 149184
rect 180892 149132 180944 149184
rect 182088 149132 182140 149184
rect 119252 149064 119304 149116
rect 119988 149064 120040 149116
rect 580264 149064 580316 149116
rect 122564 148996 122616 149048
rect 149796 148996 149848 149048
rect 160284 148996 160336 149048
rect 186964 148996 187016 149048
rect 203616 148996 203668 149048
rect 203800 148996 203852 149048
rect 113824 148928 113876 148980
rect 125140 148928 125192 148980
rect 158812 148928 158864 148980
rect 188620 148928 188672 148980
rect 115204 148860 115256 148912
rect 128360 148860 128412 148912
rect 157524 148860 157576 148912
rect 188160 148860 188212 148912
rect 116952 148792 117004 148844
rect 142528 148792 142580 148844
rect 161572 148792 161624 148844
rect 194784 148792 194836 148844
rect 122104 148724 122156 148776
rect 149704 148724 149756 148776
rect 163228 148724 163280 148776
rect 198372 148724 198424 148776
rect 112076 148656 112128 148708
rect 142712 148656 142764 148708
rect 163136 148656 163188 148708
rect 198280 148656 198332 148708
rect 114928 148588 114980 148640
rect 145472 148588 145524 148640
rect 164608 148588 164660 148640
rect 199844 148588 199896 148640
rect 115572 148520 115624 148572
rect 145564 148520 145616 148572
rect 157156 148520 157208 148572
rect 191012 148520 191064 148572
rect 116308 148452 116360 148504
rect 146668 148452 146720 148504
rect 164424 148452 164476 148504
rect 199384 148452 199436 148504
rect 112536 148384 112588 148436
rect 145196 148384 145248 148436
rect 158628 148384 158680 148436
rect 196992 148384 197044 148436
rect 98828 148316 98880 148368
rect 132960 148316 133012 148368
rect 155684 148316 155736 148368
rect 217048 148316 217100 148368
rect 164516 148248 164568 148300
rect 191104 148248 191156 148300
rect 177580 148180 177632 148232
rect 199936 148180 199988 148232
rect 180432 148112 180484 148164
rect 193956 148112 194008 148164
rect 128360 147636 128412 147688
rect 128636 147636 128688 147688
rect 136180 147636 136232 147688
rect 169852 147568 169904 147620
rect 196440 147568 196492 147620
rect 172612 147500 172664 147552
rect 198740 147500 198792 147552
rect 117688 147432 117740 147484
rect 132132 147432 132184 147484
rect 171232 147432 171284 147484
rect 180432 147432 180484 147484
rect 113732 147364 113784 147416
rect 130752 147364 130804 147416
rect 179604 147364 179656 147416
rect 197728 147364 197780 147416
rect 111892 147296 111944 147348
rect 130844 147296 130896 147348
rect 179696 147296 179748 147348
rect 199200 147296 199252 147348
rect 109684 147228 109736 147280
rect 132040 147228 132092 147280
rect 116216 147160 116268 147212
rect 143724 147160 143776 147212
rect 156236 147160 156288 147212
rect 113824 147092 113876 147144
rect 143908 147092 143960 147144
rect 178960 147228 179012 147280
rect 197912 147228 197964 147280
rect 179512 147160 179564 147212
rect 199108 147160 199160 147212
rect 180248 147092 180300 147144
rect 110788 147024 110840 147076
rect 143632 147024 143684 147076
rect 171416 147024 171468 147076
rect 198096 147092 198148 147144
rect 180432 147024 180484 147076
rect 198188 147024 198240 147076
rect 109776 146956 109828 147008
rect 143816 146956 143868 147008
rect 157248 146956 157300 147008
rect 193864 146956 193916 147008
rect 109500 146888 109552 146940
rect 145288 146888 145340 146940
rect 146208 146888 146260 146940
rect 184756 146888 184808 146940
rect 185860 146888 185912 146940
rect 186044 146888 186096 146940
rect 185676 146752 185728 146804
rect 186044 146752 186096 146804
rect 176108 146208 176160 146260
rect 194140 146208 194192 146260
rect 120356 146140 120408 146192
rect 131764 146140 131816 146192
rect 178408 146140 178460 146192
rect 196716 146140 196768 146192
rect 117964 146072 118016 146124
rect 129740 146072 129792 146124
rect 177212 146072 177264 146124
rect 199292 146072 199344 146124
rect 115388 146004 115440 146056
rect 131304 146004 131356 146056
rect 157524 146004 157576 146056
rect 188436 146004 188488 146056
rect 114008 145936 114060 145988
rect 130292 145936 130344 145988
rect 159916 145936 159968 145988
rect 192852 145936 192904 145988
rect 111064 145868 111116 145920
rect 126980 145868 127032 145920
rect 161296 145868 161348 145920
rect 194232 145868 194284 145920
rect 120632 145800 120684 145852
rect 143632 145800 143684 145852
rect 155960 145800 156012 145852
rect 189448 145800 189500 145852
rect 117964 145732 118016 145784
rect 146576 145732 146628 145784
rect 160192 145732 160244 145784
rect 195520 145732 195572 145784
rect 115204 145664 115256 145716
rect 148232 145664 148284 145716
rect 162308 145664 162360 145716
rect 196532 145664 196584 145716
rect 112812 145596 112864 145648
rect 145012 145596 145064 145648
rect 156052 145596 156104 145648
rect 191196 145596 191248 145648
rect 3516 145528 3568 145580
rect 183468 145528 183520 145580
rect 197820 145528 197872 145580
rect 178316 145460 178368 145512
rect 195980 145460 196032 145512
rect 178224 145392 178276 145444
rect 193772 145392 193824 145444
rect 179788 145324 179840 145376
rect 192668 145324 192720 145376
rect 118792 144916 118844 144968
rect 182272 144916 182324 144968
rect 183468 144916 183520 144968
rect 116676 144848 116728 144900
rect 133880 144848 133932 144900
rect 184112 144848 184164 144900
rect 196808 144848 196860 144900
rect 112444 144780 112496 144832
rect 130568 144780 130620 144832
rect 177120 144780 177172 144832
rect 195060 144780 195112 144832
rect 119528 144712 119580 144764
rect 138112 144712 138164 144764
rect 172336 144712 172388 144764
rect 185676 144712 185728 144764
rect 115480 144644 115532 144696
rect 135444 144644 135496 144696
rect 172428 144644 172480 144696
rect 196624 144644 196676 144696
rect 120264 144576 120316 144628
rect 150072 144576 150124 144628
rect 165528 144576 165580 144628
rect 193588 144576 193640 144628
rect 118884 144508 118936 144560
rect 151820 144508 151872 144560
rect 163964 144508 164016 144560
rect 192484 144508 192536 144560
rect 119620 144440 119672 144492
rect 152464 144440 152516 144492
rect 154488 144440 154540 144492
rect 187976 144440 188028 144492
rect 117872 144372 117924 144424
rect 151912 144372 151964 144424
rect 157800 144372 157852 144424
rect 192392 144372 192444 144424
rect 103980 144304 104032 144356
rect 145748 144304 145800 144356
rect 159548 144304 159600 144356
rect 193680 144304 193732 144356
rect 112628 144236 112680 144288
rect 131212 144236 131264 144288
rect 188528 144236 188580 144288
rect 116860 144168 116912 144220
rect 130200 144168 130252 144220
rect 189816 144168 189868 144220
rect 113640 144100 113692 144152
rect 130476 144100 130528 144152
rect 185676 144100 185728 144152
rect 192944 144100 192996 144152
rect 112352 144032 112404 144084
rect 122656 144032 122708 144084
rect 117596 143964 117648 144016
rect 128176 143964 128228 144016
rect 125232 143556 125284 143608
rect 126244 143556 126296 143608
rect 580540 143556 580592 143608
rect 118240 143488 118292 143540
rect 128452 143488 128504 143540
rect 147680 143488 147732 143540
rect 150808 143488 150860 143540
rect 170036 143488 170088 143540
rect 170312 143488 170364 143540
rect 172888 143488 172940 143540
rect 173532 143488 173584 143540
rect 174268 143488 174320 143540
rect 179696 143488 179748 143540
rect 185768 143488 185820 143540
rect 189356 143488 189408 143540
rect 118332 143352 118384 143404
rect 131488 143420 131540 143472
rect 176292 143420 176344 143472
rect 179604 143420 179656 143472
rect 181536 143420 181588 143472
rect 187976 143420 188028 143472
rect 188068 143420 188120 143472
rect 191380 143420 191432 143472
rect 115296 143216 115348 143268
rect 130384 143352 130436 143404
rect 131120 143352 131172 143404
rect 137560 143352 137612 143404
rect 175740 143352 175792 143404
rect 178316 143352 178368 143404
rect 178868 143352 178920 143404
rect 190276 143352 190328 143404
rect 121000 143284 121052 143336
rect 134800 143284 134852 143336
rect 170956 143284 171008 143336
rect 179512 143284 179564 143336
rect 181720 143284 181772 143336
rect 193496 143284 193548 143336
rect 129740 143216 129792 143268
rect 137008 143216 137060 143268
rect 169668 143216 169720 143268
rect 179420 143216 179472 143268
rect 184296 143216 184348 143268
rect 196440 143216 196492 143268
rect 116768 143148 116820 143200
rect 133144 143148 133196 143200
rect 173164 143148 173216 143200
rect 190644 143148 190696 143200
rect 120908 143080 120960 143132
rect 139768 143080 139820 143132
rect 168196 143080 168248 143132
rect 181352 143080 181404 143132
rect 181444 143080 181496 143132
rect 188068 143080 188120 143132
rect 119712 143012 119764 143064
rect 141424 143012 141476 143064
rect 166632 143012 166684 143064
rect 190920 143012 190972 143064
rect 119344 142944 119396 142996
rect 144920 142944 144972 142996
rect 154304 142944 154356 142996
rect 188252 142944 188304 142996
rect 119436 142876 119488 142928
rect 148048 142876 148100 142928
rect 168380 142876 168432 142928
rect 209228 142876 209280 142928
rect 116860 142808 116912 142860
rect 149704 142808 149756 142860
rect 155500 142808 155552 142860
rect 207848 142808 207900 142860
rect 186044 142740 186096 142792
rect 192668 142740 192720 142792
rect 181352 142672 181404 142724
rect 189540 142672 189592 142724
rect 188068 142604 188120 142656
rect 188712 142604 188764 142656
rect 127532 142400 127584 142452
rect 127808 142400 127860 142452
rect 123116 142332 123168 142384
rect 123944 142332 123996 142384
rect 126060 142332 126112 142384
rect 126428 142332 126480 142384
rect 40684 142264 40736 142316
rect 184296 142264 184348 142316
rect 121000 142196 121052 142248
rect 146392 142196 146444 142248
rect 184020 142196 184072 142248
rect 192576 142196 192628 142248
rect 129832 142128 129884 142180
rect 134248 142128 134300 142180
rect 117044 142060 117096 142112
rect 118056 141992 118108 142044
rect 123484 141992 123536 142044
rect 125600 142060 125652 142112
rect 150532 142128 150584 142180
rect 155868 142128 155920 142180
rect 157340 142128 157392 142180
rect 159180 142128 159232 142180
rect 192208 142060 192260 142112
rect 126520 141992 126572 142044
rect 184112 141992 184164 142044
rect 184388 141992 184440 142044
rect 184480 141992 184532 142044
rect 184848 141992 184900 142044
rect 186136 141992 186188 142044
rect 196624 141992 196676 142044
rect 114100 141924 114152 141976
rect 125600 141924 125652 141976
rect 186228 141924 186280 141976
rect 186872 141924 186924 141976
rect 187148 141924 187200 141976
rect 196716 141924 196768 141976
rect 114192 141856 114244 141908
rect 127072 141856 127124 141908
rect 180340 141856 180392 141908
rect 194968 141856 195020 141908
rect 112904 141788 112956 141840
rect 129280 141788 129332 141840
rect 176476 141788 176528 141840
rect 192300 141788 192352 141840
rect 118148 141720 118200 141772
rect 140320 141720 140372 141772
rect 170496 141720 170548 141772
rect 185308 141720 185360 141772
rect 185952 141720 186004 141772
rect 187148 141720 187200 141772
rect 123484 141652 123536 141704
rect 136640 141652 136692 141704
rect 180156 141652 180208 141704
rect 199292 141652 199344 141704
rect 113088 141584 113140 141636
rect 139400 141584 139452 141636
rect 164240 141584 164292 141636
rect 187332 141584 187384 141636
rect 119804 141516 119856 141568
rect 153752 141516 153804 141568
rect 167460 141516 167512 141568
rect 192116 141516 192168 141568
rect 119252 141448 119304 141500
rect 158076 141448 158128 141500
rect 166448 141448 166500 141500
rect 217324 141448 217376 141500
rect 119620 141380 119672 141432
rect 149888 141380 149940 141432
rect 151268 141380 151320 141432
rect 214564 141380 214616 141432
rect 116584 141312 116636 141364
rect 119988 141312 120040 141364
rect 123208 141312 123260 141364
rect 184756 141312 184808 141364
rect 195060 141312 195112 141364
rect 127992 141244 128044 141296
rect 184664 141244 184716 141296
rect 194968 141244 195020 141296
rect 185308 141176 185360 141228
rect 189816 141176 189868 141228
rect 117044 140972 117096 141024
rect 124956 140972 125008 141024
rect 116400 140904 116452 140956
rect 123300 140904 123352 140956
rect 123392 140904 123444 140956
rect 142252 140904 142304 140956
rect 97356 140836 97408 140888
rect 181720 140836 181772 140888
rect 13084 140768 13136 140820
rect 182916 140768 182968 140820
rect 120816 140700 120868 140752
rect 126612 140700 126664 140752
rect 131304 140700 131356 140752
rect 132040 140700 132092 140752
rect 145012 140700 145064 140752
rect 145840 140700 145892 140752
rect 183560 140700 183612 140752
rect 184480 140700 184532 140752
rect 120540 140632 120592 140684
rect 126428 140632 126480 140684
rect 184204 140632 184256 140684
rect 192392 140632 192444 140684
rect 118148 140564 118200 140616
rect 121736 140564 121788 140616
rect 121920 140564 121972 140616
rect 125048 140564 125100 140616
rect 184848 140564 184900 140616
rect 192300 140564 192352 140616
rect 118056 140496 118108 140548
rect 115388 140360 115440 140412
rect 118332 140360 118384 140412
rect 119804 140496 119856 140548
rect 126152 140496 126204 140548
rect 185584 140496 185636 140548
rect 195336 140496 195388 140548
rect 119160 140428 119212 140480
rect 126704 140428 126756 140480
rect 180064 140428 180116 140480
rect 190644 140428 190696 140480
rect 126336 140360 126388 140412
rect 178776 140360 178828 140412
rect 190828 140360 190880 140412
rect 125508 140292 125560 140344
rect 138388 140292 138440 140344
rect 178684 140292 178736 140344
rect 190736 140292 190788 140344
rect 115020 140224 115072 140276
rect 112260 140156 112312 140208
rect 117044 140156 117096 140208
rect 129004 140224 129056 140276
rect 164148 140224 164200 140276
rect 187148 140224 187200 140276
rect 124496 140156 124548 140208
rect 139676 140156 139728 140208
rect 162952 140156 163004 140208
rect 197912 140156 197964 140208
rect 119712 140088 119764 140140
rect 150992 140088 151044 140140
rect 157432 140088 157484 140140
rect 192576 140088 192628 140140
rect 121736 140020 121788 140072
rect 126060 140020 126112 140072
rect 118332 139952 118384 140004
rect 127624 139952 127676 140004
rect 116860 139884 116912 139936
rect 148140 140020 148192 140072
rect 156788 140020 156840 140072
rect 197820 140020 197872 140072
rect 172980 139680 173032 139732
rect 197636 139680 197688 139732
rect 161296 139612 161348 139664
rect 194876 139612 194928 139664
rect 123392 139544 123444 139596
rect 183560 139544 183612 139596
rect 118700 139476 118752 139528
rect 180064 139476 180116 139528
rect 183284 139476 183336 139528
rect 189632 139476 189684 139528
rect 125876 139408 125928 139460
rect 327724 139408 327776 139460
rect 188620 139204 188672 139256
rect 189724 139204 189776 139256
rect 189908 138660 189960 138712
rect 195244 138660 195296 138712
rect 3424 137980 3476 138032
rect 121000 137980 121052 138032
rect 3240 137912 3292 137964
rect 118700 137912 118752 137964
rect 120264 137300 120316 137352
rect 120632 137300 120684 137352
rect 117872 136144 117924 136196
rect 119804 136144 119856 136196
rect 3056 111392 3108 111444
rect 8944 111392 8996 111444
rect 467104 100648 467156 100700
rect 580172 100648 580224 100700
rect 188988 99356 189040 99408
rect 189816 99356 189868 99408
rect 190368 98200 190420 98252
rect 192668 98200 192720 98252
rect 188896 92488 188948 92540
rect 191840 92488 191892 92540
rect 464344 86912 464396 86964
rect 579988 86912 580040 86964
rect 3516 85484 3568 85536
rect 97356 85484 97408 85536
rect 186964 81472 187016 81524
rect 187424 81472 187476 81524
rect 186688 81404 186740 81456
rect 187516 81404 187568 81456
rect 112352 81064 112404 81116
rect 121828 81064 121880 81116
rect 122288 80996 122340 81048
rect 114928 80928 114980 80980
rect 117964 80860 118016 80912
rect 113916 80792 113968 80844
rect 112260 80724 112312 80776
rect 113640 80656 113692 80708
rect 121828 80588 121880 80640
rect 125600 80588 125652 80640
rect 105268 80520 105320 80572
rect 105636 80520 105688 80572
rect 130476 80588 130528 80640
rect 131120 80588 131172 80640
rect 131304 80588 131356 80640
rect 130476 80384 130528 80436
rect 130384 80316 130436 80368
rect 129004 80044 129056 80096
rect 132546 79908 132598 79960
rect 132730 79908 132782 79960
rect 132822 79908 132874 79960
rect 132914 79908 132966 79960
rect 133006 79908 133058 79960
rect 133374 79908 133426 79960
rect 133466 79908 133518 79960
rect 132500 79772 132552 79824
rect 113732 79636 113784 79688
rect 130384 79636 130436 79688
rect 133098 79840 133150 79892
rect 132776 79704 132828 79756
rect 132868 79704 132920 79756
rect 132960 79704 133012 79756
rect 133144 79704 133196 79756
rect 134386 79908 134438 79960
rect 134570 79908 134622 79960
rect 133328 79636 133380 79688
rect 133742 79840 133794 79892
rect 133834 79840 133886 79892
rect 133926 79840 133978 79892
rect 134018 79840 134070 79892
rect 109868 79568 109920 79620
rect 130292 79568 130344 79620
rect 132684 79568 132736 79620
rect 119252 79500 119304 79552
rect 130568 79500 130620 79552
rect 111156 79432 111208 79484
rect 131028 79432 131080 79484
rect 108212 79364 108264 79416
rect 129924 79364 129976 79416
rect 132868 79432 132920 79484
rect 133880 79704 133932 79756
rect 134478 79840 134530 79892
rect 134524 79704 134576 79756
rect 134064 79636 134116 79688
rect 134248 79636 134300 79688
rect 134340 79636 134392 79688
rect 133972 79500 134024 79552
rect 134708 79500 134760 79552
rect 135030 79908 135082 79960
rect 135122 79908 135174 79960
rect 135076 79704 135128 79756
rect 135398 79908 135450 79960
rect 135582 79908 135634 79960
rect 135766 79908 135818 79960
rect 135858 79908 135910 79960
rect 136042 79908 136094 79960
rect 136410 79908 136462 79960
rect 136594 79908 136646 79960
rect 136778 79908 136830 79960
rect 137146 79908 137198 79960
rect 137238 79908 137290 79960
rect 137422 79908 137474 79960
rect 137514 79908 137566 79960
rect 135260 79568 135312 79620
rect 135720 79772 135772 79824
rect 136318 79772 136370 79824
rect 135812 79704 135864 79756
rect 135352 79500 135404 79552
rect 135628 79500 135680 79552
rect 135904 79568 135956 79620
rect 136548 79636 136600 79688
rect 136732 79636 136784 79688
rect 136962 79840 137014 79892
rect 137100 79704 137152 79756
rect 137376 79772 137428 79824
rect 137606 79840 137658 79892
rect 137468 79704 137520 79756
rect 137192 79636 137244 79688
rect 138066 79908 138118 79960
rect 138158 79908 138210 79960
rect 137974 79840 138026 79892
rect 137928 79704 137980 79756
rect 138020 79636 138072 79688
rect 138296 79636 138348 79688
rect 138618 79908 138670 79960
rect 138710 79908 138762 79960
rect 138802 79908 138854 79960
rect 139262 79908 139314 79960
rect 139354 79908 139406 79960
rect 139538 79908 139590 79960
rect 139630 79908 139682 79960
rect 139814 79908 139866 79960
rect 139906 79908 139958 79960
rect 140090 79908 140142 79960
rect 140182 79908 140234 79960
rect 140366 79908 140418 79960
rect 140550 79908 140602 79960
rect 138572 79772 138624 79824
rect 138756 79772 138808 79824
rect 139078 79840 139130 79892
rect 139032 79704 139084 79756
rect 139124 79704 139176 79756
rect 139584 79704 139636 79756
rect 138572 79636 138624 79688
rect 138664 79636 138716 79688
rect 139768 79704 139820 79756
rect 136824 79568 136876 79620
rect 137652 79568 137704 79620
rect 138204 79568 138256 79620
rect 140136 79704 140188 79756
rect 140044 79636 140096 79688
rect 140412 79636 140464 79688
rect 141010 79840 141062 79892
rect 141286 79840 141338 79892
rect 141470 79840 141522 79892
rect 141746 79840 141798 79892
rect 140320 79568 140372 79620
rect 140780 79568 140832 79620
rect 140872 79568 140924 79620
rect 136364 79500 136416 79552
rect 136916 79500 136968 79552
rect 138112 79500 138164 79552
rect 140228 79500 140280 79552
rect 133880 79432 133932 79484
rect 141332 79568 141384 79620
rect 141424 79568 141476 79620
rect 141056 79500 141108 79552
rect 141240 79432 141292 79484
rect 141332 79432 141384 79484
rect 139676 79364 139728 79416
rect 140228 79364 140280 79416
rect 140504 79364 140556 79416
rect 142022 79908 142074 79960
rect 142482 79908 142534 79960
rect 142206 79840 142258 79892
rect 142390 79840 142442 79892
rect 142344 79704 142396 79756
rect 142160 79636 142212 79688
rect 142252 79568 142304 79620
rect 142850 79908 142902 79960
rect 143310 79908 143362 79960
rect 142620 79568 142672 79620
rect 143264 79568 143316 79620
rect 143862 79908 143914 79960
rect 144046 79908 144098 79960
rect 144322 79908 144374 79960
rect 144414 79908 144466 79960
rect 144506 79908 144558 79960
rect 144598 79908 144650 79960
rect 144690 79908 144742 79960
rect 144874 79908 144926 79960
rect 144138 79840 144190 79892
rect 144046 79772 144098 79824
rect 143908 79636 143960 79688
rect 143816 79568 143868 79620
rect 144000 79568 144052 79620
rect 144368 79772 144420 79824
rect 144460 79772 144512 79824
rect 144552 79636 144604 79688
rect 144644 79568 144696 79620
rect 142804 79500 142856 79552
rect 143080 79500 143132 79552
rect 144184 79500 144236 79552
rect 144920 79568 144972 79620
rect 141976 79432 142028 79484
rect 146070 79908 146122 79960
rect 146254 79908 146306 79960
rect 146346 79908 146398 79960
rect 146530 79908 146582 79960
rect 146622 79908 146674 79960
rect 145334 79840 145386 79892
rect 145518 79840 145570 79892
rect 145610 79840 145662 79892
rect 145564 79704 145616 79756
rect 146070 79772 146122 79824
rect 145932 79636 145984 79688
rect 146208 79704 146260 79756
rect 146438 79840 146490 79892
rect 146024 79568 146076 79620
rect 146300 79568 146352 79620
rect 146576 79704 146628 79756
rect 145656 79500 145708 79552
rect 146484 79500 146536 79552
rect 146300 79432 146352 79484
rect 186964 81064 187016 81116
rect 187332 81064 187384 81116
rect 195152 81064 195204 81116
rect 214564 81064 214616 81116
rect 214840 81064 214892 81116
rect 186688 80860 186740 80912
rect 215852 80860 215904 80912
rect 234620 80860 234672 80912
rect 187516 80792 187568 80844
rect 252560 80792 252612 80844
rect 146990 79908 147042 79960
rect 146898 79840 146950 79892
rect 147174 79840 147226 79892
rect 147634 79908 147686 79960
rect 148278 79908 148330 79960
rect 148370 79908 148422 79960
rect 147358 79840 147410 79892
rect 147450 79840 147502 79892
rect 148002 79840 148054 79892
rect 147634 79772 147686 79824
rect 148232 79772 148284 79824
rect 148830 79772 148882 79824
rect 147220 79568 147272 79620
rect 147404 79500 147456 79552
rect 147036 79432 147088 79484
rect 148324 79704 148376 79756
rect 147588 79500 147640 79552
rect 147772 79500 147824 79552
rect 148324 79432 148376 79484
rect 148784 79432 148836 79484
rect 147496 79364 147548 79416
rect 148600 79364 148652 79416
rect 149106 79908 149158 79960
rect 149290 79908 149342 79960
rect 149152 79772 149204 79824
rect 149244 79772 149296 79824
rect 149750 79908 149802 79960
rect 150026 79908 150078 79960
rect 150394 79908 150446 79960
rect 150670 79908 150722 79960
rect 151498 79908 151550 79960
rect 151682 79908 151734 79960
rect 151774 79908 151826 79960
rect 151958 79908 152010 79960
rect 152050 79908 152102 79960
rect 152234 79908 152286 79960
rect 149658 79840 149710 79892
rect 149842 79840 149894 79892
rect 150118 79840 150170 79892
rect 149796 79568 149848 79620
rect 149888 79568 149940 79620
rect 149980 79568 150032 79620
rect 150486 79840 150538 79892
rect 150348 79636 150400 79688
rect 149520 79500 149572 79552
rect 150072 79500 150124 79552
rect 149704 79432 149756 79484
rect 151130 79840 151182 79892
rect 150624 79772 150676 79824
rect 151636 79636 151688 79688
rect 152004 79772 152056 79824
rect 151820 79636 151872 79688
rect 152326 79840 152378 79892
rect 152096 79568 152148 79620
rect 152602 79908 152654 79960
rect 152602 79772 152654 79824
rect 152878 79908 152930 79960
rect 153246 79908 153298 79960
rect 153430 79908 153482 79960
rect 153522 79908 153574 79960
rect 153798 79908 153850 79960
rect 153982 79908 154034 79960
rect 152970 79840 153022 79892
rect 152648 79636 152700 79688
rect 152740 79636 152792 79688
rect 152832 79636 152884 79688
rect 153108 79568 153160 79620
rect 153384 79636 153436 79688
rect 153706 79840 153758 79892
rect 153660 79636 153712 79688
rect 153890 79840 153942 79892
rect 153936 79704 153988 79756
rect 153752 79568 153804 79620
rect 153660 79500 153712 79552
rect 154350 79908 154402 79960
rect 154304 79500 154356 79552
rect 151452 79432 151504 79484
rect 151728 79432 151780 79484
rect 153292 79432 153344 79484
rect 154810 79908 154862 79960
rect 155086 79908 155138 79960
rect 155178 79908 155230 79960
rect 154902 79840 154954 79892
rect 154718 79772 154770 79824
rect 154810 79772 154862 79824
rect 154948 79704 155000 79756
rect 154672 79568 154724 79620
rect 154764 79568 154816 79620
rect 155454 79908 155506 79960
rect 155638 79908 155690 79960
rect 155730 79840 155782 79892
rect 155822 79840 155874 79892
rect 155500 79772 155552 79824
rect 155592 79772 155644 79824
rect 155776 79704 155828 79756
rect 156190 79908 156242 79960
rect 156374 79908 156426 79960
rect 156834 79908 156886 79960
rect 156466 79840 156518 79892
rect 156650 79840 156702 79892
rect 156926 79840 156978 79892
rect 156236 79636 156288 79688
rect 156052 79500 156104 79552
rect 156144 79500 156196 79552
rect 156604 79568 156656 79620
rect 156788 79568 156840 79620
rect 157386 79908 157438 79960
rect 157662 79908 157714 79960
rect 157202 79772 157254 79824
rect 157754 79840 157806 79892
rect 157708 79704 157760 79756
rect 157248 79636 157300 79688
rect 157340 79636 157392 79688
rect 157616 79636 157668 79688
rect 157938 79908 157990 79960
rect 158030 79908 158082 79960
rect 158214 79908 158266 79960
rect 158398 79908 158450 79960
rect 158490 79908 158542 79960
rect 158168 79772 158220 79824
rect 157984 79704 158036 79756
rect 158076 79704 158128 79756
rect 158168 79636 158220 79688
rect 158260 79636 158312 79688
rect 157800 79500 157852 79552
rect 158858 79840 158910 79892
rect 158950 79840 159002 79892
rect 158536 79772 158588 79824
rect 158766 79772 158818 79824
rect 155132 79432 155184 79484
rect 155960 79432 156012 79484
rect 157064 79432 157116 79484
rect 158352 79432 158404 79484
rect 158536 79432 158588 79484
rect 158720 79432 158772 79484
rect 159226 79908 159278 79960
rect 159870 79908 159922 79960
rect 159686 79840 159738 79892
rect 159410 79772 159462 79824
rect 158996 79568 159048 79620
rect 159088 79568 159140 79620
rect 159456 79500 159508 79552
rect 160422 79908 160474 79960
rect 160514 79908 160566 79960
rect 160606 79908 160658 79960
rect 160376 79772 160428 79824
rect 160100 79568 160152 79620
rect 160698 79840 160750 79892
rect 160560 79500 160612 79552
rect 159640 79432 159692 79484
rect 159824 79432 159876 79484
rect 160468 79432 160520 79484
rect 161158 79908 161210 79960
rect 161526 79908 161578 79960
rect 161618 79908 161670 79960
rect 161710 79908 161762 79960
rect 161066 79840 161118 79892
rect 161250 79840 161302 79892
rect 161342 79840 161394 79892
rect 161112 79636 161164 79688
rect 161388 79636 161440 79688
rect 161894 79840 161946 79892
rect 161986 79840 162038 79892
rect 161664 79704 161716 79756
rect 161848 79704 161900 79756
rect 161480 79568 161532 79620
rect 161204 79500 161256 79552
rect 161664 79568 161716 79620
rect 161756 79500 161808 79552
rect 160928 79432 160980 79484
rect 162446 79908 162498 79960
rect 162492 79636 162544 79688
rect 182134 80588 182186 80640
rect 162860 79568 162912 79620
rect 163366 79908 163418 79960
rect 164286 79908 164338 79960
rect 163182 79840 163234 79892
rect 163274 79840 163326 79892
rect 163550 79772 163602 79824
rect 164286 79772 164338 79824
rect 163504 79568 163556 79620
rect 164056 79568 164108 79620
rect 162676 79500 162728 79552
rect 163044 79500 163096 79552
rect 163228 79500 163280 79552
rect 164240 79500 164292 79552
rect 164654 79908 164706 79960
rect 178132 80520 178184 80572
rect 187700 80724 187752 80776
rect 270500 80724 270552 80776
rect 186964 80656 187016 80708
rect 189264 80656 189316 80708
rect 288440 80656 288492 80708
rect 186688 80588 186740 80640
rect 184388 80520 184440 80572
rect 187332 80520 187384 80572
rect 187516 80452 187568 80504
rect 164838 79908 164890 79960
rect 165758 79908 165810 79960
rect 165850 79908 165902 79960
rect 165942 79908 165994 79960
rect 165390 79840 165442 79892
rect 165574 79840 165626 79892
rect 164608 79636 164660 79688
rect 165804 79704 165856 79756
rect 165712 79568 165764 79620
rect 165988 79568 166040 79620
rect 166218 79908 166270 79960
rect 166310 79908 166362 79960
rect 166402 79908 166454 79960
rect 166494 79908 166546 79960
rect 166586 79908 166638 79960
rect 167046 79908 167098 79960
rect 166264 79704 166316 79756
rect 166172 79500 166224 79552
rect 165252 79432 165304 79484
rect 165620 79432 165672 79484
rect 166770 79772 166822 79824
rect 166540 79704 166592 79756
rect 166908 79704 166960 79756
rect 167414 79908 167466 79960
rect 168334 79908 168386 79960
rect 168426 79908 168478 79960
rect 168518 79908 168570 79960
rect 168288 79704 168340 79756
rect 167368 79636 167420 79688
rect 167644 79568 167696 79620
rect 166632 79500 166684 79552
rect 166816 79500 166868 79552
rect 166908 79500 166960 79552
rect 167736 79432 167788 79484
rect 168472 79636 168524 79688
rect 168564 79636 168616 79688
rect 169346 79908 169398 79960
rect 169898 79908 169950 79960
rect 169990 79908 170042 79960
rect 170082 79908 170134 79960
rect 170450 79908 170502 79960
rect 169070 79840 169122 79892
rect 168794 79772 168846 79824
rect 168932 79636 168984 79688
rect 168656 79568 168708 79620
rect 169392 79704 169444 79756
rect 169208 79568 169260 79620
rect 170036 79772 170088 79824
rect 170266 79772 170318 79824
rect 169944 79704 169996 79756
rect 170496 79704 170548 79756
rect 170220 79636 170272 79688
rect 170910 79908 170962 79960
rect 171002 79908 171054 79960
rect 170818 79840 170870 79892
rect 170956 79636 171008 79688
rect 178592 80384 178644 80436
rect 182180 80384 182232 80436
rect 191104 80384 191156 80436
rect 177764 80248 177816 80300
rect 179512 80180 179564 80232
rect 171370 79908 171422 79960
rect 171646 79908 171698 79960
rect 171738 79908 171790 79960
rect 171922 79908 171974 79960
rect 172382 79908 172434 79960
rect 171324 79772 171376 79824
rect 170772 79568 170824 79620
rect 171140 79568 171192 79620
rect 170588 79500 170640 79552
rect 172014 79840 172066 79892
rect 172566 79908 172618 79960
rect 172658 79908 172710 79960
rect 172750 79908 172802 79960
rect 172520 79772 172572 79824
rect 172428 79704 172480 79756
rect 171784 79568 171836 79620
rect 171968 79568 172020 79620
rect 172520 79568 172572 79620
rect 177764 80112 177816 80164
rect 173026 79908 173078 79960
rect 173302 79908 173354 79960
rect 178040 80044 178092 80096
rect 178224 79976 178276 80028
rect 201224 80044 201276 80096
rect 525800 80044 525852 80096
rect 173578 79908 173630 79960
rect 173946 79908 173998 79960
rect 173394 79772 173446 79824
rect 173072 79636 173124 79688
rect 173164 79568 173216 79620
rect 173440 79568 173492 79620
rect 172152 79500 172204 79552
rect 171876 79432 171928 79484
rect 172612 79432 172664 79484
rect 173762 79840 173814 79892
rect 174222 79840 174274 79892
rect 174498 79840 174550 79892
rect 173716 79636 173768 79688
rect 173900 79500 173952 79552
rect 174544 79568 174596 79620
rect 174774 79908 174826 79960
rect 175050 79908 175102 79960
rect 175142 79908 175194 79960
rect 175234 79908 175286 79960
rect 175418 79908 175470 79960
rect 175510 79908 175562 79960
rect 175970 79908 176022 79960
rect 176982 79908 177034 79960
rect 174958 79840 175010 79892
rect 174820 79704 174872 79756
rect 175004 79704 175056 79756
rect 175188 79704 175240 79756
rect 175280 79568 175332 79620
rect 175786 79840 175838 79892
rect 176246 79840 176298 79892
rect 176338 79840 176390 79892
rect 176522 79840 176574 79892
rect 176108 79636 176160 79688
rect 176200 79636 176252 79688
rect 176384 79636 176436 79688
rect 176568 79636 176620 79688
rect 176844 79636 176896 79688
rect 177074 79840 177126 79892
rect 177764 79840 177816 79892
rect 175556 79500 175608 79552
rect 173992 79432 174044 79484
rect 175464 79432 175516 79484
rect 175924 79432 175976 79484
rect 178132 79568 178184 79620
rect 191196 79568 191248 79620
rect 178316 79500 178368 79552
rect 192576 79500 192628 79552
rect 217140 79500 217192 79552
rect 217416 79500 217468 79552
rect 178960 79432 179012 79484
rect 187148 79432 187200 79484
rect 194508 79432 194560 79484
rect 340880 79432 340932 79484
rect 120540 79296 120592 79348
rect 147772 79296 147824 79348
rect 119160 79228 119212 79280
rect 146300 79228 146352 79280
rect 146392 79228 146444 79280
rect 162124 79364 162176 79416
rect 149244 79296 149296 79348
rect 153936 79228 153988 79280
rect 154120 79228 154172 79280
rect 116308 79160 116360 79212
rect 152096 79160 152148 79212
rect 158352 79296 158404 79348
rect 162860 79296 162912 79348
rect 174360 79364 174412 79416
rect 179144 79364 179196 79416
rect 207756 79364 207808 79416
rect 376760 79364 376812 79416
rect 165252 79296 165304 79348
rect 211436 79296 211488 79348
rect 214380 79296 214432 79348
rect 448520 79296 448572 79348
rect 170864 79228 170916 79280
rect 193128 79228 193180 79280
rect 115572 79092 115624 79144
rect 142252 79092 142304 79144
rect 142804 79092 142856 79144
rect 143540 79092 143592 79144
rect 144920 79092 144972 79144
rect 146024 79092 146076 79144
rect 118056 79024 118108 79076
rect 148692 79024 148744 79076
rect 112720 78956 112772 79008
rect 144736 78956 144788 79008
rect 171232 79160 171284 79212
rect 157800 79092 157852 79144
rect 158076 79092 158128 79144
rect 162124 79092 162176 79144
rect 166172 79092 166224 79144
rect 179052 79092 179104 79144
rect 180984 79160 181036 79212
rect 198188 79160 198240 79212
rect 206192 79160 206244 79212
rect 206560 79160 206612 79212
rect 204628 79092 204680 79144
rect 156052 79024 156104 79076
rect 156696 79024 156748 79076
rect 158996 79024 159048 79076
rect 193864 79024 193916 79076
rect 194508 79024 194560 79076
rect 162676 78956 162728 79008
rect 167736 78956 167788 79008
rect 201684 78956 201736 79008
rect 115204 78888 115256 78940
rect 147680 78888 147732 78940
rect 169760 78888 169812 78940
rect 204904 78888 204956 78940
rect 112444 78820 112496 78872
rect 146116 78820 146168 78872
rect 167276 78820 167328 78872
rect 214380 78820 214432 78872
rect 130292 78752 130344 78804
rect 100300 78548 100352 78600
rect 113916 78684 113968 78736
rect 138204 78684 138256 78736
rect 138572 78684 138624 78736
rect 143632 78684 143684 78736
rect 144276 78684 144328 78736
rect 144552 78684 144604 78736
rect 144920 78684 144972 78736
rect 157156 78684 157208 78736
rect 160744 78684 160796 78736
rect 105268 78480 105320 78532
rect 138664 78616 138716 78668
rect 139952 78616 140004 78668
rect 140136 78616 140188 78668
rect 140504 78616 140556 78668
rect 145012 78616 145064 78668
rect 147956 78616 148008 78668
rect 148324 78616 148376 78668
rect 157432 78616 157484 78668
rect 157892 78616 157944 78668
rect 158168 78616 158220 78668
rect 158352 78616 158404 78668
rect 159272 78616 159324 78668
rect 159456 78616 159508 78668
rect 113916 78548 113968 78600
rect 122196 78480 122248 78532
rect 105544 78412 105596 78464
rect 105728 78412 105780 78464
rect 136916 78412 136968 78464
rect 60740 78276 60792 78328
rect 107200 78344 107252 78396
rect 137192 78344 137244 78396
rect 75920 78208 75972 78260
rect 105728 78208 105780 78260
rect 57980 78072 58032 78124
rect 107292 78072 107344 78124
rect 136272 78276 136324 78328
rect 161480 78548 161532 78600
rect 161664 78548 161716 78600
rect 185584 78752 185636 78804
rect 209228 78752 209280 78804
rect 480260 78752 480312 78804
rect 171048 78684 171100 78736
rect 174728 78684 174780 78736
rect 211804 78684 211856 78736
rect 483020 78684 483072 78736
rect 169944 78616 169996 78668
rect 171508 78548 171560 78600
rect 172244 78548 172296 78600
rect 179052 78616 179104 78668
rect 179236 78616 179288 78668
rect 200948 78616 201000 78668
rect 211804 78548 211856 78600
rect 169944 78480 169996 78532
rect 153936 78412 153988 78464
rect 161664 78412 161716 78464
rect 162492 78412 162544 78464
rect 165160 78412 165212 78464
rect 199108 78480 199160 78532
rect 199568 78480 199620 78532
rect 139584 78344 139636 78396
rect 140412 78344 140464 78396
rect 147956 78344 148008 78396
rect 149152 78344 149204 78396
rect 163136 78344 163188 78396
rect 197636 78412 197688 78464
rect 143540 78276 143592 78328
rect 53840 78004 53892 78056
rect 106924 78004 106976 78056
rect 136548 78208 136600 78260
rect 145840 78208 145892 78260
rect 160744 78208 160796 78260
rect 162492 78208 162544 78260
rect 164240 78208 164292 78260
rect 198740 78344 198792 78396
rect 171140 78276 171192 78328
rect 203524 78276 203576 78328
rect 172428 78208 172480 78260
rect 180064 78208 180116 78260
rect 46940 77936 46992 77988
rect 107016 77936 107068 77988
rect 135260 78140 135312 78192
rect 136732 78140 136784 78192
rect 137284 78140 137336 78192
rect 140136 78140 140188 78192
rect 140780 78140 140832 78192
rect 142252 78140 142304 78192
rect 145288 78140 145340 78192
rect 152924 78140 152976 78192
rect 156236 78140 156288 78192
rect 164148 78140 164200 78192
rect 178776 78140 178828 78192
rect 179144 78140 179196 78192
rect 179328 78140 179380 78192
rect 213092 78140 213144 78192
rect 120724 78072 120776 78124
rect 145656 78072 145708 78124
rect 164240 78072 164292 78124
rect 164792 78072 164844 78124
rect 169392 78072 169444 78124
rect 169576 78072 169628 78124
rect 171140 78072 171192 78124
rect 171324 78072 171376 78124
rect 187700 78072 187752 78124
rect 197636 78072 197688 78124
rect 198464 78072 198516 78124
rect 393320 78072 393372 78124
rect 108304 78004 108356 78056
rect 129832 78004 129884 78056
rect 130660 78004 130712 78056
rect 130752 78004 130804 78056
rect 142068 78004 142120 78056
rect 152924 78004 152976 78056
rect 153200 78004 153252 78056
rect 158444 78004 158496 78056
rect 162216 78004 162268 78056
rect 164056 78004 164108 78056
rect 178684 78004 178736 78056
rect 178960 78004 179012 78056
rect 198740 78004 198792 78056
rect 199476 78004 199528 78056
rect 415492 78004 415544 78056
rect 108396 77936 108448 77988
rect 131212 77936 131264 77988
rect 142528 77936 142580 77988
rect 156512 77936 156564 77988
rect 156880 77936 156932 77988
rect 166908 77936 166960 77988
rect 170496 77936 170548 77988
rect 175556 77936 175608 77988
rect 176108 77936 176160 77988
rect 177948 77936 178000 77988
rect 181996 77936 182048 77988
rect 199108 77936 199160 77988
rect 422300 77936 422352 77988
rect 109500 77868 109552 77920
rect 129740 77868 129792 77920
rect 130660 77868 130712 77920
rect 137376 77868 137428 77920
rect 138756 77868 138808 77920
rect 139308 77868 139360 77920
rect 143816 77868 143868 77920
rect 144460 77868 144512 77920
rect 168288 77868 168340 77920
rect 180616 77868 180668 77920
rect 201776 77868 201828 77920
rect 108120 77800 108172 77852
rect 128544 77800 128596 77852
rect 129924 77800 129976 77852
rect 133880 77800 133932 77852
rect 134524 77800 134576 77852
rect 142252 77800 142304 77852
rect 170496 77800 170548 77852
rect 179144 77800 179196 77852
rect 179328 77800 179380 77852
rect 179972 77800 180024 77852
rect 191288 77800 191340 77852
rect 99840 77732 99892 77784
rect 130936 77732 130988 77784
rect 139492 77732 139544 77784
rect 162400 77732 162452 77784
rect 162768 77732 162820 77784
rect 167184 77732 167236 77784
rect 179052 77732 179104 77784
rect 130660 77664 130712 77716
rect 131028 77664 131080 77716
rect 144092 77664 144144 77716
rect 148416 77664 148468 77716
rect 207848 77664 207900 77716
rect 132868 77596 132920 77648
rect 133880 77596 133932 77648
rect 134340 77596 134392 77648
rect 140412 77596 140464 77648
rect 140688 77596 140740 77648
rect 150900 77596 150952 77648
rect 169944 77596 169996 77648
rect 175740 77596 175792 77648
rect 176200 77596 176252 77648
rect 176660 77596 176712 77648
rect 176844 77596 176896 77648
rect 177764 77596 177816 77648
rect 211712 77596 211764 77648
rect 145012 77528 145064 77580
rect 145564 77528 145616 77580
rect 157524 77528 157576 77580
rect 170864 77528 170916 77580
rect 174360 77528 174412 77580
rect 178868 77528 178920 77580
rect 146300 77460 146352 77512
rect 146852 77460 146904 77512
rect 148692 77460 148744 77512
rect 148968 77460 149020 77512
rect 161848 77460 161900 77512
rect 162400 77460 162452 77512
rect 167368 77460 167420 77512
rect 178500 77460 178552 77512
rect 133052 77392 133104 77444
rect 146024 77392 146076 77444
rect 146944 77392 146996 77444
rect 169944 77392 169996 77444
rect 170680 77392 170732 77444
rect 132592 77324 132644 77376
rect 132776 77324 132828 77376
rect 133236 77324 133288 77376
rect 135628 77324 135680 77376
rect 136272 77324 136324 77376
rect 175832 77324 175884 77376
rect 176568 77324 176620 77376
rect 109040 77256 109092 77308
rect 109500 77256 109552 77308
rect 132500 77256 132552 77308
rect 133420 77256 133472 77308
rect 135812 77256 135864 77308
rect 136180 77256 136232 77308
rect 138296 77256 138348 77308
rect 138480 77256 138532 77308
rect 154948 77256 155000 77308
rect 164884 77256 164936 77308
rect 174176 77256 174228 77308
rect 177580 77256 177632 77308
rect 187700 77256 187752 77308
rect 500960 77256 501012 77308
rect 111248 77188 111300 77240
rect 145104 77188 145156 77240
rect 146024 77188 146076 77240
rect 155500 77188 155552 77240
rect 217140 77188 217192 77240
rect 124864 77120 124916 77172
rect 125600 77120 125652 77172
rect 141884 77120 141936 77172
rect 145932 77120 145984 77172
rect 148324 77120 148376 77172
rect 102140 77052 102192 77104
rect 102876 77052 102928 77104
rect 137468 77052 137520 77104
rect 114468 76984 114520 77036
rect 147128 76984 147180 77036
rect 114284 76916 114336 76968
rect 146760 76916 146812 76968
rect 115296 76848 115348 76900
rect 149704 76848 149756 76900
rect 152188 76848 152240 76900
rect 213184 77120 213236 77172
rect 164884 77052 164936 77104
rect 170036 76984 170088 77036
rect 170772 76984 170824 77036
rect 171232 76984 171284 77036
rect 171416 76984 171468 77036
rect 174176 76984 174228 77036
rect 174912 76984 174964 77036
rect 175464 76984 175516 77036
rect 210516 76984 210568 77036
rect 165344 76916 165396 76968
rect 199384 76916 199436 76968
rect 160192 76848 160244 76900
rect 160744 76848 160796 76900
rect 161572 76848 161624 76900
rect 164148 76848 164200 76900
rect 165804 76848 165856 76900
rect 166172 76848 166224 76900
rect 169852 76848 169904 76900
rect 170312 76848 170364 76900
rect 172704 76848 172756 76900
rect 173532 76848 173584 76900
rect 175464 76848 175516 76900
rect 176384 76848 176436 76900
rect 177856 76848 177908 76900
rect 210424 76848 210476 76900
rect 112996 76780 113048 76832
rect 144368 76780 144420 76832
rect 153292 76780 153344 76832
rect 154028 76780 154080 76832
rect 114376 76712 114428 76764
rect 145748 76712 145800 76764
rect 152556 76712 152608 76764
rect 99380 76644 99432 76696
rect 110880 76644 110932 76696
rect 140044 76644 140096 76696
rect 140964 76644 141016 76696
rect 141240 76644 141292 76696
rect 150532 76644 150584 76696
rect 151636 76644 151688 76696
rect 151912 76644 151964 76696
rect 152464 76644 152516 76696
rect 159824 76644 159876 76696
rect 189264 76780 189316 76832
rect 193128 76780 193180 76832
rect 214564 76780 214616 76832
rect 247684 76848 247736 76900
rect 162860 76712 162912 76764
rect 163688 76712 163740 76764
rect 164332 76712 164384 76764
rect 164792 76712 164844 76764
rect 167368 76712 167420 76764
rect 167552 76712 167604 76764
rect 174268 76712 174320 76764
rect 175188 76712 175240 76764
rect 176016 76712 176068 76764
rect 176200 76712 176252 76764
rect 177212 76712 177264 76764
rect 206652 76712 206704 76764
rect 160192 76644 160244 76696
rect 160376 76644 160428 76696
rect 160836 76644 160888 76696
rect 161296 76644 161348 76696
rect 161572 76644 161624 76696
rect 161940 76644 161992 76696
rect 163228 76644 163280 76696
rect 163412 76644 163464 76696
rect 164700 76644 164752 76696
rect 165068 76644 165120 76696
rect 165896 76644 165948 76696
rect 166080 76644 166132 76696
rect 167184 76644 167236 76696
rect 167460 76644 167512 76696
rect 168564 76644 168616 76696
rect 169116 76644 169168 76696
rect 171140 76644 171192 76696
rect 171968 76644 172020 76696
rect 172428 76644 172480 76696
rect 198096 76644 198148 76696
rect 217324 76780 217376 76832
rect 289820 76780 289872 76832
rect 217140 76712 217192 76764
rect 296720 76712 296772 76764
rect 324320 76644 324372 76696
rect 66260 76576 66312 76628
rect 102140 76576 102192 76628
rect 113824 76576 113876 76628
rect 141148 76576 141200 76628
rect 147312 76576 147364 76628
rect 181444 76576 181496 76628
rect 189264 76576 189316 76628
rect 189724 76576 189776 76628
rect 353300 76576 353352 76628
rect 59360 76508 59412 76560
rect 102968 76508 103020 76560
rect 114560 76508 114612 76560
rect 132776 76508 132828 76560
rect 132960 76508 133012 76560
rect 133788 76508 133840 76560
rect 135628 76508 135680 76560
rect 136088 76508 136140 76560
rect 136640 76508 136692 76560
rect 137468 76508 137520 76560
rect 146760 76508 146812 76560
rect 184940 76508 184992 76560
rect 111708 76440 111760 76492
rect 137652 76440 137704 76492
rect 154948 76440 155000 76492
rect 155408 76440 155460 76492
rect 155960 76440 156012 76492
rect 157064 76440 157116 76492
rect 158720 76440 158772 76492
rect 159088 76440 159140 76492
rect 163228 76440 163280 76492
rect 163964 76440 164016 76492
rect 164332 76440 164384 76492
rect 164516 76440 164568 76492
rect 178592 76440 178644 76492
rect 187700 76440 187752 76492
rect 110972 76372 111024 76424
rect 126980 76372 127032 76424
rect 134340 76372 134392 76424
rect 135168 76372 135220 76424
rect 135444 76372 135496 76424
rect 136088 76372 136140 76424
rect 150440 76372 150492 76424
rect 151268 76372 151320 76424
rect 163780 76372 163832 76424
rect 166356 76372 166408 76424
rect 136824 76304 136876 76356
rect 161020 76304 161072 76356
rect 187424 76304 187476 76356
rect 367100 76508 367152 76560
rect 164516 76236 164568 76288
rect 165436 76236 165488 76288
rect 166080 76236 166132 76288
rect 166816 76236 166868 76288
rect 132776 76168 132828 76220
rect 140872 76168 140924 76220
rect 171784 76100 171836 76152
rect 172428 76100 172480 76152
rect 132776 76032 132828 76084
rect 133604 76032 133656 76084
rect 144368 75964 144420 76016
rect 146300 75964 146352 76016
rect 173348 75896 173400 75948
rect 173624 75896 173676 75948
rect 177212 75896 177264 75948
rect 177672 75896 177724 75948
rect 210516 75896 210568 75948
rect 553400 75896 553452 75948
rect 103060 75828 103112 75880
rect 103888 75760 103940 75812
rect 104072 75760 104124 75812
rect 138940 75760 138992 75812
rect 140044 75828 140096 75880
rect 140228 75828 140280 75880
rect 166632 75828 166684 75880
rect 200764 75828 200816 75880
rect 144828 75760 144880 75812
rect 111892 75692 111944 75744
rect 100760 75624 100812 75676
rect 101220 75624 101272 75676
rect 135076 75624 135128 75676
rect 135352 75624 135404 75676
rect 135904 75624 135956 75676
rect 104440 75556 104492 75608
rect 137560 75556 137612 75608
rect 138204 75692 138256 75744
rect 139216 75692 139268 75744
rect 139768 75692 139820 75744
rect 140228 75692 140280 75744
rect 142528 75624 142580 75676
rect 142804 75624 142856 75676
rect 93860 75488 93912 75540
rect 105268 75488 105320 75540
rect 116584 75488 116636 75540
rect 104256 75420 104308 75472
rect 131028 75420 131080 75472
rect 131120 75420 131172 75472
rect 132592 75420 132644 75472
rect 85580 75352 85632 75404
rect 103888 75352 103940 75404
rect 117228 75352 117280 75404
rect 146484 75556 146536 75608
rect 158628 75556 158680 75608
rect 175096 75760 175148 75812
rect 204904 75760 204956 75812
rect 172980 75692 173032 75744
rect 207572 75692 207624 75744
rect 208308 75692 208360 75744
rect 170588 75624 170640 75676
rect 171048 75624 171100 75676
rect 204720 75624 204772 75676
rect 144828 75488 144880 75540
rect 147036 75488 147088 75540
rect 154580 75488 154632 75540
rect 155500 75488 155552 75540
rect 156144 75488 156196 75540
rect 156788 75488 156840 75540
rect 180800 75556 180852 75608
rect 179972 75488 180024 75540
rect 180708 75488 180760 75540
rect 216680 75488 216732 75540
rect 146668 75420 146720 75472
rect 176752 75420 176804 75472
rect 176936 75420 176988 75472
rect 177120 75420 177172 75472
rect 99012 75284 99064 75336
rect 131120 75284 131172 75336
rect 137008 75284 137060 75336
rect 137192 75284 137244 75336
rect 145472 75284 145524 75336
rect 71044 75216 71096 75268
rect 104440 75216 104492 75268
rect 118608 75216 118660 75268
rect 138020 75216 138072 75268
rect 138112 75216 138164 75268
rect 138480 75216 138532 75268
rect 141240 75216 141292 75268
rect 141608 75216 141660 75268
rect 142896 75216 142948 75268
rect 143356 75216 143408 75268
rect 143908 75216 143960 75268
rect 144092 75216 144144 75268
rect 145196 75216 145248 75268
rect 145748 75216 145800 75268
rect 35900 75148 35952 75200
rect 100760 75148 100812 75200
rect 112444 75148 112496 75200
rect 97908 75080 97960 75132
rect 114560 75080 114612 75132
rect 121092 75080 121144 75132
rect 141148 75148 141200 75200
rect 141976 75148 142028 75200
rect 142712 75148 142764 75200
rect 143172 75148 143224 75200
rect 151084 75352 151136 75404
rect 216680 75352 216732 75404
rect 149704 75284 149756 75336
rect 187700 75284 187752 75336
rect 191748 75284 191800 75336
rect 305000 75284 305052 75336
rect 147496 75216 147548 75268
rect 193864 75216 193916 75268
rect 204904 75216 204956 75268
rect 442264 75216 442316 75268
rect 148048 75148 148100 75200
rect 108580 75012 108632 75064
rect 130568 75012 130620 75064
rect 130936 75012 130988 75064
rect 140964 75080 141016 75132
rect 142436 75080 142488 75132
rect 143264 75080 143316 75132
rect 149336 75080 149388 75132
rect 149980 75080 150032 75132
rect 152004 75148 152056 75200
rect 153016 75148 153068 75200
rect 156052 75148 156104 75200
rect 156972 75148 157024 75200
rect 201684 75148 201736 75200
rect 208308 75148 208360 75200
rect 521660 75148 521712 75200
rect 158720 75080 158772 75132
rect 160008 75080 160060 75132
rect 165712 75080 165764 75132
rect 189632 75080 189684 75132
rect 146576 75012 146628 75064
rect 151636 75012 151688 75064
rect 151820 75012 151872 75064
rect 154672 75012 154724 75064
rect 155592 75012 155644 75064
rect 158904 75012 158956 75064
rect 159916 75012 159968 75064
rect 131304 74944 131356 74996
rect 137008 74944 137060 74996
rect 137744 74944 137796 74996
rect 138020 74944 138072 74996
rect 145196 74944 145248 74996
rect 139308 74876 139360 74928
rect 143724 74876 143776 74928
rect 144736 74876 144788 74928
rect 131028 74808 131080 74860
rect 135352 74808 135404 74860
rect 156328 74808 156380 74860
rect 191380 75012 191432 75064
rect 191748 75012 191800 75064
rect 173164 74944 173216 74996
rect 173532 74944 173584 74996
rect 176752 74944 176804 74996
rect 185032 74944 185084 74996
rect 181996 74876 182048 74928
rect 210792 74944 210844 74996
rect 173072 74808 173124 74860
rect 177948 74808 178000 74860
rect 211344 74876 211396 74928
rect 161756 74740 161808 74792
rect 162676 74740 162728 74792
rect 130660 74672 130712 74724
rect 131028 74672 131080 74724
rect 167092 74536 167144 74588
rect 167736 74536 167788 74588
rect 128544 74468 128596 74520
rect 139584 74468 139636 74520
rect 142252 74468 142304 74520
rect 143080 74468 143132 74520
rect 152648 74468 152700 74520
rect 218336 74468 218388 74520
rect 119436 74400 119488 74452
rect 153844 74400 153896 74452
rect 159640 74400 159692 74452
rect 218152 74400 218204 74452
rect 106740 74332 106792 74384
rect 140596 74332 140648 74384
rect 153752 74332 153804 74384
rect 154488 74332 154540 74384
rect 156236 74332 156288 74384
rect 188528 74332 188580 74384
rect 115388 74264 115440 74316
rect 147864 74264 147916 74316
rect 148692 74264 148744 74316
rect 165068 74264 165120 74316
rect 165712 74264 165764 74316
rect 168288 74264 168340 74316
rect 202328 74264 202380 74316
rect 109960 74196 110012 74248
rect 142528 74196 142580 74248
rect 153844 74196 153896 74248
rect 154396 74196 154448 74248
rect 155868 74196 155920 74248
rect 156972 74196 157024 74248
rect 108488 74128 108540 74180
rect 140412 74128 140464 74180
rect 149152 74128 149204 74180
rect 156788 74128 156840 74180
rect 159456 74196 159508 74248
rect 194048 74196 194100 74248
rect 189080 74128 189132 74180
rect 218244 74128 218296 74180
rect 218612 74128 218664 74180
rect 121184 74060 121236 74112
rect 152924 74060 152976 74112
rect 163136 74060 163188 74112
rect 163872 74060 163924 74112
rect 165712 74060 165764 74112
rect 166540 74060 166592 74112
rect 167276 74060 167328 74112
rect 168196 74060 168248 74112
rect 119068 73992 119120 74044
rect 151636 73992 151688 74044
rect 159732 73992 159784 74044
rect 159916 73992 159968 74044
rect 164148 73992 164200 74044
rect 196992 74060 197044 74112
rect 175280 73992 175332 74044
rect 206376 73992 206428 74044
rect 218336 73992 218388 74044
rect 255320 73992 255372 74044
rect 111340 73924 111392 73976
rect 142252 73924 142304 73976
rect 158536 73924 158588 73976
rect 159824 73924 159876 73976
rect 163504 73924 163556 73976
rect 168196 73924 168248 73976
rect 170220 73924 170272 73976
rect 180524 73924 180576 73976
rect 188528 73924 188580 73976
rect 261484 73924 261536 73976
rect 89720 73856 89772 73908
rect 8944 73788 8996 73840
rect 119344 73856 119396 73908
rect 149244 73856 149296 73908
rect 149980 73856 150032 73908
rect 173716 73856 173768 73908
rect 203616 73856 203668 73908
rect 218152 73856 218204 73908
rect 347780 73856 347832 73908
rect 107200 73788 107252 73840
rect 136364 73788 136416 73840
rect 159364 73788 159416 73840
rect 160008 73788 160060 73840
rect 162216 73788 162268 73840
rect 192944 73788 192996 73840
rect 322940 73788 322992 73840
rect 104348 73720 104400 73772
rect 139124 73720 139176 73772
rect 157984 73720 158036 73772
rect 158536 73720 158588 73772
rect 180524 73720 180576 73772
rect 208860 73720 208912 73772
rect 105912 73652 105964 73704
rect 132408 73652 132460 73704
rect 179052 73652 179104 73704
rect 201500 73652 201552 73704
rect 122012 73584 122064 73636
rect 128452 73584 128504 73636
rect 129648 73584 129700 73636
rect 152280 73584 152332 73636
rect 153016 73584 153068 73636
rect 162124 73584 162176 73636
rect 167920 73584 167972 73636
rect 106280 73176 106332 73228
rect 106740 73176 106792 73228
rect 107660 73176 107712 73228
rect 108488 73176 108540 73228
rect 121368 73108 121420 73160
rect 149612 73108 149664 73160
rect 149888 73108 149940 73160
rect 161112 73108 161164 73160
rect 195244 73108 195296 73160
rect 327724 73108 327776 73160
rect 579620 73108 579672 73160
rect 121276 73040 121328 73092
rect 129924 73040 129976 73092
rect 130752 73040 130804 73092
rect 131396 73040 131448 73092
rect 132500 73040 132552 73092
rect 142344 73040 142396 73092
rect 143448 73040 143500 73092
rect 159088 73040 159140 73092
rect 194140 73040 194192 73092
rect 115664 72972 115716 73024
rect 147864 72972 147916 73024
rect 148508 72972 148560 73024
rect 156696 72972 156748 73024
rect 157156 72972 157208 73024
rect 210332 72972 210384 73024
rect 52460 72564 52512 72616
rect 102600 72904 102652 72956
rect 136456 72904 136508 72956
rect 157248 72904 157300 72956
rect 191012 72904 191064 72956
rect 107108 72836 107160 72888
rect 140320 72836 140372 72888
rect 157708 72836 157760 72888
rect 192484 72836 192536 72888
rect 110236 72768 110288 72820
rect 142160 72768 142212 72820
rect 158260 72768 158312 72820
rect 191840 72768 191892 72820
rect 117136 72700 117188 72752
rect 148416 72700 148468 72752
rect 150900 72700 150952 72752
rect 154488 72700 154540 72752
rect 187240 72700 187292 72752
rect 218152 72836 218204 72888
rect 218612 72836 218664 72888
rect 229744 72836 229796 72888
rect 216956 72768 217008 72820
rect 342904 72768 342956 72820
rect 318800 72700 318852 72752
rect 96620 72632 96672 72684
rect 107108 72632 107160 72684
rect 111524 72632 111576 72684
rect 142344 72632 142396 72684
rect 155868 72632 155920 72684
rect 188344 72632 188396 72684
rect 192484 72632 192536 72684
rect 323584 72632 323636 72684
rect 118516 72564 118568 72616
rect 148140 72564 148192 72616
rect 148600 72564 148652 72616
rect 158352 72564 158404 72616
rect 188160 72564 188212 72616
rect 332600 72564 332652 72616
rect 9680 72496 9732 72548
rect 98828 72496 98880 72548
rect 99104 72496 99156 72548
rect 131396 72496 131448 72548
rect 156420 72496 156472 72548
rect 157156 72496 157208 72548
rect 190276 72496 190328 72548
rect 194140 72496 194192 72548
rect 340972 72496 341024 72548
rect 4160 72428 4212 72480
rect 99196 72428 99248 72480
rect 109684 72428 109736 72480
rect 138204 72428 138256 72480
rect 146576 72428 146628 72480
rect 182180 72428 182232 72480
rect 195244 72428 195296 72480
rect 368480 72428 368532 72480
rect 109776 72360 109828 72412
rect 121460 72360 121512 72412
rect 141516 72360 141568 72412
rect 161388 72360 161440 72412
rect 194232 72360 194284 72412
rect 98828 72292 98880 72344
rect 133144 72292 133196 72344
rect 159180 72292 159232 72344
rect 216956 72292 217008 72344
rect 99196 72224 99248 72276
rect 132592 72224 132644 72276
rect 155684 72224 155736 72276
rect 218152 72224 218204 72276
rect 3516 71680 3568 71732
rect 13084 71680 13136 71732
rect 121920 71680 121972 71732
rect 149796 71680 149848 71732
rect 161112 71680 161164 71732
rect 192300 71680 192352 71732
rect 105820 71612 105872 71664
rect 140044 71612 140096 71664
rect 157524 71612 157576 71664
rect 158260 71612 158312 71664
rect 159916 71612 159968 71664
rect 193772 71612 193824 71664
rect 104532 71544 104584 71596
rect 137928 71544 137980 71596
rect 192392 71544 192444 71596
rect 118148 71476 118200 71528
rect 147956 71476 148008 71528
rect 150164 71476 150216 71528
rect 157340 71476 157392 71528
rect 158444 71476 158496 71528
rect 160744 71476 160796 71528
rect 195060 71476 195112 71528
rect 116860 71408 116912 71460
rect 148232 71408 148284 71460
rect 148508 71408 148560 71460
rect 159824 71408 159876 71460
rect 193680 71408 193732 71460
rect 134984 71340 135036 71392
rect 157340 71340 157392 71392
rect 157800 71340 157852 71392
rect 158444 71340 158496 71392
rect 161112 71340 161164 71392
rect 162768 71340 162820 71392
rect 196532 71340 196584 71392
rect 71780 71136 71832 71188
rect 104532 71136 104584 71188
rect 35164 71068 35216 71120
rect 103244 71068 103296 71120
rect 119620 71272 119672 71324
rect 150072 71272 150124 71324
rect 166264 71272 166316 71324
rect 166908 71272 166960 71324
rect 200672 71272 200724 71324
rect 112076 71204 112128 71256
rect 142804 71204 142856 71256
rect 160928 71204 160980 71256
rect 195520 71204 195572 71256
rect 122104 71136 122156 71188
rect 151452 71136 151504 71188
rect 153568 71136 153620 71188
rect 187056 71136 187108 71188
rect 27620 71000 27672 71052
rect 99932 71000 99984 71052
rect 107384 71000 107436 71052
rect 133420 71068 133472 71120
rect 147128 71068 147180 71120
rect 184204 71068 184256 71120
rect 111708 71000 111760 71052
rect 128360 71000 128412 71052
rect 129556 71000 129608 71052
rect 150900 71000 150952 71052
rect 200120 71000 200172 71052
rect 134432 70932 134484 70984
rect 160008 70932 160060 70984
rect 192852 70932 192904 70984
rect 157064 70864 157116 70916
rect 188620 70864 188672 70916
rect 158536 70796 158588 70848
rect 188068 70796 188120 70848
rect 169208 70728 169260 70780
rect 169392 70728 169444 70780
rect 149796 70592 149848 70644
rect 150256 70592 150308 70644
rect 103520 70388 103572 70440
rect 105820 70388 105872 70440
rect 113180 70388 113232 70440
rect 115112 70388 115164 70440
rect 100760 70320 100812 70372
rect 101312 70320 101364 70372
rect 135996 70320 136048 70372
rect 168012 70320 168064 70372
rect 214288 70320 214340 70372
rect 118884 70252 118936 70304
rect 152096 70252 152148 70304
rect 152648 70252 152700 70304
rect 164056 70252 164108 70304
rect 204996 70252 205048 70304
rect 104164 70184 104216 70236
rect 137192 70184 137244 70236
rect 161848 70184 161900 70236
rect 196624 70184 196676 70236
rect 85672 69776 85724 69828
rect 106004 70116 106056 70168
rect 139032 70116 139084 70168
rect 162308 70116 162360 70168
rect 196716 70116 196768 70168
rect 108396 70048 108448 70100
rect 108672 70048 108724 70100
rect 139952 70048 140004 70100
rect 160468 70048 160520 70100
rect 161204 70048 161256 70100
rect 194968 70048 195020 70100
rect 120816 69980 120868 70032
rect 150992 69980 151044 70032
rect 163964 69980 164016 70032
rect 197912 69980 197964 70032
rect 111984 69912 112036 69964
rect 142436 69912 142488 69964
rect 163320 69912 163372 69964
rect 164056 69912 164108 69964
rect 165160 69912 165212 69964
rect 199292 69912 199344 69964
rect 113548 69844 113600 69896
rect 142988 69844 143040 69896
rect 151360 69844 151412 69896
rect 242164 69844 242216 69896
rect 115112 69776 115164 69828
rect 141332 69776 141384 69828
rect 150992 69776 151044 69828
rect 151544 69776 151596 69828
rect 160376 69776 160428 69828
rect 194692 69776 194744 69828
rect 362960 69776 363012 69828
rect 60832 69708 60884 69760
rect 104164 69708 104216 69760
rect 117320 69708 117372 69760
rect 117780 69708 117832 69760
rect 141056 69708 141108 69760
rect 163412 69708 163464 69760
rect 163964 69708 164016 69760
rect 164792 69708 164844 69760
rect 165160 69708 165212 69760
rect 166172 69708 166224 69760
rect 45560 69640 45612 69692
rect 100760 69640 100812 69692
rect 102876 69640 102928 69692
rect 108396 69640 108448 69692
rect 148600 69640 148652 69692
rect 189724 69640 189776 69692
rect 214288 69708 214340 69760
rect 397460 69708 397512 69760
rect 201132 69640 201184 69692
rect 430580 69640 430632 69692
rect 161940 69572 161992 69624
rect 162676 69572 162728 69624
rect 166080 69572 166132 69624
rect 166724 69572 166776 69624
rect 194784 69572 194836 69624
rect 178868 69504 178920 69556
rect 210332 69504 210384 69556
rect 210700 69504 210752 69556
rect 166724 69436 166776 69488
rect 186872 69436 186924 69488
rect 140044 69028 140096 69080
rect 142160 69028 142212 69080
rect 110052 68960 110104 69012
rect 143908 68960 143960 69012
rect 155040 68960 155092 69012
rect 155868 68960 155920 69012
rect 197820 68960 197872 69012
rect 100760 68892 100812 68944
rect 101588 68892 101640 68944
rect 135628 68892 135680 68944
rect 163228 68892 163280 68944
rect 163872 68892 163924 68944
rect 164700 68892 164752 68944
rect 165436 68892 165488 68944
rect 165988 68892 166040 68944
rect 166816 68892 166868 68944
rect 167368 68892 167420 68944
rect 168196 68892 168248 68944
rect 202236 68892 202288 68944
rect 108764 68824 108816 68876
rect 142160 68824 142212 68876
rect 142712 68824 142764 68876
rect 167460 68824 167512 68876
rect 168104 68824 168156 68876
rect 202144 68824 202196 68876
rect 108948 68756 109000 68808
rect 142896 68756 142948 68808
rect 166816 68756 166868 68808
rect 200580 68756 200632 68808
rect 112536 68688 112588 68740
rect 144092 68688 144144 68740
rect 168748 68688 168800 68740
rect 169392 68688 169444 68740
rect 203340 68688 203392 68740
rect 106832 68620 106884 68672
rect 138020 68620 138072 68672
rect 138572 68620 138624 68672
rect 175924 68620 175976 68672
rect 199844 68620 199896 68672
rect 102140 68552 102192 68604
rect 103060 68552 103112 68604
rect 134248 68552 134300 68604
rect 163872 68552 163924 68604
rect 198280 68552 198332 68604
rect 114008 68484 114060 68536
rect 144000 68484 144052 68536
rect 160192 68484 160244 68536
rect 194600 68484 194652 68536
rect 195060 68484 195112 68536
rect 102232 68416 102284 68468
rect 132776 68416 132828 68468
rect 165436 68416 165488 68468
rect 175924 68416 175976 68468
rect 176568 68416 176620 68468
rect 210424 68416 210476 68468
rect 116216 68348 116268 68400
rect 141424 68348 141476 68400
rect 164608 68348 164660 68400
rect 189080 68348 189132 68400
rect 48320 68280 48372 68332
rect 100760 68280 100812 68332
rect 110788 68280 110840 68332
rect 120172 68280 120224 68332
rect 141240 68280 141292 68332
rect 160284 68280 160336 68332
rect 161112 68280 161164 68332
rect 184388 68280 184440 68332
rect 195060 68280 195112 68332
rect 358820 68280 358872 68332
rect 175832 68212 175884 68264
rect 176568 68212 176620 68264
rect 177580 68212 177632 68264
rect 200764 68212 200816 68264
rect 201408 68212 201460 68264
rect 189080 67736 189132 67788
rect 422944 67736 422996 67788
rect 188436 67668 188488 67720
rect 507860 67668 507912 67720
rect 141424 67600 141476 67652
rect 142252 67600 142304 67652
rect 144092 67600 144144 67652
rect 144368 67600 144420 67652
rect 201408 67600 201460 67652
rect 536840 67600 536892 67652
rect 99288 67532 99340 67584
rect 132684 67532 132736 67584
rect 133236 67532 133288 67584
rect 150624 67532 150676 67584
rect 151084 67532 151136 67584
rect 172612 67532 172664 67584
rect 212908 67532 212960 67584
rect 213828 67532 213880 67584
rect 108856 67464 108908 67516
rect 135260 67464 135312 67516
rect 142620 67464 142672 67516
rect 172796 67464 172848 67516
rect 173624 67464 173676 67516
rect 174268 67464 174320 67516
rect 174728 67464 174780 67516
rect 175648 67464 175700 67516
rect 215576 67464 215628 67516
rect 120356 67396 120408 67448
rect 151912 67396 151964 67448
rect 152556 67396 152608 67448
rect 172704 67396 172756 67448
rect 173440 67396 173492 67448
rect 174176 67396 174228 67448
rect 175004 67396 175056 67448
rect 175740 67396 175792 67448
rect 176292 67396 176344 67448
rect 117596 67328 117648 67380
rect 149152 67328 149204 67380
rect 174084 67328 174136 67380
rect 174820 67328 174872 67380
rect 175556 67328 175608 67380
rect 176476 67328 176528 67380
rect 104532 67260 104584 67312
rect 136088 67260 136140 67312
rect 175004 67260 175056 67312
rect 208952 67396 209004 67448
rect 177212 67328 177264 67380
rect 207480 67328 207532 67380
rect 80060 66852 80112 66904
rect 107292 67192 107344 67244
rect 138296 67192 138348 67244
rect 174820 67192 174872 67244
rect 208768 67260 208820 67312
rect 177120 67192 177172 67244
rect 207296 67192 207348 67244
rect 108304 67124 108356 67176
rect 138848 67124 138900 67176
rect 122472 67056 122524 67108
rect 150624 67124 150676 67176
rect 176476 67124 176528 67176
rect 210056 67124 210108 67176
rect 149152 67056 149204 67108
rect 149888 67056 149940 67108
rect 154396 67056 154448 67108
rect 274640 67056 274692 67108
rect 162492 66988 162544 67040
rect 189448 66988 189500 67040
rect 317420 66988 317472 67040
rect 176292 66920 176344 66972
rect 209964 66920 210016 66972
rect 213828 66920 213880 66972
rect 529940 66920 529992 66972
rect 147864 66852 147916 66904
rect 203524 66852 203576 66904
rect 215576 66852 215628 66904
rect 545764 66852 545816 66904
rect 153476 66784 153528 66836
rect 154488 66784 154540 66836
rect 174728 66784 174780 66836
rect 207388 66784 207440 66836
rect 173624 66716 173676 66768
rect 177120 66716 177172 66768
rect 173440 66648 173492 66700
rect 177212 66648 177264 66700
rect 144000 66512 144052 66564
rect 147220 66512 147272 66564
rect 141516 66240 141568 66292
rect 142344 66240 142396 66292
rect 100760 66172 100812 66224
rect 101680 66172 101732 66224
rect 134340 66172 134392 66224
rect 161756 66172 161808 66224
rect 162492 66172 162544 66224
rect 164516 66172 164568 66224
rect 165252 66172 165304 66224
rect 168656 66172 168708 66224
rect 169576 66172 169628 66224
rect 100024 66104 100076 66156
rect 134156 66104 134208 66156
rect 142344 66104 142396 66156
rect 142988 66104 143040 66156
rect 210148 66172 210200 66224
rect 170220 66104 170272 66156
rect 209044 66104 209096 66156
rect 100116 66036 100168 66088
rect 134064 66036 134116 66088
rect 134800 66036 134852 66088
rect 161664 66036 161716 66088
rect 162584 66036 162636 66088
rect 165252 66036 165304 66088
rect 205824 66036 205876 66088
rect 102692 65968 102744 66020
rect 135536 65968 135588 66020
rect 165896 65968 165948 66020
rect 200304 65968 200356 66020
rect 201408 65968 201460 66020
rect 99472 65900 99524 65952
rect 100484 65900 100536 65952
rect 133052 65900 133104 65952
rect 154948 65900 155000 65952
rect 189080 65900 189132 65952
rect 119712 65832 119764 65884
rect 150532 65832 150584 65884
rect 162584 65832 162636 65884
rect 170220 65832 170272 65884
rect 185584 65832 185636 65884
rect 214840 65832 214892 65884
rect 108948 65764 109000 65816
rect 140136 65764 140188 65816
rect 177028 65764 177080 65816
rect 203616 65764 203668 65816
rect 204168 65764 204220 65816
rect 124128 65696 124180 65748
rect 161572 65696 161624 65748
rect 162124 65696 162176 65748
rect 169576 65696 169628 65748
rect 186780 65696 186832 65748
rect 238760 65696 238812 65748
rect 149428 65628 149480 65680
rect 223580 65628 223632 65680
rect 35992 65560 36044 65612
rect 100760 65560 100812 65612
rect 189080 65560 189132 65612
rect 295340 65560 295392 65612
rect 8300 65492 8352 65544
rect 99472 65492 99524 65544
rect 112168 65492 112220 65544
rect 131488 65492 131540 65544
rect 141148 65492 141200 65544
rect 201408 65492 201460 65544
rect 432604 65492 432656 65544
rect 150532 65424 150584 65476
rect 151268 65424 151320 65476
rect 142528 65356 142580 65408
rect 142804 65356 142856 65408
rect 204168 64880 204220 64932
rect 570604 64880 570656 64932
rect 104256 64812 104308 64864
rect 137468 64812 137520 64864
rect 165712 64812 165764 64864
rect 200856 64812 200908 64864
rect 104624 64744 104676 64796
rect 137100 64744 137152 64796
rect 153108 64744 153160 64796
rect 186596 64744 186648 64796
rect 165344 64676 165396 64728
rect 199936 64676 199988 64728
rect 166540 64608 166592 64660
rect 200396 64608 200448 64660
rect 158996 64540 159048 64592
rect 193312 64540 193364 64592
rect 168564 64472 168616 64524
rect 202880 64472 202932 64524
rect 171416 64404 171468 64456
rect 187148 64404 187200 64456
rect 186596 64336 186648 64388
rect 256700 64336 256752 64388
rect 149612 64268 149664 64320
rect 220084 64268 220136 64320
rect 193312 64200 193364 64252
rect 345020 64200 345072 64252
rect 62120 64132 62172 64184
rect 104624 64132 104676 64184
rect 146852 64132 146904 64184
rect 183560 64132 183612 64184
rect 202880 64132 202932 64184
rect 472624 64132 472676 64184
rect 165804 63996 165856 64048
rect 166540 63996 166592 64048
rect 164424 63860 164476 63912
rect 165344 63860 165396 63912
rect 146024 63588 146076 63640
rect 149796 63588 149848 63640
rect 165712 63520 165764 63572
rect 166448 63520 166500 63572
rect 187148 63520 187200 63572
rect 512000 63520 512052 63572
rect 164332 63452 164384 63504
rect 199016 63452 199068 63504
rect 199200 63452 199252 63504
rect 143816 63384 143868 63436
rect 148416 63384 148468 63436
rect 154764 63384 154816 63436
rect 189080 63384 189132 63436
rect 151728 62908 151780 62960
rect 245660 62908 245712 62960
rect 189080 62840 189132 62892
rect 190000 62840 190052 62892
rect 292580 62840 292632 62892
rect 199200 62772 199252 62824
rect 412640 62772 412692 62824
rect 102232 62024 102284 62076
rect 103336 62024 103388 62076
rect 136180 62024 136232 62076
rect 167276 62024 167328 62076
rect 202052 62024 202104 62076
rect 202788 62024 202840 62076
rect 102140 61956 102192 62008
rect 102692 61956 102744 62008
rect 134432 61956 134484 62008
rect 156144 61956 156196 62008
rect 190552 61956 190604 62008
rect 191748 61956 191800 62008
rect 163044 61888 163096 61940
rect 197360 61888 197412 61940
rect 175464 61820 175516 61872
rect 199108 61820 199160 61872
rect 148968 61616 149020 61668
rect 197636 61616 197688 61668
rect 191748 61548 191800 61600
rect 313280 61548 313332 61600
rect 154212 61480 154264 61532
rect 277400 61480 277452 61532
rect 197360 61412 197412 61464
rect 398840 61412 398892 61464
rect 43444 61344 43496 61396
rect 102232 61344 102284 61396
rect 202788 61344 202840 61396
rect 459560 61344 459612 61396
rect 199108 60732 199160 60784
rect 563704 60732 563756 60784
rect 98920 60664 98972 60716
rect 132960 60664 133012 60716
rect 154672 60664 154724 60716
rect 214196 60664 214248 60716
rect 214472 60664 214524 60716
rect 102140 60596 102192 60648
rect 103428 60596 103480 60648
rect 135720 60596 135772 60648
rect 158904 60596 158956 60648
rect 193404 60596 193456 60648
rect 194508 60596 194560 60648
rect 111800 60528 111852 60580
rect 112260 60528 112312 60580
rect 139860 60528 139912 60580
rect 166356 60528 166408 60580
rect 196256 60528 196308 60580
rect 214472 60120 214524 60172
rect 299480 60120 299532 60172
rect 44180 60052 44232 60104
rect 102140 60052 102192 60104
rect 194508 60052 194560 60104
rect 351920 60052 351972 60104
rect 21364 59984 21416 60036
rect 98920 59984 98972 60036
rect 196256 59984 196308 60036
rect 196900 59984 196952 60036
rect 402980 59984 403032 60036
rect 3516 59304 3568 59356
rect 40684 59304 40736 59356
rect 109868 59304 109920 59356
rect 110420 59304 110472 59356
rect 104164 59168 104216 59220
rect 135812 59304 135864 59356
rect 161480 59304 161532 59356
rect 196256 59304 196308 59356
rect 196532 59304 196584 59356
rect 106004 59100 106056 59152
rect 106188 59100 106240 59152
rect 137008 59236 137060 59288
rect 157432 59236 157484 59288
rect 192116 59236 192168 59288
rect 193036 59236 193088 59288
rect 148692 58896 148744 58948
rect 198740 58896 198792 58948
rect 151636 58828 151688 58880
rect 249800 58828 249852 58880
rect 154120 58760 154172 58812
rect 281540 58760 281592 58812
rect 193036 58692 193088 58744
rect 327080 58692 327132 58744
rect 69020 58624 69072 58676
rect 106004 58624 106056 58676
rect 196256 58624 196308 58676
rect 380900 58624 380952 58676
rect 158812 57876 158864 57928
rect 193220 57876 193272 57928
rect 194508 57876 194560 57928
rect 170128 57808 170180 57860
rect 196256 57808 196308 57860
rect 194508 57196 194560 57248
rect 349160 57196 349212 57248
rect 196256 56584 196308 56636
rect 484400 56584 484452 56636
rect 113548 56516 113600 56568
rect 138388 56516 138440 56568
rect 167184 56516 167236 56568
rect 201592 56516 201644 56568
rect 202788 56516 202840 56568
rect 145104 55836 145156 55888
rect 170404 55836 170456 55888
rect 202788 55836 202840 55888
rect 450544 55836 450596 55888
rect 138664 55224 138716 55276
rect 142344 55224 142396 55276
rect 156052 55156 156104 55208
rect 190460 55156 190512 55208
rect 191748 55156 191800 55208
rect 176936 55088 176988 55140
rect 203340 55088 203392 55140
rect 167920 55020 167972 55072
rect 189356 55020 189408 55072
rect 151544 54612 151596 54664
rect 239404 54612 239456 54664
rect 191748 54544 191800 54596
rect 315304 54544 315356 54596
rect 189356 54476 189408 54528
rect 382280 54476 382332 54528
rect 203984 53796 204036 53848
rect 571984 53796 572036 53848
rect 162952 53728 163004 53780
rect 198372 53728 198424 53780
rect 172520 53660 172572 53712
rect 207204 53660 207256 53712
rect 165620 53592 165672 53644
rect 198924 53592 198976 53644
rect 199108 53592 199160 53644
rect 198372 53184 198424 53236
rect 391940 53184 391992 53236
rect 199108 53116 199160 53168
rect 437480 53116 437532 53168
rect 145748 53048 145800 53100
rect 163504 53048 163556 53100
rect 207204 53048 207256 53100
rect 516784 53048 516836 53100
rect 158720 52368 158772 52420
rect 193220 52368 193272 52420
rect 194508 52368 194560 52420
rect 162860 52300 162912 52352
rect 197544 52300 197596 52352
rect 198096 52300 198148 52352
rect 168380 52232 168432 52284
rect 201960 52232 202012 52284
rect 202788 52232 202840 52284
rect 143724 51688 143776 51740
rect 157432 51688 157484 51740
rect 198096 51688 198148 51740
rect 400864 51688 400916 51740
rect 194508 51144 194560 51196
rect 356060 51144 356112 51196
rect 202788 51076 202840 51128
rect 464344 51076 464396 51128
rect 176844 51008 176896 51060
rect 207204 51008 207256 51060
rect 150348 50328 150400 50380
rect 225604 50328 225656 50380
rect 207204 49716 207256 49768
rect 569960 49716 570012 49768
rect 167000 49648 167052 49700
rect 201868 49648 201920 49700
rect 202788 49648 202840 49700
rect 147404 49172 147456 49224
rect 186320 49172 186372 49224
rect 150256 49104 150308 49156
rect 222200 49104 222252 49156
rect 147772 49036 147824 49088
rect 201592 49036 201644 49088
rect 202788 49036 202840 49088
rect 448612 49036 448664 49088
rect 133972 48968 134024 49020
rect 142528 48968 142580 49020
rect 145012 48968 145064 49020
rect 168380 48968 168432 49020
rect 172060 48968 172112 49020
rect 502984 48968 503036 49020
rect 144368 48220 144420 48272
rect 147680 48220 147732 48272
rect 147772 47676 147824 47728
rect 208400 47676 208452 47728
rect 150164 47608 150216 47660
rect 215300 47608 215352 47660
rect 169300 47540 169352 47592
rect 468484 47540 468536 47592
rect 154580 46860 154632 46912
rect 216772 46860 216824 46912
rect 217048 46860 217100 46912
rect 176752 46792 176804 46844
rect 207204 46792 207256 46844
rect 145656 46180 145708 46232
rect 167000 46180 167052 46232
rect 216772 46180 216824 46232
rect 292672 46180 292724 46232
rect 207940 45568 207992 45620
rect 560944 45568 560996 45620
rect 152924 44820 152976 44872
rect 267740 44820 267792 44872
rect 177396 44072 177448 44124
rect 211252 44072 211304 44124
rect 212448 44072 212500 44124
rect 151452 43460 151504 43512
rect 233240 43460 233292 43512
rect 212448 43392 212500 43444
rect 578240 43392 578292 43444
rect 149060 42304 149112 42356
rect 218152 42304 218204 42356
rect 155316 42236 155368 42288
rect 285680 42236 285732 42288
rect 165068 42168 165120 42220
rect 426440 42168 426492 42220
rect 170036 42100 170088 42152
rect 495440 42100 495492 42152
rect 70400 42032 70452 42084
rect 136916 42032 136968 42084
rect 172152 42032 172204 42084
rect 503720 42032 503772 42084
rect 148600 41012 148652 41064
rect 204352 41012 204404 41064
rect 156696 40944 156748 40996
rect 309140 40944 309192 40996
rect 158352 40876 158404 40928
rect 332692 40876 332744 40928
rect 169944 40808 169996 40860
rect 491300 40808 491352 40860
rect 171324 40740 171376 40792
rect 498292 40740 498344 40792
rect 74540 40672 74592 40724
rect 138112 40672 138164 40724
rect 174728 40672 174780 40724
rect 549260 40672 549312 40724
rect 138112 39992 138164 40044
rect 142252 39992 142304 40044
rect 150440 39584 150492 39636
rect 236000 39584 236052 39636
rect 158260 39516 158312 39568
rect 324412 39516 324464 39568
rect 169392 39448 169444 39500
rect 463700 39448 463752 39500
rect 167092 39380 167144 39432
rect 462320 39380 462372 39432
rect 77392 39312 77444 39364
rect 138020 39312 138072 39364
rect 173532 39312 173584 39364
rect 516140 39312 516192 39364
rect 145564 38156 145616 38208
rect 168564 38156 168616 38208
rect 153016 38088 153068 38140
rect 251272 38088 251324 38140
rect 169484 38020 169536 38072
rect 470600 38020 470652 38072
rect 168472 37952 168524 38004
rect 476120 37952 476172 38004
rect 13820 37884 13872 37936
rect 132868 37884 132920 37936
rect 174912 37884 174964 37936
rect 534080 37884 534132 37936
rect 154028 36660 154080 36712
rect 267832 36660 267884 36712
rect 170864 36592 170916 36644
rect 481640 36592 481692 36644
rect 95240 36524 95292 36576
rect 139584 36524 139636 36576
rect 173440 36524 173492 36576
rect 527824 36524 527876 36576
rect 158444 35368 158496 35420
rect 321560 35368 321612 35420
rect 166448 35300 166500 35352
rect 440332 35300 440384 35352
rect 174820 35232 174872 35284
rect 538864 35232 538916 35284
rect 23480 35164 23532 35216
rect 134156 35164 134208 35216
rect 176384 35164 176436 35216
rect 558920 35164 558972 35216
rect 160836 33940 160888 33992
rect 357440 33940 357492 33992
rect 162124 33872 162176 33924
rect 378784 33872 378836 33924
rect 169852 33804 169904 33856
rect 488540 33804 488592 33856
rect 31760 33736 31812 33788
rect 134064 33736 134116 33788
rect 144276 33736 144328 33788
rect 160100 33736 160152 33788
rect 177672 33736 177724 33788
rect 576860 33736 576912 33788
rect 3516 33056 3568 33108
rect 97264 33056 97316 33108
rect 148508 32648 148560 32700
rect 205732 32648 205784 32700
rect 152832 32580 152884 32632
rect 264980 32580 265032 32632
rect 159732 32512 159784 32564
rect 346400 32512 346452 32564
rect 163780 32444 163832 32496
rect 404360 32444 404412 32496
rect 170956 32376 171008 32428
rect 492680 32376 492732 32428
rect 155776 31288 155828 31340
rect 299572 31288 299624 31340
rect 160928 31220 160980 31272
rect 360200 31220 360252 31272
rect 163872 31152 163924 31204
rect 407212 31152 407264 31204
rect 184296 31084 184348 31136
rect 561680 31084 561732 31136
rect 42800 31016 42852 31068
rect 135536 31016 135588 31068
rect 176292 31016 176344 31068
rect 564532 31016 564584 31068
rect 150072 29928 150124 29980
rect 229100 29928 229152 29980
rect 156972 29860 157024 29912
rect 303620 29860 303672 29912
rect 165160 29792 165212 29844
rect 409880 29792 409932 29844
rect 169576 29724 169628 29776
rect 474740 29724 474792 29776
rect 171232 29656 171284 29708
rect 502340 29656 502392 29708
rect 177764 29588 177816 29640
rect 574100 29588 574152 29640
rect 151360 28500 151412 28552
rect 242992 28500 243044 28552
rect 159824 28432 159876 28484
rect 339500 28432 339552 28484
rect 161020 28364 161072 28416
rect 360844 28364 360896 28416
rect 166632 28296 166684 28348
rect 438860 28296 438912 28348
rect 172428 28228 172480 28280
rect 506572 28228 506624 28280
rect 154396 27072 154448 27124
rect 275284 27072 275336 27124
rect 162308 27004 162360 27056
rect 374092 27004 374144 27056
rect 171140 26936 171192 26988
rect 509240 26936 509292 26988
rect 172244 26868 172296 26920
rect 510620 26868 510672 26920
rect 153292 25712 153344 25764
rect 278780 25712 278832 25764
rect 144184 25644 144236 25696
rect 144920 25644 144972 25696
rect 162400 25644 162452 25696
rect 378140 25644 378192 25696
rect 172336 25576 172388 25628
rect 513380 25576 513432 25628
rect 146024 25508 146076 25560
rect 171784 25508 171836 25560
rect 173624 25508 173676 25560
rect 531412 25508 531464 25560
rect 153200 24352 153252 24404
rect 282920 24352 282972 24404
rect 163964 24284 164016 24336
rect 396080 24284 396132 24336
rect 165252 24216 165304 24268
rect 425060 24216 425112 24268
rect 173808 24148 173860 24200
rect 520280 24148 520332 24200
rect 175004 24080 175056 24132
rect 546500 24080 546552 24132
rect 157064 22924 157116 22976
rect 310520 22924 310572 22976
rect 164056 22856 164108 22908
rect 398932 22856 398984 22908
rect 173716 22788 173768 22840
rect 527180 22788 527232 22840
rect 176476 22720 176528 22772
rect 552664 22720 552716 22772
rect 166540 21360 166592 21412
rect 431960 21360 432012 21412
rect 574744 20612 574796 20664
rect 580172 20612 580224 20664
rect 153844 20136 153896 20188
rect 280160 20136 280212 20188
rect 155868 20068 155920 20120
rect 287060 20068 287112 20120
rect 155224 20000 155276 20052
rect 291200 20000 291252 20052
rect 144828 19932 144880 19984
rect 154580 19932 154632 19984
rect 161112 19932 161164 19984
rect 357532 19932 357584 19984
rect 152740 18776 152792 18828
rect 266360 18776 266412 18828
rect 157340 18708 157392 18760
rect 329840 18708 329892 18760
rect 176568 18640 176620 18692
rect 567200 18640 567252 18692
rect 177856 18572 177908 18624
rect 571340 18572 571392 18624
rect 149980 17416 150032 17468
rect 219440 17416 219492 17468
rect 168104 17348 168156 17400
rect 445760 17348 445812 17400
rect 169208 17280 169260 17332
rect 477500 17280 477552 17332
rect 177948 17212 178000 17264
rect 518900 17212 518952 17264
rect 151268 16056 151320 16108
rect 248420 16056 248472 16108
rect 161204 15988 161256 16040
rect 364616 15988 364668 16040
rect 165436 15920 165488 15972
rect 420920 15920 420972 15972
rect 87512 15852 87564 15904
rect 138204 15852 138256 15904
rect 166724 15852 166776 15904
rect 442172 15852 442224 15904
rect 153936 14696 153988 14748
rect 272432 14696 272484 14748
rect 155960 14628 156012 14680
rect 314660 14628 314712 14680
rect 162768 14560 162820 14612
rect 385960 14560 386012 14612
rect 165344 14492 165396 14544
rect 411904 14492 411956 14544
rect 169760 14424 169812 14476
rect 486424 14424 486476 14476
rect 152648 13336 152700 13388
rect 258264 13336 258316 13388
rect 157156 13268 157208 13320
rect 307944 13268 307996 13320
rect 162676 13200 162728 13252
rect 382372 13200 382424 13252
rect 162492 13132 162544 13184
rect 390652 13132 390704 13184
rect 171048 13064 171100 13116
rect 482192 13064 482244 13116
rect 151176 11976 151228 12028
rect 245200 11976 245252 12028
rect 158536 11908 158588 11960
rect 328736 11908 328788 11960
rect 164148 11840 164200 11892
rect 376024 11840 376076 11892
rect 164240 11772 164292 11824
rect 417424 11772 417476 11824
rect 143540 11704 143592 11756
rect 144736 11704 144788 11756
rect 175096 11704 175148 11756
rect 545488 11704 545540 11756
rect 184940 11636 184992 11688
rect 186136 11636 186188 11688
rect 234620 11636 234672 11688
rect 235816 11636 235868 11688
rect 151084 10548 151136 10600
rect 241704 10548 241756 10600
rect 158628 10480 158680 10532
rect 336280 10480 336332 10532
rect 162584 10412 162636 10464
rect 386696 10412 386748 10464
rect 166816 10344 166868 10396
rect 432052 10344 432104 10396
rect 175188 10276 175240 10328
rect 548432 10276 548484 10328
rect 157248 9052 157300 9104
rect 316224 9052 316276 9104
rect 165528 8984 165580 9036
rect 414296 8984 414348 9036
rect 52552 8916 52604 8968
rect 135352 8916 135404 8968
rect 175372 8916 175424 8968
rect 556160 8916 556212 8968
rect 142804 8236 142856 8288
rect 143540 8236 143592 8288
rect 149888 7828 149940 7880
rect 227536 7828 227588 7880
rect 159916 7760 159968 7812
rect 343364 7760 343416 7812
rect 161296 7692 161348 7744
rect 365812 7692 365864 7744
rect 166908 7624 166960 7676
rect 435548 7624 435600 7676
rect 25320 7556 25372 7608
rect 133880 7556 133932 7608
rect 173992 7556 174044 7608
rect 538404 7556 538456 7608
rect 152556 6536 152608 6588
rect 259552 6536 259604 6588
rect 160008 6468 160060 6520
rect 350448 6468 350500 6520
rect 179144 6400 179196 6452
rect 443828 6400 443880 6452
rect 180616 6332 180668 6384
rect 450912 6332 450964 6384
rect 168196 6264 168248 6316
rect 453304 6264 453356 6316
rect 176200 6196 176252 6248
rect 563244 6196 563296 6248
rect 103336 6128 103388 6180
rect 139768 6128 139820 6180
rect 182088 6128 182140 6180
rect 583392 6128 583444 6180
rect 154488 4972 154540 5024
rect 273628 4972 273680 5024
rect 161388 4904 161440 4956
rect 371700 4904 371752 4956
rect 168288 4836 168340 4888
rect 456892 4836 456944 4888
rect 6460 4768 6512 4820
rect 132684 4768 132736 4820
rect 173900 4768 173952 4820
rect 541992 4768 542044 4820
rect 572 4088 624 4140
rect 7564 4088 7616 4140
rect 73804 4088 73856 4140
rect 75184 4088 75236 4140
rect 112812 4088 112864 4140
rect 113824 4088 113876 4140
rect 141240 4088 141292 4140
rect 142344 4088 142396 4140
rect 149704 4088 149756 4140
rect 153016 4088 153068 4140
rect 189816 4088 189868 4140
rect 203892 4088 203944 4140
rect 211804 4088 211856 4140
rect 217324 4088 217376 4140
rect 229744 4088 229796 4140
rect 230940 4088 230992 4140
rect 181444 4020 181496 4072
rect 190828 4020 190880 4072
rect 193864 4020 193916 4072
rect 195612 4020 195664 4072
rect 195704 4020 195756 4072
rect 216496 4020 216548 4072
rect 216680 4020 216732 4072
rect 247592 4088 247644 4140
rect 247684 4088 247736 4140
rect 254676 4088 254728 4140
rect 315304 4088 315356 4140
rect 317328 4088 317380 4140
rect 323584 4088 323636 4140
rect 326804 4088 326856 4140
rect 450544 4088 450596 4140
rect 452108 4088 452160 4140
rect 486516 4088 486568 4140
rect 489920 4088 489972 4140
rect 527916 4088 527968 4140
rect 529020 4088 529072 4140
rect 251180 4020 251232 4072
rect 252376 4020 252428 4072
rect 181536 3952 181588 4004
rect 212172 3952 212224 4004
rect 217324 3952 217376 4004
rect 231032 3952 231084 4004
rect 231124 3952 231176 4004
rect 298468 3952 298520 4004
rect 299572 3952 299624 4004
rect 300768 3952 300820 4004
rect 311164 3952 311216 4004
rect 312636 3952 312688 4004
rect 360844 3952 360896 4004
rect 362316 3952 362368 4004
rect 122288 3680 122340 3732
rect 127072 3884 127124 3936
rect 152464 3884 152516 3936
rect 161388 3884 161440 3936
rect 178684 3884 178736 3936
rect 401324 3884 401376 3936
rect 65524 3612 65576 3664
rect 17040 3544 17092 3596
rect 18604 3544 18656 3596
rect 19432 3544 19484 3596
rect 21364 3544 21416 3596
rect 27620 3544 27672 3596
rect 28540 3544 28592 3596
rect 51356 3544 51408 3596
rect 54484 3544 54536 3596
rect 56048 3544 56100 3596
rect 57244 3544 57296 3596
rect 60740 3544 60792 3596
rect 61660 3544 61712 3596
rect 69112 3544 69164 3596
rect 71044 3544 71096 3596
rect 83280 3612 83332 3664
rect 131304 3816 131356 3868
rect 132960 3816 133012 3868
rect 140044 3816 140096 3868
rect 146944 3816 146996 3868
rect 149612 3816 149664 3868
rect 149796 3816 149848 3868
rect 163688 3816 163740 3868
rect 170404 3816 170456 3868
rect 173164 3816 173216 3868
rect 178776 3816 178828 3868
rect 408408 3816 408460 3868
rect 129832 3748 129884 3800
rect 131028 3748 131080 3800
rect 150624 3748 150676 3800
rect 160100 3748 160152 3800
rect 161296 3748 161348 3800
rect 161388 3748 161440 3800
rect 171968 3748 172020 3800
rect 179328 3748 179380 3800
rect 429660 3748 429712 3800
rect 15936 3476 15988 3528
rect 130844 3680 130896 3732
rect 162492 3680 162544 3732
rect 131396 3612 131448 3664
rect 137652 3612 137704 3664
rect 138664 3612 138716 3664
rect 147036 3612 147088 3664
rect 149520 3612 149572 3664
rect 149612 3612 149664 3664
rect 170772 3680 170824 3732
rect 179236 3680 179288 3732
rect 436744 3680 436796 3732
rect 442264 3680 442316 3732
rect 497096 3680 497148 3732
rect 125876 3544 125928 3596
rect 129924 3544 129976 3596
rect 130936 3544 130988 3596
rect 166080 3612 166132 3664
rect 179052 3612 179104 3664
rect 447416 3612 447468 3664
rect 163504 3544 163556 3596
rect 164884 3544 164936 3596
rect 168380 3544 168432 3596
rect 169576 3544 169628 3596
rect 186228 3544 186280 3596
rect 468300 3544 468352 3596
rect 468484 3544 468536 3596
rect 469864 3544 469916 3596
rect 123484 3476 123536 3528
rect 124864 3476 124916 3528
rect 128176 3476 128228 3528
rect 129004 3476 129056 3528
rect 140044 3476 140096 3528
rect 141516 3476 141568 3528
rect 147220 3476 147272 3528
rect 175464 3476 175516 3528
rect 180708 3476 180760 3528
rect 472624 3476 472676 3528
rect 473452 3476 473504 3528
rect 478236 3544 478288 3596
rect 498200 3544 498252 3596
rect 516784 3544 516836 3596
rect 518348 3544 518400 3596
rect 479340 3476 479392 3528
rect 482284 3476 482336 3528
rect 507676 3476 507728 3528
rect 526444 3476 526496 3528
rect 533712 3476 533764 3528
rect 538864 3476 538916 3528
rect 539600 3476 539652 3528
rect 540244 3476 540296 3528
rect 547880 3476 547932 3528
rect 552756 3476 552808 3528
rect 560852 3476 560904 3528
rect 563704 3476 563756 3528
rect 565636 3476 565688 3528
rect 567844 3476 567896 3528
rect 569132 3476 569184 3528
rect 1676 3408 1728 3460
rect 8944 3408 8996 3460
rect 11152 3408 11204 3460
rect 91560 3340 91612 3392
rect 93124 3340 93176 3392
rect 101036 3340 101088 3392
rect 102876 3340 102928 3392
rect 105728 3340 105780 3392
rect 106924 3340 106976 3392
rect 111616 3340 111668 3392
rect 112444 3340 112496 3392
rect 120080 3340 120132 3392
rect 120724 3340 120776 3392
rect 148324 3408 148376 3460
rect 176660 3408 176712 3460
rect 180524 3408 180576 3460
rect 487620 3408 487672 3460
rect 498844 3408 498896 3460
rect 540796 3408 540848 3460
rect 545764 3408 545816 3460
rect 554964 3408 555016 3460
rect 560944 3408 560996 3460
rect 573916 3408 573968 3460
rect 131120 3340 131172 3392
rect 147312 3340 147364 3392
rect 151820 3340 151872 3392
rect 182824 3340 182876 3392
rect 193220 3340 193272 3392
rect 210424 3340 210476 3392
rect 218060 3340 218112 3392
rect 225604 3340 225656 3392
rect 226340 3340 226392 3392
rect 239404 3340 239456 3392
rect 240508 3340 240560 3392
rect 242164 3340 242216 3392
rect 242900 3340 242952 3392
rect 259460 3340 259512 3392
rect 260656 3340 260708 3392
rect 261484 3340 261536 3392
rect 262956 3340 263008 3392
rect 275284 3340 275336 3392
rect 276020 3340 276072 3392
rect 307024 3340 307076 3392
rect 309048 3340 309100 3392
rect 324412 3340 324464 3392
rect 325608 3340 325660 3392
rect 332600 3340 332652 3392
rect 333888 3340 333940 3392
rect 340880 3340 340932 3392
rect 342168 3340 342220 3392
rect 342904 3340 342956 3392
rect 344560 3340 344612 3392
rect 357532 3340 357584 3392
rect 358728 3340 358780 3392
rect 364984 3340 365036 3392
rect 367008 3340 367060 3392
rect 374092 3340 374144 3392
rect 375288 3340 375340 3392
rect 378784 3340 378836 3392
rect 379980 3340 380032 3392
rect 382280 3340 382332 3392
rect 383568 3340 383620 3392
rect 398932 3340 398984 3392
rect 400128 3340 400180 3392
rect 400864 3340 400916 3392
rect 402520 3340 402572 3392
rect 414664 3340 414716 3392
rect 416688 3340 416740 3392
rect 418804 3340 418856 3392
rect 420184 3340 420236 3392
rect 422944 3340 422996 3392
rect 424968 3340 425020 3392
rect 432604 3340 432656 3392
rect 434444 3340 434496 3392
rect 440240 3340 440292 3392
rect 441528 3340 441580 3392
rect 448612 3340 448664 3392
rect 449808 3340 449860 3392
rect 456800 3340 456852 3392
rect 458088 3340 458140 3392
rect 571984 3340 572036 3392
rect 576308 3340 576360 3392
rect 126980 3272 127032 3324
rect 128452 3272 128504 3324
rect 193128 3272 193180 3324
rect 195704 3272 195756 3324
rect 207756 3272 207808 3324
rect 210976 3272 211028 3324
rect 431960 3272 432012 3324
rect 433248 3272 433300 3324
rect 184204 3204 184256 3256
rect 189724 3204 189776 3256
rect 520924 3204 520976 3256
rect 524236 3204 524288 3256
rect 33600 3136 33652 3188
rect 35164 3136 35216 3188
rect 38384 3136 38436 3188
rect 39304 3136 39356 3188
rect 41880 3136 41932 3188
rect 43444 3136 43496 3188
rect 136456 3136 136508 3188
rect 141424 3136 141476 3188
rect 548524 3136 548576 3188
rect 551468 3136 551520 3188
rect 12348 3068 12400 3120
rect 17224 3068 17276 3120
rect 30104 3068 30156 3120
rect 32404 3068 32456 3120
rect 124680 3068 124732 3120
rect 131488 3068 131540 3120
rect 171876 3068 171928 3120
rect 174268 3068 174320 3120
rect 382924 3068 382976 3120
rect 384764 3068 384816 3120
rect 570604 3068 570656 3120
rect 572720 3068 572772 3120
rect 20628 3000 20680 3052
rect 22744 3000 22796 3052
rect 23020 3000 23072 3052
rect 25504 3000 25556 3052
rect 118792 3000 118844 3052
rect 121460 3000 121512 3052
rect 148416 3000 148468 3052
rect 154212 3000 154264 3052
rect 464344 3000 464396 3052
rect 466276 3000 466328 3052
rect 503076 3000 503128 3052
rect 505376 3000 505428 3052
rect 514024 3000 514076 3052
rect 515956 3000 516008 3052
rect 203524 2932 203576 2984
rect 207388 2932 207440 2984
rect 220084 2932 220136 2984
rect 225144 2932 225196 2984
rect 509884 2932 509936 2984
rect 514760 2932 514812 2984
rect 171784 2864 171836 2916
rect 177856 2864 177908 2916
rect 260104 2864 260156 2916
rect 261760 2864 261812 2916
rect 390560 1776 390612 1828
rect 391848 1776 391900 1828
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 700534 8156 703520
rect 24320 700602 24348 703520
rect 24308 700596 24360 700602
rect 24308 700538 24360 700544
rect 8116 700528 8168 700534
rect 8116 700470 8168 700476
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683262 3464 684247
rect 3424 683256 3476 683262
rect 3424 683198 3476 683204
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 3476 632088 3478 632097
rect 3422 632023 3478 632032
rect 3146 619168 3202 619177
rect 3146 619103 3202 619112
rect 3160 618322 3188 619103
rect 3148 618316 3200 618322
rect 3148 618258 3200 618264
rect 3238 606112 3294 606121
rect 3238 606047 3294 606056
rect 3252 605878 3280 606047
rect 3240 605872 3292 605878
rect 3240 605814 3292 605820
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 3436 565894 3464 566879
rect 3424 565888 3476 565894
rect 3424 565830 3476 565836
rect 3422 553888 3478 553897
rect 3422 553823 3478 553832
rect 3436 553450 3464 553823
rect 3424 553444 3476 553450
rect 3424 553386 3476 553392
rect 3422 527912 3478 527921
rect 3422 527847 3478 527856
rect 3436 527202 3464 527847
rect 3424 527196 3476 527202
rect 3424 527138 3476 527144
rect 3422 514856 3478 514865
rect 3422 514791 3424 514800
rect 3476 514791 3478 514800
rect 8944 514820 8996 514826
rect 3424 514762 3476 514768
rect 8944 514762 8996 514768
rect 3054 501800 3110 501809
rect 3054 501735 3110 501744
rect 3068 501022 3096 501735
rect 3056 501016 3108 501022
rect 3056 500958 3108 500964
rect 3422 475688 3478 475697
rect 3422 475623 3478 475632
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 2870 410544 2926 410553
rect 2870 410479 2926 410488
rect 2884 409902 2912 410479
rect 2872 409896 2924 409902
rect 2872 409838 2924 409844
rect 2778 371376 2834 371385
rect 2778 371311 2780 371320
rect 2832 371311 2834 371320
rect 2780 371282 2832 371288
rect 3146 358456 3202 358465
rect 3146 358391 3202 358400
rect 3160 357474 3188 358391
rect 3148 357468 3200 357474
rect 3148 357410 3200 357416
rect 3330 319288 3386 319297
rect 3330 319223 3386 319232
rect 3344 318850 3372 319223
rect 3332 318844 3384 318850
rect 3332 318786 3384 318792
rect 3054 267200 3110 267209
rect 3054 267135 3110 267144
rect 3068 266422 3096 267135
rect 3056 266416 3108 266422
rect 3056 266358 3108 266364
rect 3436 265674 3464 475623
rect 3514 462632 3570 462641
rect 3514 462567 3570 462576
rect 3528 462398 3556 462567
rect 3516 462392 3568 462398
rect 3516 462334 3568 462340
rect 3514 423600 3570 423609
rect 3514 423535 3570 423544
rect 3528 422346 3556 423535
rect 3516 422340 3568 422346
rect 3516 422282 3568 422288
rect 3516 397520 3568 397526
rect 3514 397488 3516 397497
rect 3568 397488 3570 397497
rect 3514 397423 3570 397432
rect 4804 371340 4856 371346
rect 4804 371282 4856 371288
rect 3514 345400 3570 345409
rect 3514 345335 3570 345344
rect 3528 345234 3556 345335
rect 3516 345228 3568 345234
rect 3516 345170 3568 345176
rect 3514 306232 3570 306241
rect 3514 306167 3570 306176
rect 3528 305046 3556 306167
rect 3516 305040 3568 305046
rect 3516 304982 3568 304988
rect 3514 293176 3570 293185
rect 3514 293111 3570 293120
rect 3528 292602 3556 293111
rect 3516 292596 3568 292602
rect 3516 292538 3568 292544
rect 4816 268394 4844 371282
rect 7564 345228 7616 345234
rect 7564 345170 7616 345176
rect 7576 271250 7604 345170
rect 8956 274038 8984 514762
rect 10324 357468 10376 357474
rect 10324 357410 10376 357416
rect 10336 289134 10364 357410
rect 10324 289128 10376 289134
rect 10324 289070 10376 289076
rect 40052 279478 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218072 703582 218836 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 40040 279472 40092 279478
rect 40040 279414 40092 279420
rect 8944 274032 8996 274038
rect 8944 273974 8996 273980
rect 7564 271244 7616 271250
rect 7564 271186 7616 271192
rect 71792 269890 71820 702986
rect 89180 700738 89208 703520
rect 89168 700732 89220 700738
rect 89168 700674 89220 700680
rect 105464 699718 105492 703520
rect 137848 700874 137876 703520
rect 154132 702434 154160 703520
rect 170324 702434 170352 703520
rect 153212 702406 154160 702434
rect 169772 702406 170352 702434
rect 137836 700868 137888 700874
rect 137836 700810 137888 700816
rect 152464 700392 152516 700398
rect 152464 700334 152516 700340
rect 148324 700324 148376 700330
rect 148324 700266 148376 700272
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 106924 699712 106976 699718
rect 106924 699654 106976 699660
rect 71780 269884 71832 269890
rect 71780 269826 71832 269832
rect 4804 268388 4856 268394
rect 4804 268330 4856 268336
rect 3424 265668 3476 265674
rect 3424 265610 3476 265616
rect 106936 264246 106964 699654
rect 146944 696992 146996 696998
rect 146944 696934 146996 696940
rect 143540 616888 143592 616894
rect 143540 616830 143592 616836
rect 142160 590708 142212 590714
rect 142160 590650 142212 590656
rect 139400 484424 139452 484430
rect 139400 484366 139452 484372
rect 138664 430636 138716 430642
rect 138664 430578 138716 430584
rect 135260 351960 135312 351966
rect 135260 351902 135312 351908
rect 134524 324352 134576 324358
rect 134524 324294 134576 324300
rect 133144 271924 133196 271930
rect 133144 271866 133196 271872
rect 113088 265192 113140 265198
rect 113088 265134 113140 265140
rect 112812 265056 112864 265062
rect 112812 264998 112864 265004
rect 106924 264240 106976 264246
rect 106924 264182 106976 264188
rect 3424 263084 3476 263090
rect 3424 263026 3476 263032
rect 2780 241256 2832 241262
rect 2780 241198 2832 241204
rect 2792 241097 2820 241198
rect 2778 241088 2834 241097
rect 2778 241023 2834 241032
rect 3436 201929 3464 263026
rect 3516 262472 3568 262478
rect 3516 262414 3568 262420
rect 3528 254153 3556 262414
rect 112534 262304 112590 262313
rect 112534 262239 112590 262248
rect 111064 261044 111116 261050
rect 111064 260986 111116 260992
rect 4804 260976 4856 260982
rect 4804 260918 4856 260924
rect 3514 254144 3570 254153
rect 3514 254079 3570 254088
rect 4816 241262 4844 260918
rect 7564 260364 7616 260370
rect 7564 260306 7616 260312
rect 4804 241256 4856 241262
rect 4804 241198 4856 241204
rect 7576 215150 7604 260306
rect 3516 215144 3568 215150
rect 3516 215086 3568 215092
rect 7564 215144 7616 215150
rect 7564 215086 7616 215092
rect 3528 214985 3556 215086
rect 3514 214976 3570 214985
rect 3514 214911 3570 214920
rect 3422 201920 3478 201929
rect 3422 201855 3478 201864
rect 107292 200592 107344 200598
rect 107292 200534 107344 200540
rect 104808 200524 104860 200530
rect 104808 200466 104860 200472
rect 103152 198076 103204 198082
rect 103152 198018 103204 198024
rect 97908 196648 97960 196654
rect 97908 196590 97960 196596
rect 3424 189032 3476 189038
rect 3424 188974 3476 188980
rect 3436 188873 3464 188974
rect 3422 188864 3478 188873
rect 3422 188799 3478 188808
rect 3514 162888 3570 162897
rect 3514 162823 3570 162832
rect 3146 149832 3202 149841
rect 3146 149767 3202 149776
rect 3160 149190 3188 149767
rect 3148 149184 3200 149190
rect 3148 149126 3200 149132
rect 3528 145586 3556 162823
rect 97264 153264 97316 153270
rect 97264 153206 97316 153212
rect 3516 145580 3568 145586
rect 3516 145522 3568 145528
rect 40684 142316 40736 142322
rect 40684 142258 40736 142264
rect 13084 140820 13136 140826
rect 13084 140762 13136 140768
rect 8942 139496 8998 139505
rect 8942 139431 8998 139440
rect 3424 138032 3476 138038
rect 3424 137974 3476 137980
rect 3240 137964 3292 137970
rect 3240 137906 3292 137912
rect 3252 136785 3280 137906
rect 3238 136776 3294 136785
rect 3238 136711 3294 136720
rect 3056 111444 3108 111450
rect 3056 111386 3108 111392
rect 3068 110673 3096 111386
rect 3054 110664 3110 110673
rect 3054 110599 3110 110608
rect 2778 77888 2834 77897
rect 2778 77823 2834 77832
rect 2792 6914 2820 77823
rect 2870 62792 2926 62801
rect 2870 62727 2926 62736
rect 2884 16574 2912 62727
rect 3436 19417 3464 137974
rect 8956 111450 8984 139431
rect 8944 111444 8996 111450
rect 8944 111386 8996 111392
rect 3516 85536 3568 85542
rect 3516 85478 3568 85484
rect 3528 84697 3556 85478
rect 3514 84688 3570 84697
rect 3514 84623 3570 84632
rect 6918 78024 6974 78033
rect 6918 77959 6974 77968
rect 4160 72480 4212 72486
rect 4160 72422 4212 72428
rect 3516 71732 3568 71738
rect 3516 71674 3568 71680
rect 3528 71641 3556 71674
rect 3514 71632 3570 71641
rect 3514 71567 3570 71576
rect 3516 59356 3568 59362
rect 3516 59298 3568 59304
rect 3528 58585 3556 59298
rect 3514 58576 3570 58585
rect 3514 58511 3570 58520
rect 3516 33108 3568 33114
rect 3516 33050 3568 33056
rect 3528 32473 3556 33050
rect 3514 32464 3570 32473
rect 3514 32399 3570 32408
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 4172 16574 4200 72422
rect 6932 16574 6960 77959
rect 7562 75168 7618 75177
rect 7562 75103 7618 75112
rect 2884 16546 3372 16574
rect 4172 16546 5304 16574
rect 6932 16546 7512 16574
rect 2792 6886 2912 6914
rect 572 4140 624 4146
rect 572 4082 624 4088
rect 584 480 612 4082
rect 1676 3460 1728 3466
rect 1676 3402 1728 3408
rect 1688 480 1716 3402
rect 2884 480 2912 6886
rect 3344 490 3372 16546
rect 3422 10296 3478 10305
rect 3422 10231 3478 10240
rect 3436 6497 3464 10231
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 3344 462 3740 490
rect 5276 480 5304 16546
rect 6460 4820 6512 4826
rect 6460 4762 6512 4768
rect 6472 480 6500 4762
rect 7484 3482 7512 16546
rect 7576 4146 7604 75103
rect 8944 73840 8996 73846
rect 8944 73782 8996 73788
rect 8300 65544 8352 65550
rect 8300 65486 8352 65492
rect 8312 16574 8340 65486
rect 8312 16546 8800 16574
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7484 3454 7696 3482
rect 7668 480 7696 3454
rect 8772 480 8800 16546
rect 8956 3466 8984 73782
rect 9680 72548 9732 72554
rect 9680 72490 9732 72496
rect 8944 3460 8996 3466
rect 8944 3402 8996 3408
rect 3712 354 3740 462
rect 4038 354 4150 480
rect 3712 326 4150 354
rect 4038 -960 4150 326
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 72490
rect 13096 71738 13124 140762
rect 20718 78160 20774 78169
rect 20718 78095 20774 78104
rect 13084 71732 13136 71738
rect 13084 71674 13136 71680
rect 17222 71088 17278 71097
rect 17222 71023 17278 71032
rect 12438 55856 12494 55865
rect 12438 55791 12494 55800
rect 12452 16574 12480 55791
rect 13820 37936 13872 37942
rect 13820 37878 13872 37884
rect 13832 16574 13860 37878
rect 12452 16546 13584 16574
rect 13832 16546 14320 16574
rect 11152 3460 11204 3466
rect 11152 3402 11204 3408
rect 11164 480 11192 3402
rect 12348 3120 12400 3126
rect 12348 3062 12400 3068
rect 12360 480 12388 3062
rect 13556 480 13584 16546
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 17040 3596 17092 3602
rect 17040 3538 17092 3544
rect 15936 3528 15988 3534
rect 15936 3470 15988 3476
rect 15948 480 15976 3470
rect 17052 480 17080 3538
rect 17236 3126 17264 71023
rect 18602 68232 18658 68241
rect 18602 68167 18658 68176
rect 17958 51776 18014 51785
rect 17958 51711 18014 51720
rect 17224 3120 17276 3126
rect 17224 3062 17276 3068
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 51711
rect 18616 3602 18644 68167
rect 20732 16574 20760 78095
rect 34518 76528 34574 76537
rect 34518 76463 34574 76472
rect 22742 73808 22798 73817
rect 22742 73743 22798 73752
rect 21364 60036 21416 60042
rect 21364 59978 21416 59984
rect 20732 16546 21312 16574
rect 18604 3596 18656 3602
rect 18604 3538 18656 3544
rect 19432 3596 19484 3602
rect 19432 3538 19484 3544
rect 19444 480 19472 3538
rect 21284 3482 21312 16546
rect 21376 3602 21404 59978
rect 21364 3596 21416 3602
rect 21364 3538 21416 3544
rect 21284 3454 21864 3482
rect 20628 3052 20680 3058
rect 20628 2994 20680 3000
rect 20640 480 20668 2994
rect 21836 480 21864 3454
rect 22756 3058 22784 73743
rect 27620 71052 27672 71058
rect 27620 70994 27672 71000
rect 26238 68368 26294 68377
rect 26238 68303 26294 68312
rect 25502 57216 25558 57225
rect 25502 57151 25558 57160
rect 23480 35216 23532 35222
rect 23480 35158 23532 35164
rect 23492 16574 23520 35158
rect 23492 16546 24256 16574
rect 22744 3052 22796 3058
rect 22744 2994 22796 3000
rect 23020 3052 23072 3058
rect 23020 2994 23072 3000
rect 23032 480 23060 2994
rect 24228 480 24256 16546
rect 25320 7608 25372 7614
rect 25320 7550 25372 7556
rect 25332 480 25360 7550
rect 25516 3058 25544 57151
rect 25504 3052 25556 3058
rect 25504 2994 25556 3000
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 68303
rect 27632 3602 27660 70994
rect 32402 61432 32458 61441
rect 32402 61367 32458 61376
rect 27710 50280 27766 50289
rect 27710 50215 27766 50224
rect 27620 3596 27672 3602
rect 27620 3538 27672 3544
rect 27724 480 27752 50215
rect 30378 48920 30434 48929
rect 30378 48855 30434 48864
rect 30392 16574 30420 48855
rect 31760 33788 31812 33794
rect 31760 33730 31812 33736
rect 31772 16574 31800 33730
rect 30392 16546 30880 16574
rect 31772 16546 31984 16574
rect 28540 3596 28592 3602
rect 28540 3538 28592 3544
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28552 354 28580 3538
rect 30104 3120 30156 3126
rect 30104 3062 30156 3068
rect 30116 480 30144 3062
rect 28878 354 28990 480
rect 28552 326 28990 354
rect 28878 -960 28990 326
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31956 354 31984 16546
rect 32416 3126 32444 61367
rect 33600 3188 33652 3194
rect 33600 3130 33652 3136
rect 32404 3120 32456 3126
rect 32404 3062 32456 3068
rect 33612 480 33640 3130
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 31270 -960 31382 326
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34532 354 34560 76463
rect 35900 75200 35952 75206
rect 35900 75142 35952 75148
rect 35164 71120 35216 71126
rect 35164 71062 35216 71068
rect 35176 3194 35204 71062
rect 35912 6914 35940 75142
rect 40038 66872 40094 66881
rect 40038 66807 40094 66816
rect 35992 65612 36044 65618
rect 35992 65554 36044 65560
rect 36004 16574 36032 65554
rect 38658 64152 38714 64161
rect 38658 64087 38714 64096
rect 38672 16574 38700 64087
rect 39302 47560 39358 47569
rect 39302 47495 39358 47504
rect 36004 16546 36768 16574
rect 38672 16546 39160 16574
rect 35912 6886 36032 6914
rect 35164 3188 35216 3194
rect 35164 3130 35216 3136
rect 36004 480 36032 6886
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36740 354 36768 16546
rect 38384 3188 38436 3194
rect 38384 3130 38436 3136
rect 38396 480 38424 3130
rect 37158 354 37270 480
rect 36740 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39132 354 39160 16546
rect 39316 3194 39344 47495
rect 40052 16574 40080 66807
rect 40696 59362 40724 142258
rect 60740 78328 60792 78334
rect 60740 78270 60792 78276
rect 57980 78124 58032 78130
rect 57980 78066 58032 78072
rect 53840 78056 53892 78062
rect 53840 77998 53892 78004
rect 46940 77988 46992 77994
rect 46940 77930 46992 77936
rect 45560 69692 45612 69698
rect 45560 69634 45612 69640
rect 43444 61396 43496 61402
rect 43444 61338 43496 61344
rect 40684 59356 40736 59362
rect 40684 59298 40736 59304
rect 42800 31068 42852 31074
rect 42800 31010 42852 31016
rect 40052 16546 40264 16574
rect 39304 3188 39356 3194
rect 39304 3130 39356 3136
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 40236 354 40264 16546
rect 41880 3188 41932 3194
rect 41880 3130 41932 3136
rect 41892 480 41920 3130
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 39550 -960 39662 326
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 42812 354 42840 31010
rect 43456 3194 43484 61338
rect 44180 60104 44232 60110
rect 44180 60046 44232 60052
rect 44192 6914 44220 60046
rect 44270 46200 44326 46209
rect 44270 46135 44326 46144
rect 44284 16574 44312 46135
rect 45572 16574 45600 69634
rect 46952 16574 46980 77930
rect 52460 72616 52512 72622
rect 52460 72558 52512 72564
rect 48320 68332 48372 68338
rect 48320 68274 48372 68280
rect 48332 16574 48360 68274
rect 49698 58576 49754 58585
rect 49698 58511 49754 58520
rect 49712 16574 49740 58511
rect 52472 16574 52500 72558
rect 53852 16574 53880 77998
rect 54482 73944 54538 73953
rect 54482 73879 54538 73888
rect 44284 16546 45048 16574
rect 45572 16546 46704 16574
rect 46952 16546 47440 16574
rect 48332 16546 48544 16574
rect 49712 16546 50200 16574
rect 52472 16546 53328 16574
rect 53852 16546 54432 16574
rect 44192 6886 44312 6914
rect 43444 3188 43496 3194
rect 43444 3130 43496 3136
rect 44284 480 44312 6886
rect 43046 354 43158 480
rect 42812 326 43158 354
rect 43046 -960 43158 326
rect 44242 -960 44354 480
rect 45020 354 45048 16546
rect 46676 480 46704 16546
rect 45438 354 45550 480
rect 45020 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 48516 354 48544 16546
rect 50172 480 50200 16546
rect 52552 8968 52604 8974
rect 52552 8910 52604 8916
rect 51356 3596 51408 3602
rect 51356 3538 51408 3544
rect 51368 480 51396 3538
rect 52564 480 52592 8910
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 47830 -960 47942 326
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53300 354 53328 16546
rect 54404 3482 54432 16546
rect 54496 3602 54524 73879
rect 57242 64288 57298 64297
rect 57242 64223 57298 64232
rect 56598 53136 56654 53145
rect 56598 53071 56654 53080
rect 56612 16574 56640 53071
rect 56612 16546 56824 16574
rect 54484 3596 54536 3602
rect 54484 3538 54536 3544
rect 56048 3596 56100 3602
rect 56048 3538 56100 3544
rect 54404 3454 54984 3482
rect 54956 480 54984 3454
rect 56060 480 56088 3538
rect 53718 354 53830 480
rect 53300 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 57256 3602 57284 64223
rect 57992 16574 58020 78066
rect 59360 76560 59412 76566
rect 59360 76502 59412 76508
rect 57992 16546 58480 16574
rect 57244 3596 57296 3602
rect 57244 3538 57296 3544
rect 58452 480 58480 16546
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59372 354 59400 76502
rect 60752 3602 60780 78270
rect 75920 78260 75972 78266
rect 75920 78202 75972 78208
rect 67638 76664 67694 76673
rect 66260 76628 66312 76634
rect 67638 76599 67694 76608
rect 66260 76570 66312 76576
rect 60832 69760 60884 69766
rect 60832 69702 60884 69708
rect 60740 3596 60792 3602
rect 60740 3538 60792 3544
rect 60844 480 60872 69702
rect 62120 64184 62172 64190
rect 62120 64126 62172 64132
rect 62132 16574 62160 64126
rect 63498 43480 63554 43489
rect 63498 43415 63554 43424
rect 63512 16574 63540 43415
rect 66272 16574 66300 76570
rect 62132 16546 63264 16574
rect 63512 16546 64368 16574
rect 66272 16546 66760 16574
rect 61660 3596 61712 3602
rect 61660 3538 61712 3544
rect 59606 354 59718 480
rect 59372 326 59718 354
rect 59606 -960 59718 326
rect 60802 -960 60914 480
rect 61672 354 61700 3538
rect 63236 480 63264 16546
rect 64340 480 64368 16546
rect 65524 3664 65576 3670
rect 65524 3606 65576 3612
rect 65536 480 65564 3606
rect 66732 480 66760 16546
rect 61998 354 62110 480
rect 61672 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67652 354 67680 76599
rect 71044 75268 71096 75274
rect 71044 75210 71096 75216
rect 69020 58676 69072 58682
rect 69020 58618 69072 58624
rect 69032 16574 69060 58618
rect 70400 42084 70452 42090
rect 70400 42026 70452 42032
rect 70412 16574 70440 42026
rect 69032 16546 69888 16574
rect 70412 16546 70992 16574
rect 69112 3596 69164 3602
rect 69112 3538 69164 3544
rect 69124 480 69152 3538
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 69860 354 69888 16546
rect 70964 3482 70992 16546
rect 71056 3602 71084 75210
rect 71780 71188 71832 71194
rect 71780 71130 71832 71136
rect 71792 16574 71820 71130
rect 75182 62928 75238 62937
rect 75182 62863 75238 62872
rect 74540 40724 74592 40730
rect 74540 40666 74592 40672
rect 74552 16574 74580 40666
rect 71792 16546 72648 16574
rect 74552 16546 75040 16574
rect 71044 3596 71096 3602
rect 71044 3538 71096 3544
rect 70964 3454 71544 3482
rect 71516 480 71544 3454
rect 72620 480 72648 16546
rect 73804 4140 73856 4146
rect 73804 4082 73856 4088
rect 73816 480 73844 4082
rect 75012 480 75040 16546
rect 75196 4146 75224 62863
rect 75184 4140 75236 4146
rect 75184 4082 75236 4088
rect 70278 354 70390 480
rect 69860 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 75932 354 75960 78202
rect 93860 75540 93912 75546
rect 93860 75482 93912 75488
rect 85580 75404 85632 75410
rect 85580 75346 85632 75352
rect 84198 67008 84254 67017
rect 84198 66943 84254 66952
rect 80060 66904 80112 66910
rect 80060 66846 80112 66852
rect 77298 57352 77354 57361
rect 77298 57287 77354 57296
rect 77312 6914 77340 57287
rect 78678 50416 78734 50425
rect 78678 50351 78734 50360
rect 77392 39364 77444 39370
rect 77392 39306 77444 39312
rect 77404 16574 77432 39306
rect 78692 16574 78720 50351
rect 80072 16574 80100 66846
rect 81438 63064 81494 63073
rect 81438 62999 81494 63008
rect 81452 16574 81480 62999
rect 77404 16546 78168 16574
rect 78692 16546 79272 16574
rect 80072 16546 80928 16574
rect 81452 16546 81664 16574
rect 77312 6886 77432 6914
rect 77404 480 77432 6886
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78140 354 78168 16546
rect 78558 354 78670 480
rect 78140 326 78670 354
rect 79244 354 79272 16546
rect 80900 480 80928 16546
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 78558 -960 78670 326
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 83280 3664 83332 3670
rect 83280 3606 83332 3612
rect 83292 480 83320 3606
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84212 354 84240 66943
rect 85592 6914 85620 75346
rect 89720 73908 89772 73914
rect 89720 73850 89772 73856
rect 85672 69828 85724 69834
rect 85672 69770 85724 69776
rect 85684 16574 85712 69770
rect 88338 55992 88394 56001
rect 88338 55927 88394 55936
rect 88352 16574 88380 55927
rect 89732 16574 89760 73850
rect 93122 65512 93178 65521
rect 93122 65447 93178 65456
rect 92478 54496 92534 54505
rect 92478 54431 92534 54440
rect 85684 16546 86448 16574
rect 88352 16546 89208 16574
rect 89732 16546 89944 16574
rect 85592 6886 85712 6914
rect 85684 480 85712 6886
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86420 354 86448 16546
rect 87512 15904 87564 15910
rect 87512 15846 87564 15852
rect 86838 354 86950 480
rect 86420 326 86950 354
rect 87524 354 87552 15846
rect 89180 480 89208 16546
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 86838 -960 86950 326
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91560 3392 91612 3398
rect 91560 3334 91612 3340
rect 91572 480 91600 3334
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 54431
rect 93136 3398 93164 65447
rect 93872 6914 93900 75482
rect 96620 72684 96672 72690
rect 96620 72626 96672 72632
rect 93950 61568 94006 61577
rect 93950 61503 94006 61512
rect 93964 16574 93992 61503
rect 95240 36576 95292 36582
rect 95240 36518 95292 36524
rect 95252 16574 95280 36518
rect 96632 16574 96660 72626
rect 97276 33114 97304 153206
rect 97356 140888 97408 140894
rect 97356 140830 97408 140836
rect 97368 85542 97396 140830
rect 97356 85536 97408 85542
rect 97356 85478 97408 85484
rect 97920 75138 97948 196590
rect 100298 195392 100354 195401
rect 100298 195327 100354 195336
rect 99196 191276 99248 191282
rect 99196 191218 99248 191224
rect 99104 187196 99156 187202
rect 99104 187138 99156 187144
rect 99012 187060 99064 187066
rect 99012 187002 99064 187008
rect 98920 154080 98972 154086
rect 98920 154022 98972 154028
rect 98828 148368 98880 148374
rect 98828 148310 98880 148316
rect 97908 75132 97960 75138
rect 97908 75074 97960 75080
rect 98840 72554 98868 148310
rect 98828 72548 98880 72554
rect 98828 72490 98880 72496
rect 98840 72350 98868 72490
rect 98828 72344 98880 72350
rect 98828 72286 98880 72292
rect 98932 60722 98960 154022
rect 99024 75342 99052 187002
rect 99012 75336 99064 75342
rect 99012 75278 99064 75284
rect 99116 72554 99144 187138
rect 99104 72548 99156 72554
rect 99104 72490 99156 72496
rect 99208 72486 99236 191218
rect 99288 187128 99340 187134
rect 99288 187070 99340 187076
rect 99196 72480 99248 72486
rect 99196 72422 99248 72428
rect 99208 72282 99236 72422
rect 99196 72276 99248 72282
rect 99196 72218 99248 72224
rect 99300 67590 99328 187070
rect 100208 186992 100260 186998
rect 100208 186934 100260 186940
rect 100024 154012 100076 154018
rect 100024 153954 100076 153960
rect 99932 153876 99984 153882
rect 99932 153818 99984 153824
rect 99840 151292 99892 151298
rect 99840 151234 99892 151240
rect 99852 77790 99880 151234
rect 99840 77784 99892 77790
rect 99840 77726 99892 77732
rect 99380 76696 99432 76702
rect 99380 76638 99432 76644
rect 99288 67584 99340 67590
rect 99288 67526 99340 67532
rect 98920 60716 98972 60722
rect 98920 60658 98972 60664
rect 98932 60042 98960 60658
rect 98920 60036 98972 60042
rect 98920 59978 98972 59984
rect 97998 59936 98054 59945
rect 97998 59871 98054 59880
rect 97264 33108 97316 33114
rect 97264 33050 97316 33056
rect 98012 16574 98040 59871
rect 99392 16574 99420 76638
rect 99944 71058 99972 153818
rect 99932 71052 99984 71058
rect 99932 70994 99984 71000
rect 100036 66162 100064 153954
rect 100116 153944 100168 153950
rect 100116 153886 100168 153892
rect 100024 66156 100076 66162
rect 100024 66098 100076 66104
rect 100128 66094 100156 153886
rect 100220 78985 100248 186934
rect 100206 78976 100262 78985
rect 100206 78911 100262 78920
rect 100312 78606 100340 195327
rect 101678 194032 101734 194041
rect 101678 193967 101734 193976
rect 100484 192908 100536 192914
rect 100484 192850 100536 192856
rect 100392 191208 100444 191214
rect 100392 191150 100444 191156
rect 100300 78600 100352 78606
rect 100300 78542 100352 78548
rect 100404 74225 100432 191150
rect 100390 74216 100446 74225
rect 100390 74151 100446 74160
rect 100404 73817 100432 74151
rect 100390 73808 100446 73817
rect 100390 73743 100446 73752
rect 100116 66088 100168 66094
rect 100116 66030 100168 66036
rect 100496 65958 100524 192850
rect 100666 191312 100722 191321
rect 100666 191247 100722 191256
rect 100576 190188 100628 190194
rect 100576 190130 100628 190136
rect 99472 65952 99524 65958
rect 99472 65894 99524 65900
rect 100484 65952 100536 65958
rect 100484 65894 100536 65900
rect 99484 65550 99512 65894
rect 99472 65544 99524 65550
rect 99472 65486 99524 65492
rect 100588 52465 100616 190130
rect 99470 52456 99526 52465
rect 99470 52391 99526 52400
rect 100574 52456 100630 52465
rect 100574 52391 100630 52400
rect 99484 51785 99512 52391
rect 99470 51776 99526 51785
rect 99470 51711 99526 51720
rect 100680 49609 100708 191247
rect 101588 189780 101640 189786
rect 101588 189722 101640 189728
rect 101496 187264 101548 187270
rect 101496 187206 101548 187212
rect 101220 154148 101272 154154
rect 101220 154090 101272 154096
rect 100758 77072 100814 77081
rect 100758 77007 100814 77016
rect 100772 76537 100800 77007
rect 100758 76528 100814 76537
rect 100758 76463 100814 76472
rect 101232 75682 101260 154090
rect 101312 149728 101364 149734
rect 101312 149670 101364 149676
rect 101402 149696 101458 149705
rect 100760 75676 100812 75682
rect 100760 75618 100812 75624
rect 101220 75676 101272 75682
rect 101220 75618 101272 75624
rect 100772 75206 100800 75618
rect 100760 75200 100812 75206
rect 100760 75142 100812 75148
rect 101324 70378 101352 149670
rect 101402 149631 101458 149640
rect 100760 70372 100812 70378
rect 100760 70314 100812 70320
rect 101312 70372 101364 70378
rect 101312 70314 101364 70320
rect 100772 69698 100800 70314
rect 100760 69692 100812 69698
rect 100760 69634 100812 69640
rect 100760 68944 100812 68950
rect 100760 68886 100812 68892
rect 100772 68338 100800 68886
rect 100760 68332 100812 68338
rect 100760 68274 100812 68280
rect 100760 66224 100812 66230
rect 100760 66166 100812 66172
rect 100772 65618 100800 66166
rect 100760 65612 100812 65618
rect 100760 65554 100812 65560
rect 101416 64705 101444 149631
rect 101508 77081 101536 187206
rect 101494 77072 101550 77081
rect 101494 77007 101550 77016
rect 101600 68950 101628 189722
rect 101588 68944 101640 68950
rect 101588 68886 101640 68892
rect 101692 66230 101720 193967
rect 101862 191720 101918 191729
rect 101862 191655 101918 191664
rect 101770 191584 101826 191593
rect 101770 191519 101826 191528
rect 101680 66224 101732 66230
rect 101680 66166 101732 66172
rect 101402 64696 101458 64705
rect 101402 64631 101458 64640
rect 101416 64161 101444 64631
rect 101402 64152 101458 64161
rect 101402 64087 101458 64096
rect 101784 57769 101812 191519
rect 100758 57760 100814 57769
rect 100758 57695 100814 57704
rect 101770 57760 101826 57769
rect 101770 57695 101826 57704
rect 100772 57225 100800 57695
rect 100758 57216 100814 57225
rect 100758 57151 100814 57160
rect 101876 50289 101904 191655
rect 102046 191448 102102 191457
rect 102046 191383 102102 191392
rect 101954 191040 102010 191049
rect 101954 190975 102010 190984
rect 101862 50280 101918 50289
rect 101862 50215 101918 50224
rect 99470 49600 99526 49609
rect 99470 49535 99526 49544
rect 100666 49600 100722 49609
rect 100666 49535 100722 49544
rect 99484 48929 99512 49535
rect 99470 48920 99526 48929
rect 99470 48855 99526 48864
rect 101968 48249 101996 190975
rect 100758 48240 100814 48249
rect 100758 48175 100814 48184
rect 101954 48240 102010 48249
rect 101954 48175 102010 48184
rect 100772 47569 100800 48175
rect 100758 47560 100814 47569
rect 100758 47495 100814 47504
rect 102060 46889 102088 191383
rect 103060 191140 103112 191146
rect 103060 191082 103112 191088
rect 102876 189916 102928 189922
rect 102876 189858 102928 189864
rect 102600 151156 102652 151162
rect 102600 151098 102652 151104
rect 102140 77104 102192 77110
rect 102140 77046 102192 77052
rect 102152 76634 102180 77046
rect 102140 76628 102192 76634
rect 102140 76570 102192 76576
rect 102612 72962 102640 151098
rect 102782 151056 102838 151065
rect 102782 150991 102838 151000
rect 102692 149796 102744 149802
rect 102692 149738 102744 149744
rect 102600 72956 102652 72962
rect 102600 72898 102652 72904
rect 102140 68604 102192 68610
rect 102140 68546 102192 68552
rect 102152 68377 102180 68546
rect 102232 68468 102284 68474
rect 102232 68410 102284 68416
rect 102138 68368 102194 68377
rect 102138 68303 102194 68312
rect 102244 68241 102272 68410
rect 102230 68232 102286 68241
rect 102230 68167 102286 68176
rect 102704 66026 102732 149738
rect 102692 66020 102744 66026
rect 102692 65962 102744 65968
rect 102690 62112 102746 62121
rect 102232 62076 102284 62082
rect 102690 62047 102746 62056
rect 102232 62018 102284 62024
rect 102140 62008 102192 62014
rect 102140 61950 102192 61956
rect 102152 61441 102180 61950
rect 102138 61432 102194 61441
rect 102244 61402 102272 62018
rect 102704 62014 102732 62047
rect 102692 62008 102744 62014
rect 102692 61950 102744 61956
rect 102138 61367 102194 61376
rect 102232 61396 102284 61402
rect 102232 61338 102284 61344
rect 102140 60648 102192 60654
rect 102140 60590 102192 60596
rect 102152 60110 102180 60590
rect 102140 60104 102192 60110
rect 102140 60046 102192 60052
rect 102138 54632 102194 54641
rect 102138 54567 102194 54576
rect 100758 46880 100814 46889
rect 100758 46815 100814 46824
rect 102046 46880 102102 46889
rect 102046 46815 102102 46824
rect 100772 46209 100800 46815
rect 100758 46200 100814 46209
rect 100758 46135 100814 46144
rect 102152 16574 102180 54567
rect 102796 44169 102824 150991
rect 102888 77110 102916 189858
rect 102968 189848 103020 189854
rect 102968 189790 103020 189796
rect 102876 77104 102928 77110
rect 102876 77046 102928 77052
rect 102980 76566 103008 189790
rect 102968 76560 103020 76566
rect 102968 76502 103020 76508
rect 103072 75886 103100 191082
rect 103164 78577 103192 198018
rect 104440 195492 104492 195498
rect 104440 195434 104492 195440
rect 103242 194304 103298 194313
rect 103242 194239 103298 194248
rect 103150 78568 103206 78577
rect 103150 78503 103206 78512
rect 103060 75880 103112 75886
rect 103060 75822 103112 75828
rect 103256 71126 103284 194239
rect 104348 192568 104400 192574
rect 104348 192510 104400 192516
rect 103336 191344 103388 191350
rect 103336 191286 103388 191292
rect 103244 71120 103296 71126
rect 103244 71062 103296 71068
rect 102876 69692 102928 69698
rect 102876 69634 102928 69640
rect 102230 44160 102286 44169
rect 102230 44095 102286 44104
rect 102782 44160 102838 44169
rect 102782 44095 102838 44104
rect 102244 43489 102272 44095
rect 102230 43480 102286 43489
rect 102230 43415 102286 43424
rect 93964 16546 94728 16574
rect 95252 16546 95832 16574
rect 96632 16546 97488 16574
rect 98012 16546 98224 16574
rect 99392 16546 99880 16574
rect 102152 16546 102272 16574
rect 93872 6886 93992 6914
rect 93124 3392 93176 3398
rect 93124 3334 93176 3340
rect 93964 480 93992 6886
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 94700 354 94728 16546
rect 95118 354 95230 480
rect 94700 326 95230 354
rect 95804 354 95832 16546
rect 97460 480 97488 16546
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 95118 -960 95230 326
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98196 354 98224 16546
rect 99852 480 99880 16546
rect 101036 3392 101088 3398
rect 101036 3334 101088 3340
rect 101048 480 101076 3334
rect 102244 480 102272 16546
rect 102888 3398 102916 69634
rect 103058 68912 103114 68921
rect 103058 68847 103114 68856
rect 103072 68610 103100 68847
rect 103060 68604 103112 68610
rect 103060 68546 103112 68552
rect 103348 62082 103376 191286
rect 104256 190256 104308 190262
rect 104256 190198 104308 190204
rect 103428 190120 103480 190126
rect 103428 190062 103480 190068
rect 103336 62076 103388 62082
rect 103336 62018 103388 62024
rect 103440 60654 103468 190062
rect 104164 151360 104216 151366
rect 104164 151302 104216 151308
rect 104072 151088 104124 151094
rect 104072 151030 104124 151036
rect 103980 144356 104032 144362
rect 103980 144298 104032 144304
rect 103992 81977 104020 144298
rect 103978 81968 104034 81977
rect 103978 81903 104034 81912
rect 104084 75818 104112 151030
rect 103888 75812 103940 75818
rect 103888 75754 103940 75760
rect 104072 75812 104124 75818
rect 104072 75754 104124 75760
rect 103900 75410 103928 75754
rect 103888 75404 103940 75410
rect 103888 75346 103940 75352
rect 103520 70440 103572 70446
rect 103520 70382 103572 70388
rect 103428 60648 103480 60654
rect 103428 60590 103480 60596
rect 103532 16574 103560 70382
rect 104176 70242 104204 151302
rect 104268 75478 104296 190198
rect 104256 75472 104308 75478
rect 104256 75414 104308 75420
rect 104360 73778 104388 192510
rect 104452 75614 104480 195434
rect 104532 195424 104584 195430
rect 104532 195366 104584 195372
rect 104440 75608 104492 75614
rect 104440 75550 104492 75556
rect 104452 75274 104480 75550
rect 104440 75268 104492 75274
rect 104440 75210 104492 75216
rect 104348 73772 104400 73778
rect 104348 73714 104400 73720
rect 104544 71602 104572 195366
rect 104624 189984 104676 189990
rect 104624 189926 104676 189932
rect 104532 71596 104584 71602
rect 104532 71538 104584 71544
rect 104544 71194 104572 71538
rect 104532 71188 104584 71194
rect 104532 71130 104584 71136
rect 104164 70236 104216 70242
rect 104164 70178 104216 70184
rect 104176 69766 104204 70178
rect 104164 69760 104216 69766
rect 104164 69702 104216 69708
rect 104532 67312 104584 67318
rect 104532 67254 104584 67260
rect 104544 66881 104572 67254
rect 104530 66872 104586 66881
rect 104530 66807 104586 66816
rect 104256 64864 104308 64870
rect 104256 64806 104308 64812
rect 104268 64705 104296 64806
rect 104636 64802 104664 189926
rect 104714 189680 104770 189689
rect 104714 189615 104770 189624
rect 104624 64796 104676 64802
rect 104624 64738 104676 64744
rect 104254 64696 104310 64705
rect 104254 64631 104310 64640
rect 104268 64297 104296 64631
rect 104254 64288 104310 64297
rect 104254 64223 104310 64232
rect 104636 64190 104664 64738
rect 104624 64184 104676 64190
rect 104624 64126 104676 64132
rect 104162 59256 104218 59265
rect 104162 59191 104164 59200
rect 104216 59191 104218 59200
rect 104164 59162 104216 59168
rect 104176 58585 104204 59162
rect 104162 58576 104218 58585
rect 104162 58511 104218 58520
rect 104728 57905 104756 189615
rect 103794 57896 103850 57905
rect 103794 57831 103850 57840
rect 104714 57896 104770 57905
rect 104714 57831 104770 57840
rect 103808 57361 103836 57831
rect 103794 57352 103850 57361
rect 103794 57287 103850 57296
rect 104820 50969 104848 200466
rect 107198 199200 107254 199209
rect 107198 199135 107254 199144
rect 105728 198280 105780 198286
rect 105728 198222 105780 198228
rect 105910 198248 105966 198257
rect 105636 197328 105688 197334
rect 105636 197270 105688 197276
rect 105544 196716 105596 196722
rect 105544 196658 105596 196664
rect 105450 151328 105506 151337
rect 105450 151263 105506 151272
rect 105358 151192 105414 151201
rect 105358 151127 105414 151136
rect 105268 80572 105320 80578
rect 105268 80514 105320 80520
rect 105280 78538 105308 80514
rect 105268 78532 105320 78538
rect 105268 78474 105320 78480
rect 105280 75546 105308 78474
rect 105268 75540 105320 75546
rect 105268 75482 105320 75488
rect 105372 63481 105400 151127
rect 105358 63472 105414 63481
rect 105358 63407 105414 63416
rect 105464 53825 105492 151263
rect 105556 78470 105584 196658
rect 105648 80578 105676 197270
rect 105636 80572 105688 80578
rect 105636 80514 105688 80520
rect 105740 80458 105768 198222
rect 105910 198183 105966 198192
rect 107016 198212 107068 198218
rect 105820 193044 105872 193050
rect 105820 192986 105872 192992
rect 105648 80430 105768 80458
rect 105544 78464 105596 78470
rect 105544 78406 105596 78412
rect 105648 78033 105676 80430
rect 105728 78464 105780 78470
rect 105728 78406 105780 78412
rect 105740 78266 105768 78406
rect 105728 78260 105780 78266
rect 105728 78202 105780 78208
rect 105634 78024 105690 78033
rect 105634 77959 105690 77968
rect 105832 71670 105860 192986
rect 105924 73710 105952 198183
rect 107016 198154 107068 198160
rect 106922 196888 106978 196897
rect 106922 196823 106978 196832
rect 106002 194168 106058 194177
rect 106002 194103 106058 194112
rect 105912 73704 105964 73710
rect 105912 73646 105964 73652
rect 105820 71664 105872 71670
rect 105820 71606 105872 71612
rect 105832 70446 105860 71606
rect 105820 70440 105872 70446
rect 105820 70382 105872 70388
rect 106016 70174 106044 194103
rect 106094 191176 106150 191185
rect 106094 191111 106150 191120
rect 106004 70168 106056 70174
rect 106004 70110 106056 70116
rect 106108 62121 106136 191111
rect 106188 190324 106240 190330
rect 106188 190266 106240 190272
rect 106094 62112 106150 62121
rect 106094 62047 106150 62056
rect 106200 59158 106228 190266
rect 106832 151496 106884 151502
rect 106832 151438 106884 151444
rect 106740 151224 106792 151230
rect 106740 151166 106792 151172
rect 106752 74390 106780 151166
rect 106740 74384 106792 74390
rect 106740 74326 106792 74332
rect 106752 73234 106780 74326
rect 106280 73228 106332 73234
rect 106280 73170 106332 73176
rect 106740 73228 106792 73234
rect 106740 73170 106792 73176
rect 106004 59152 106056 59158
rect 106004 59094 106056 59100
rect 106188 59152 106240 59158
rect 106188 59094 106240 59100
rect 106016 58682 106044 59094
rect 106004 58676 106056 58682
rect 106004 58618 106056 58624
rect 105450 53816 105506 53825
rect 105450 53751 105506 53760
rect 105464 53145 105492 53751
rect 105450 53136 105506 53145
rect 105450 53071 105506 53080
rect 104806 50960 104862 50969
rect 104806 50895 104862 50904
rect 106292 16574 106320 73170
rect 106844 68678 106872 151438
rect 106936 78062 106964 196823
rect 106924 78056 106976 78062
rect 106924 77998 106976 78004
rect 107028 77994 107056 198154
rect 107108 193112 107160 193118
rect 107108 193054 107160 193060
rect 107016 77988 107068 77994
rect 107016 77930 107068 77936
rect 107120 72894 107148 193054
rect 107212 78402 107240 199135
rect 107200 78396 107252 78402
rect 107200 78338 107252 78344
rect 107304 78130 107332 200534
rect 110236 200252 110288 200258
rect 110236 200194 110288 200200
rect 109868 199640 109920 199646
rect 109868 199582 109920 199588
rect 108580 199096 108632 199102
rect 108580 199038 108632 199044
rect 108396 197872 108448 197878
rect 108396 197814 108448 197820
rect 108304 197192 108356 197198
rect 108304 197134 108356 197140
rect 108210 195528 108266 195537
rect 108210 195463 108266 195472
rect 107384 190392 107436 190398
rect 107384 190334 107436 190340
rect 107292 78124 107344 78130
rect 107292 78066 107344 78072
rect 107396 74534 107424 190334
rect 107474 190088 107530 190097
rect 107474 190023 107530 190032
rect 107304 74506 107424 74534
rect 107198 74080 107254 74089
rect 107198 74015 107254 74024
rect 107212 73846 107240 74015
rect 107200 73840 107252 73846
rect 107200 73782 107252 73788
rect 107108 72888 107160 72894
rect 107108 72830 107160 72836
rect 107120 72690 107148 72830
rect 107108 72684 107160 72690
rect 107108 72626 107160 72632
rect 106832 68672 106884 68678
rect 106832 68614 106884 68620
rect 107304 67250 107332 74506
rect 107382 71088 107438 71097
rect 107382 71023 107384 71032
rect 107436 71023 107438 71032
rect 107384 70994 107436 71000
rect 107292 67244 107344 67250
rect 107292 67186 107344 67192
rect 106922 66192 106978 66201
rect 106922 66127 106978 66136
rect 103532 16546 104112 16574
rect 106292 16546 106504 16574
rect 103336 6180 103388 6186
rect 103336 6122 103388 6128
rect 102876 3392 102928 3398
rect 102876 3334 102928 3340
rect 103348 480 103376 6122
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16546
rect 105728 3392 105780 3398
rect 105728 3334 105780 3340
rect 105740 480 105768 3334
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 106936 3398 106964 66127
rect 107488 63209 107516 190023
rect 107566 186960 107622 186969
rect 107566 186895 107622 186904
rect 107474 63200 107530 63209
rect 107474 63135 107530 63144
rect 107580 55185 107608 186895
rect 108118 137864 108174 137873
rect 108118 137799 108174 137808
rect 108132 77858 108160 137799
rect 108224 79422 108252 195463
rect 108212 79416 108264 79422
rect 108212 79358 108264 79364
rect 108316 78062 108344 197134
rect 108304 78056 108356 78062
rect 108304 77998 108356 78004
rect 108408 77994 108436 197814
rect 108488 194132 108540 194138
rect 108488 194074 108540 194080
rect 108396 77988 108448 77994
rect 108396 77930 108448 77936
rect 108120 77852 108172 77858
rect 108120 77794 108172 77800
rect 108500 74186 108528 194074
rect 108592 75070 108620 199038
rect 108948 198144 109000 198150
rect 108948 198086 109000 198092
rect 108856 195288 108908 195294
rect 108856 195230 108908 195236
rect 108672 194064 108724 194070
rect 108672 194006 108724 194012
rect 108580 75064 108632 75070
rect 108580 75006 108632 75012
rect 108488 74180 108540 74186
rect 108488 74122 108540 74128
rect 108500 73234 108528 74122
rect 107660 73228 107712 73234
rect 107660 73170 107712 73176
rect 108488 73228 108540 73234
rect 108488 73170 108540 73176
rect 107566 55176 107622 55185
rect 107566 55111 107622 55120
rect 107580 54641 107608 55111
rect 107566 54632 107622 54641
rect 107566 54567 107622 54576
rect 107672 16574 107700 73170
rect 108684 70106 108712 194006
rect 108764 192636 108816 192642
rect 108764 192578 108816 192584
rect 108396 70100 108448 70106
rect 108396 70042 108448 70048
rect 108672 70100 108724 70106
rect 108672 70042 108724 70048
rect 108408 69698 108436 70042
rect 108396 69692 108448 69698
rect 108396 69634 108448 69640
rect 108776 68882 108804 192578
rect 108764 68876 108816 68882
rect 108764 68818 108816 68824
rect 108868 67522 108896 195230
rect 108960 68814 108988 198086
rect 109592 151428 109644 151434
rect 109592 151370 109644 151376
rect 109500 146940 109552 146946
rect 109500 146882 109552 146888
rect 109512 77926 109540 146882
rect 109500 77920 109552 77926
rect 109500 77862 109552 77868
rect 109512 77314 109540 77862
rect 109040 77308 109092 77314
rect 109040 77250 109092 77256
rect 109500 77308 109552 77314
rect 109500 77250 109552 77256
rect 108948 68808 109000 68814
rect 108948 68750 109000 68756
rect 108856 67516 108908 67522
rect 108856 67458 108908 67464
rect 108304 67176 108356 67182
rect 108304 67118 108356 67124
rect 108316 67017 108344 67118
rect 108302 67008 108358 67017
rect 108302 66943 108358 66952
rect 108946 66192 109002 66201
rect 108946 66127 109002 66136
rect 108960 65822 108988 66127
rect 108948 65816 109000 65822
rect 108948 65758 109000 65764
rect 107672 16546 108160 16574
rect 106924 3392 106976 3398
rect 106924 3334 106976 3340
rect 108132 480 108160 16546
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109052 354 109080 77250
rect 109604 76945 109632 151370
rect 109684 147280 109736 147286
rect 109684 147222 109736 147228
rect 109590 76936 109646 76945
rect 109590 76871 109646 76880
rect 109604 64874 109632 76871
rect 109696 72486 109724 147222
rect 109776 147008 109828 147014
rect 109776 146950 109828 146956
rect 109684 72480 109736 72486
rect 109684 72422 109736 72428
rect 109788 72418 109816 146950
rect 109880 79626 109908 199582
rect 109960 195356 110012 195362
rect 109960 195298 110012 195304
rect 109868 79620 109920 79626
rect 109868 79562 109920 79568
rect 109972 74254 110000 195298
rect 110144 192772 110196 192778
rect 110144 192714 110196 192720
rect 110052 192500 110104 192506
rect 110052 192442 110104 192448
rect 109960 74248 110012 74254
rect 109960 74190 110012 74196
rect 109776 72412 109828 72418
rect 109776 72354 109828 72360
rect 110064 69018 110092 192442
rect 110052 69012 110104 69018
rect 110052 68954 110104 68960
rect 110156 67561 110184 192714
rect 110248 72826 110276 200194
rect 110328 192840 110380 192846
rect 110328 192782 110380 192788
rect 110236 72820 110288 72826
rect 110236 72762 110288 72768
rect 110142 67552 110198 67561
rect 110142 67487 110198 67496
rect 109604 64846 109908 64874
rect 109880 59362 109908 64846
rect 110340 64705 110368 192782
rect 110788 147076 110840 147082
rect 110788 147018 110840 147024
rect 110800 68338 110828 147018
rect 110970 146976 111026 146985
rect 110970 146911 111026 146920
rect 110878 139088 110934 139097
rect 110878 139023 110934 139032
rect 110892 76702 110920 139023
rect 110880 76696 110932 76702
rect 110880 76638 110932 76644
rect 110984 76430 111012 146911
rect 111076 145926 111104 260986
rect 112444 260024 112496 260030
rect 112444 259966 112496 259972
rect 111708 199708 111760 199714
rect 111708 199650 111760 199656
rect 111524 196988 111576 196994
rect 111524 196930 111576 196936
rect 111156 196784 111208 196790
rect 111156 196726 111208 196732
rect 111064 145920 111116 145926
rect 111064 145862 111116 145868
rect 111168 79490 111196 196726
rect 111340 195628 111392 195634
rect 111340 195570 111392 195576
rect 111248 193860 111300 193866
rect 111248 193802 111300 193808
rect 111156 79484 111208 79490
rect 111156 79426 111208 79432
rect 111260 77246 111288 193802
rect 111248 77240 111300 77246
rect 111248 77182 111300 77188
rect 110972 76424 111024 76430
rect 110972 76366 111024 76372
rect 111352 73982 111380 195570
rect 111432 193928 111484 193934
rect 111432 193870 111484 193876
rect 111340 73976 111392 73982
rect 111340 73918 111392 73924
rect 111444 73137 111472 193870
rect 111430 73128 111486 73137
rect 111430 73063 111486 73072
rect 111536 72690 111564 196930
rect 111616 190052 111668 190058
rect 111616 189994 111668 190000
rect 111524 72684 111576 72690
rect 111524 72626 111576 72632
rect 110788 68332 110840 68338
rect 110788 68274 110840 68280
rect 110326 64696 110382 64705
rect 110326 64631 110382 64640
rect 111628 64569 111656 189994
rect 111720 76786 111748 199650
rect 112456 154426 112484 259966
rect 112444 154420 112496 154426
rect 112444 154362 112496 154368
rect 111984 151564 112036 151570
rect 111984 151506 112036 151512
rect 111892 147348 111944 147354
rect 111892 147290 111944 147296
rect 111720 76758 111840 76786
rect 111706 76664 111762 76673
rect 111706 76599 111762 76608
rect 111720 76498 111748 76599
rect 111708 76492 111760 76498
rect 111708 76434 111760 76440
rect 111812 76378 111840 76758
rect 111720 76350 111840 76378
rect 111720 71058 111748 76350
rect 111904 75750 111932 147290
rect 111892 75744 111944 75750
rect 111892 75686 111944 75692
rect 111708 71052 111760 71058
rect 111708 70994 111760 71000
rect 111996 69970 112024 151506
rect 112168 149864 112220 149870
rect 112168 149806 112220 149812
rect 112076 148708 112128 148714
rect 112076 148650 112128 148656
rect 112088 71262 112116 148650
rect 112076 71256 112128 71262
rect 112076 71198 112128 71204
rect 111984 69964 112036 69970
rect 111984 69906 112036 69912
rect 112180 65550 112208 149806
rect 112548 148442 112576 262239
rect 112628 260908 112680 260914
rect 112628 260850 112680 260856
rect 112536 148436 112588 148442
rect 112536 148378 112588 148384
rect 112444 144832 112496 144838
rect 112444 144774 112496 144780
rect 112352 144084 112404 144090
rect 112352 144026 112404 144032
rect 112260 140208 112312 140214
rect 112260 140150 112312 140156
rect 112272 80782 112300 140150
rect 112364 81122 112392 144026
rect 112352 81116 112404 81122
rect 112352 81058 112404 81064
rect 112260 80776 112312 80782
rect 112260 80718 112312 80724
rect 112456 78878 112484 144774
rect 112640 144294 112668 260850
rect 112720 196920 112772 196926
rect 112720 196862 112772 196868
rect 112628 144288 112680 144294
rect 112628 144230 112680 144236
rect 112534 138680 112590 138689
rect 112534 138615 112590 138624
rect 112444 78872 112496 78878
rect 112444 78814 112496 78820
rect 112442 75304 112498 75313
rect 112442 75239 112498 75248
rect 112456 75206 112484 75239
rect 112444 75200 112496 75206
rect 112444 75142 112496 75148
rect 112168 65544 112220 65550
rect 112168 65486 112220 65492
rect 111614 64560 111670 64569
rect 111614 64495 111670 64504
rect 112258 60616 112314 60625
rect 111800 60580 111852 60586
rect 112258 60551 112260 60560
rect 111800 60522 111852 60528
rect 112312 60551 112314 60560
rect 112260 60522 112312 60528
rect 111812 59945 111840 60522
rect 111798 59936 111854 59945
rect 111798 59871 111854 59880
rect 109868 59356 109920 59362
rect 109868 59298 109920 59304
rect 110420 59356 110472 59362
rect 110420 59298 110472 59304
rect 110432 16574 110460 59298
rect 110432 16546 110552 16574
rect 110524 480 110552 16546
rect 112456 3398 112484 75142
rect 112548 68746 112576 138615
rect 112732 79014 112760 196862
rect 112824 145654 112852 264998
rect 112904 261180 112956 261186
rect 112904 261122 112956 261128
rect 112812 145648 112864 145654
rect 112812 145590 112864 145596
rect 112916 141846 112944 261122
rect 112996 197056 113048 197062
rect 112996 196998 113048 197004
rect 112904 141840 112956 141846
rect 112904 141782 112956 141788
rect 112720 79008 112772 79014
rect 112720 78950 112772 78956
rect 113008 76838 113036 196998
rect 113100 141642 113128 265134
rect 116584 265124 116636 265130
rect 116584 265066 116636 265072
rect 115388 262880 115440 262886
rect 115388 262822 115440 262828
rect 114008 262608 114060 262614
rect 114008 262550 114060 262556
rect 113732 260160 113784 260166
rect 113732 260102 113784 260108
rect 113744 154290 113772 260102
rect 113824 259684 113876 259690
rect 113824 259626 113876 259632
rect 113732 154284 113784 154290
rect 113732 154226 113784 154232
rect 113548 151632 113600 151638
rect 113548 151574 113600 151580
rect 113088 141636 113140 141642
rect 113088 141578 113140 141584
rect 112996 76832 113048 76838
rect 112996 76774 113048 76780
rect 113180 70440 113232 70446
rect 113180 70382 113232 70388
rect 112536 68740 112588 68746
rect 112536 68682 112588 68688
rect 113192 16574 113220 70382
rect 113560 69902 113588 151574
rect 113836 148986 113864 259626
rect 113916 193996 113968 194002
rect 113916 193938 113968 193944
rect 113824 148980 113876 148986
rect 113824 148922 113876 148928
rect 113732 147416 113784 147422
rect 113732 147358 113784 147364
rect 113640 144152 113692 144158
rect 113640 144094 113692 144100
rect 113652 80714 113680 144094
rect 113640 80708 113692 80714
rect 113640 80650 113692 80656
rect 113744 79694 113772 147358
rect 113824 147144 113876 147150
rect 113824 147086 113876 147092
rect 113732 79688 113784 79694
rect 113732 79630 113784 79636
rect 113836 76634 113864 147086
rect 113928 80850 113956 193938
rect 114020 145994 114048 262550
rect 115110 262440 115166 262449
rect 115110 262375 115166 262384
rect 114192 260296 114244 260302
rect 114192 260238 114244 260244
rect 114100 259548 114152 259554
rect 114100 259490 114152 259496
rect 114008 145988 114060 145994
rect 114008 145930 114060 145936
rect 114112 141982 114140 259490
rect 114100 141976 114152 141982
rect 114100 141918 114152 141924
rect 114204 141914 114232 260238
rect 115020 259752 115072 259758
rect 115020 259694 115072 259700
rect 114468 199572 114520 199578
rect 114468 199514 114520 199520
rect 114376 199504 114428 199510
rect 114376 199446 114428 199452
rect 114284 196852 114336 196858
rect 114284 196794 114336 196800
rect 114192 141908 114244 141914
rect 114192 141850 114244 141856
rect 114006 138952 114062 138961
rect 114006 138887 114062 138896
rect 113916 80844 113968 80850
rect 113916 80786 113968 80792
rect 113916 78736 113968 78742
rect 113916 78678 113968 78684
rect 113928 78606 113956 78678
rect 113916 78600 113968 78606
rect 113916 78542 113968 78548
rect 113824 76628 113876 76634
rect 113824 76570 113876 76576
rect 113548 69896 113600 69902
rect 113548 69838 113600 69844
rect 113548 56568 113600 56574
rect 113548 56510 113600 56516
rect 113560 56001 113588 56510
rect 113546 55992 113602 56001
rect 113546 55927 113602 55936
rect 113192 16546 113772 16574
rect 112812 4140 112864 4146
rect 112812 4082 112864 4088
rect 111616 3392 111668 3398
rect 111616 3334 111668 3340
rect 112444 3392 112496 3398
rect 112444 3334 112496 3340
rect 111628 480 111656 3334
rect 112824 480 112852 4082
rect 113744 3482 113772 16546
rect 113836 4146 113864 76570
rect 114020 68542 114048 138887
rect 114098 138408 114154 138417
rect 114098 138343 114154 138352
rect 114008 68536 114060 68542
rect 114112 68513 114140 138343
rect 114296 76974 114324 196794
rect 114284 76968 114336 76974
rect 114284 76910 114336 76916
rect 114388 76770 114416 199446
rect 114480 77042 114508 199514
rect 114928 148640 114980 148646
rect 114928 148582 114980 148588
rect 114940 80986 114968 148582
rect 115032 142089 115060 259694
rect 115124 154222 115152 262375
rect 115294 259720 115350 259729
rect 115294 259655 115350 259664
rect 115204 259480 115256 259486
rect 115204 259422 115256 259428
rect 115112 154216 115164 154222
rect 115112 154158 115164 154164
rect 115112 151700 115164 151706
rect 115112 151642 115164 151648
rect 115018 142080 115074 142089
rect 115018 142015 115074 142024
rect 115020 140276 115072 140282
rect 115020 140218 115072 140224
rect 114928 80980 114980 80986
rect 114928 80922 114980 80928
rect 115032 78713 115060 140218
rect 115018 78704 115074 78713
rect 115018 78639 115074 78648
rect 114468 77036 114520 77042
rect 114468 76978 114520 76984
rect 114376 76764 114428 76770
rect 114376 76706 114428 76712
rect 114560 76560 114612 76566
rect 114560 76502 114612 76508
rect 114572 75138 114600 76502
rect 114560 75132 114612 75138
rect 114560 75074 114612 75080
rect 114008 68478 114060 68484
rect 114098 68504 114154 68513
rect 114098 68439 114154 68448
rect 114572 16574 114600 75074
rect 115124 70446 115152 151642
rect 115216 148918 115244 259422
rect 115204 148912 115256 148918
rect 115204 148854 115256 148860
rect 115204 145716 115256 145722
rect 115204 145658 115256 145664
rect 115216 78946 115244 145658
rect 115308 144129 115336 259655
rect 115400 146062 115428 262822
rect 115480 262812 115532 262818
rect 115480 262754 115532 262760
rect 115388 146056 115440 146062
rect 115388 145998 115440 146004
rect 115492 144702 115520 262754
rect 116492 262268 116544 262274
rect 116492 262210 116544 262216
rect 115756 199164 115808 199170
rect 115756 199106 115808 199112
rect 115664 195560 115716 195566
rect 115664 195502 115716 195508
rect 115572 148572 115624 148578
rect 115572 148514 115624 148520
rect 115480 144696 115532 144702
rect 115480 144638 115532 144644
rect 115294 144120 115350 144129
rect 115294 144055 115350 144064
rect 115296 143268 115348 143274
rect 115296 143210 115348 143216
rect 115204 78940 115256 78946
rect 115204 78882 115256 78888
rect 115308 76906 115336 143210
rect 115388 140412 115440 140418
rect 115388 140354 115440 140360
rect 115296 76900 115348 76906
rect 115296 76842 115348 76848
rect 115400 74322 115428 140354
rect 115584 79150 115612 148514
rect 115572 79144 115624 79150
rect 115572 79086 115624 79092
rect 115388 74316 115440 74322
rect 115388 74258 115440 74264
rect 115676 73030 115704 195502
rect 115768 75449 115796 199106
rect 115848 199028 115900 199034
rect 115848 198970 115900 198976
rect 115754 75440 115810 75449
rect 115754 75375 115810 75384
rect 115664 73024 115716 73030
rect 115860 73001 115888 198970
rect 116308 148504 116360 148510
rect 116308 148446 116360 148452
rect 116216 147212 116268 147218
rect 116216 147154 116268 147160
rect 115664 72966 115716 72972
rect 115846 72992 115902 73001
rect 115846 72927 115902 72936
rect 115112 70440 115164 70446
rect 115112 70382 115164 70388
rect 115124 69834 115152 70382
rect 115112 69828 115164 69834
rect 115112 69770 115164 69776
rect 116228 68406 116256 147154
rect 116320 79218 116348 148446
rect 116504 142225 116532 262210
rect 116596 154358 116624 265066
rect 119620 264988 119672 264994
rect 119620 264930 119672 264936
rect 118700 264240 118752 264246
rect 118700 264182 118752 264188
rect 117964 263764 118016 263770
rect 117964 263706 118016 263712
rect 116860 263152 116912 263158
rect 116860 263094 116912 263100
rect 116676 262948 116728 262954
rect 116676 262890 116728 262896
rect 116584 154352 116636 154358
rect 116584 154294 116636 154300
rect 116688 144906 116716 262890
rect 116768 261112 116820 261118
rect 116768 261054 116820 261060
rect 116676 144900 116728 144906
rect 116676 144842 116728 144848
rect 116780 143206 116808 261054
rect 116872 144226 116900 263094
rect 117044 263016 117096 263022
rect 117044 262958 117096 262964
rect 116952 148844 117004 148850
rect 116952 148786 117004 148792
rect 116860 144220 116912 144226
rect 116860 144162 116912 144168
rect 116858 143984 116914 143993
rect 116858 143919 116914 143928
rect 116768 143200 116820 143206
rect 116768 143142 116820 143148
rect 116872 142866 116900 143919
rect 116860 142860 116912 142866
rect 116860 142802 116912 142808
rect 116490 142216 116546 142225
rect 116490 142151 116546 142160
rect 116584 141364 116636 141370
rect 116584 141306 116636 141312
rect 116400 140956 116452 140962
rect 116400 140898 116452 140904
rect 116412 80889 116440 140898
rect 116490 139904 116546 139913
rect 116490 139839 116546 139848
rect 116398 80880 116454 80889
rect 116398 80815 116454 80824
rect 116308 79212 116360 79218
rect 116308 79154 116360 79160
rect 116504 78849 116532 139839
rect 116490 78840 116546 78849
rect 116490 78775 116546 78784
rect 116596 75546 116624 141306
rect 116860 139936 116912 139942
rect 116860 139878 116912 139884
rect 116674 138136 116730 138145
rect 116674 138071 116730 138080
rect 116584 75540 116636 75546
rect 116584 75482 116636 75488
rect 116688 72865 116716 138071
rect 116674 72856 116730 72865
rect 116674 72791 116730 72800
rect 116872 71466 116900 139878
rect 116964 75313 116992 148786
rect 117056 142118 117084 262958
rect 117872 259820 117924 259826
rect 117872 259762 117924 259768
rect 117780 259616 117832 259622
rect 117780 259558 117832 259564
rect 117228 199232 117280 199238
rect 117228 199174 117280 199180
rect 117136 195696 117188 195702
rect 117136 195638 117188 195644
rect 117044 142112 117096 142118
rect 117044 142054 117096 142060
rect 117044 141024 117096 141030
rect 117044 140966 117096 140972
rect 117056 140214 117084 140966
rect 117044 140208 117096 140214
rect 117044 140150 117096 140156
rect 116950 75304 117006 75313
rect 116950 75239 117006 75248
rect 117148 72758 117176 195638
rect 117240 75410 117268 199174
rect 117792 189038 117820 259558
rect 117780 189032 117832 189038
rect 117780 188974 117832 188980
rect 117688 147484 117740 147490
rect 117688 147426 117740 147432
rect 117596 144016 117648 144022
rect 117596 143958 117648 143964
rect 117228 75404 117280 75410
rect 117228 75346 117280 75352
rect 117136 72752 117188 72758
rect 117136 72694 117188 72700
rect 116860 71460 116912 71466
rect 116860 71402 116912 71408
rect 117320 69760 117372 69766
rect 117320 69702 117372 69708
rect 116216 68400 116268 68406
rect 116216 68342 116268 68348
rect 116228 64874 116256 68342
rect 115952 64846 116256 64874
rect 115952 16574 115980 64846
rect 114572 16546 114784 16574
rect 115952 16546 116440 16574
rect 113824 4140 113876 4146
rect 113824 4082 113876 4088
rect 113744 3454 114048 3482
rect 114020 480 114048 3454
rect 109286 354 109398 480
rect 109052 326 109398 354
rect 109286 -960 109398 326
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 116412 480 116440 16546
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117332 354 117360 69702
rect 117608 67386 117636 143958
rect 117700 69737 117728 147426
rect 117884 144430 117912 259762
rect 117976 146130 118004 263706
rect 118712 263634 118740 264182
rect 119528 263900 119580 263906
rect 119528 263842 119580 263848
rect 118700 263628 118752 263634
rect 118700 263570 118752 263576
rect 118332 262744 118384 262750
rect 118332 262686 118384 262692
rect 118240 262676 118292 262682
rect 118240 262618 118292 262624
rect 118148 260228 118200 260234
rect 118148 260170 118200 260176
rect 118056 260092 118108 260098
rect 118056 260034 118108 260040
rect 117964 146124 118016 146130
rect 117964 146066 118016 146072
rect 117964 145784 118016 145790
rect 117964 145726 118016 145732
rect 117872 144424 117924 144430
rect 117872 144366 117924 144372
rect 117872 136196 117924 136202
rect 117872 136138 117924 136144
rect 117778 92440 117834 92449
rect 117778 92375 117834 92384
rect 117792 69766 117820 92375
rect 117884 81161 117912 136138
rect 117870 81152 117926 81161
rect 117870 81087 117926 81096
rect 117976 80918 118004 145726
rect 118068 142050 118096 260034
rect 118056 142044 118108 142050
rect 118056 141986 118108 141992
rect 118160 141778 118188 260170
rect 118252 143546 118280 262618
rect 118240 143540 118292 143546
rect 118240 143482 118292 143488
rect 118344 143410 118372 262686
rect 119252 260772 119304 260778
rect 119252 260714 119304 260720
rect 118608 199368 118660 199374
rect 118608 199310 118660 199316
rect 118424 199300 118476 199306
rect 118424 199242 118476 199248
rect 118332 143404 118384 143410
rect 118332 143346 118384 143352
rect 118148 141772 118200 141778
rect 118148 141714 118200 141720
rect 118148 140616 118200 140622
rect 118148 140558 118200 140564
rect 118056 140548 118108 140554
rect 118056 140490 118108 140496
rect 117964 80912 118016 80918
rect 117964 80854 118016 80860
rect 118068 79082 118096 140490
rect 118056 79076 118108 79082
rect 118056 79018 118108 79024
rect 118160 71534 118188 140558
rect 118332 140412 118384 140418
rect 118332 140354 118384 140360
rect 118344 140010 118372 140354
rect 118332 140004 118384 140010
rect 118332 139946 118384 139952
rect 118436 76809 118464 199242
rect 118516 195764 118568 195770
rect 118516 195706 118568 195712
rect 118422 76800 118478 76809
rect 118422 76735 118478 76744
rect 118528 72622 118556 195706
rect 118620 75274 118648 199310
rect 119068 197124 119120 197130
rect 119068 197066 119120 197072
rect 118792 144968 118844 144974
rect 118792 144910 118844 144916
rect 118804 140729 118832 144910
rect 118884 144560 118936 144566
rect 118884 144502 118936 144508
rect 118790 140720 118846 140729
rect 118790 140655 118846 140664
rect 118700 139528 118752 139534
rect 118700 139470 118752 139476
rect 118712 137970 118740 139470
rect 118700 137964 118752 137970
rect 118700 137906 118752 137912
rect 118608 75268 118660 75274
rect 118608 75210 118660 75216
rect 118516 72616 118568 72622
rect 118516 72558 118568 72564
rect 118148 71528 118200 71534
rect 118148 71470 118200 71476
rect 118896 70310 118924 144502
rect 119080 74050 119108 197066
rect 119264 149122 119292 260714
rect 119344 259888 119396 259894
rect 119344 259830 119396 259836
rect 119434 259856 119490 259865
rect 119252 149116 119304 149122
rect 119252 149058 119304 149064
rect 119356 143002 119384 259830
rect 119434 259791 119490 259800
rect 119344 142996 119396 143002
rect 119344 142938 119396 142944
rect 119448 142934 119476 259791
rect 119540 144770 119568 263842
rect 119528 144764 119580 144770
rect 119528 144706 119580 144712
rect 119632 144498 119660 264930
rect 121000 263968 121052 263974
rect 121000 263910 121052 263916
rect 120908 263832 120960 263838
rect 120908 263774 120960 263780
rect 119712 263696 119764 263702
rect 119712 263638 119764 263644
rect 119620 144492 119672 144498
rect 119620 144434 119672 144440
rect 119724 143070 119752 263638
rect 119988 263628 120040 263634
rect 119988 263570 120040 263576
rect 119804 262540 119856 262546
rect 119804 262482 119856 262488
rect 119712 143064 119764 143070
rect 119712 143006 119764 143012
rect 119436 142928 119488 142934
rect 119436 142870 119488 142876
rect 119816 141574 119844 262482
rect 119896 260840 119948 260846
rect 119896 260782 119948 260788
rect 119908 199918 119936 260782
rect 119896 199912 119948 199918
rect 119896 199854 119948 199860
rect 119896 195832 119948 195838
rect 120000 195809 120028 263570
rect 120814 262712 120870 262721
rect 120814 262647 120870 262656
rect 120632 259956 120684 259962
rect 120632 259898 120684 259904
rect 119896 195774 119948 195780
rect 119986 195800 120042 195809
rect 119804 141568 119856 141574
rect 119804 141510 119856 141516
rect 119252 141500 119304 141506
rect 119252 141442 119304 141448
rect 119160 140480 119212 140486
rect 119160 140422 119212 140428
rect 119172 79286 119200 140422
rect 119264 79558 119292 141442
rect 119620 141432 119672 141438
rect 119620 141374 119672 141380
rect 119434 140584 119490 140593
rect 119434 140519 119490 140528
rect 119342 136640 119398 136649
rect 119342 136575 119398 136584
rect 119252 79552 119304 79558
rect 119252 79494 119304 79500
rect 119160 79280 119212 79286
rect 119160 79222 119212 79228
rect 119068 74044 119120 74050
rect 119068 73986 119120 73992
rect 119356 73914 119384 136575
rect 119448 74458 119476 140519
rect 119526 140176 119582 140185
rect 119526 140111 119582 140120
rect 119436 74452 119488 74458
rect 119436 74394 119488 74400
rect 119344 73908 119396 73914
rect 119344 73850 119396 73856
rect 119540 71369 119568 140111
rect 119526 71360 119582 71369
rect 119632 71330 119660 141374
rect 119804 140548 119856 140554
rect 119804 140490 119856 140496
rect 119712 140140 119764 140146
rect 119712 140082 119764 140088
rect 119526 71295 119582 71304
rect 119620 71324 119672 71330
rect 119620 71266 119672 71272
rect 118884 70304 118936 70310
rect 118884 70246 118936 70252
rect 117780 69760 117832 69766
rect 117686 69728 117742 69737
rect 117780 69702 117832 69708
rect 117686 69663 117742 69672
rect 117596 67380 117648 67386
rect 117596 67322 117648 67328
rect 119724 65890 119752 140082
rect 119816 136202 119844 140490
rect 119804 136196 119856 136202
rect 119804 136138 119856 136144
rect 119908 72729 119936 195774
rect 119986 195735 120042 195744
rect 119988 149116 120040 149122
rect 119988 149058 120040 149064
rect 120000 141370 120028 149058
rect 120446 147656 120502 147665
rect 120446 147591 120502 147600
rect 120356 146192 120408 146198
rect 120356 146134 120408 146140
rect 120264 144628 120316 144634
rect 120264 144570 120316 144576
rect 119988 141364 120040 141370
rect 119988 141306 120040 141312
rect 120276 137358 120304 144570
rect 120264 137352 120316 137358
rect 120264 137294 120316 137300
rect 119894 72720 119950 72729
rect 119894 72655 119950 72664
rect 120172 68332 120224 68338
rect 120172 68274 120224 68280
rect 119712 65884 119764 65890
rect 119712 65826 119764 65832
rect 120078 52592 120134 52601
rect 120078 52527 120134 52536
rect 120092 3398 120120 52527
rect 120080 3392 120132 3398
rect 120080 3334 120132 3340
rect 120184 3210 120212 68274
rect 120368 67454 120396 146134
rect 120356 67448 120408 67454
rect 120356 67390 120408 67396
rect 120460 55049 120488 147591
rect 120644 145858 120672 259898
rect 120724 195968 120776 195974
rect 120724 195910 120776 195916
rect 120632 145852 120684 145858
rect 120632 145794 120684 145800
rect 120540 140684 120592 140690
rect 120540 140626 120592 140632
rect 120552 79354 120580 140626
rect 120632 137352 120684 137358
rect 120632 137294 120684 137300
rect 120540 79348 120592 79354
rect 120540 79290 120592 79296
rect 120644 74633 120672 137294
rect 120736 78130 120764 195910
rect 120828 144537 120856 262647
rect 120814 144528 120870 144537
rect 120814 144463 120870 144472
rect 120920 143138 120948 263774
rect 121012 143342 121040 263910
rect 129280 263152 129332 263158
rect 129280 263094 129332 263100
rect 125968 263016 126020 263022
rect 125968 262958 126020 262964
rect 122840 262744 122892 262750
rect 122840 262686 122892 262692
rect 122852 262410 122880 262686
rect 122840 262404 122892 262410
rect 122840 262346 122892 262352
rect 122748 262268 122800 262274
rect 122748 262210 122800 262216
rect 122760 260710 122788 262210
rect 125598 261216 125654 261225
rect 125598 261151 125654 261160
rect 124312 260840 124364 260846
rect 124312 260782 124364 260788
rect 122840 260772 122892 260778
rect 122840 260714 122892 260720
rect 122748 260704 122800 260710
rect 122748 260646 122800 260652
rect 122852 259978 122880 260714
rect 123208 260704 123260 260710
rect 123208 260646 123260 260652
rect 123220 259978 123248 260646
rect 124324 259978 124352 260782
rect 125612 259978 125640 261151
rect 125980 259978 126008 262958
rect 127532 262948 127584 262954
rect 127532 262890 127584 262896
rect 127544 262750 127572 262890
rect 127532 262744 127584 262750
rect 127532 262686 127584 262692
rect 127624 262676 127676 262682
rect 127624 262618 127676 262624
rect 127072 261044 127124 261050
rect 127072 260986 127124 260992
rect 126520 260296 126572 260302
rect 126520 260238 126572 260244
rect 126532 259978 126560 260238
rect 127084 259978 127112 260986
rect 127636 259978 127664 262618
rect 128728 261180 128780 261186
rect 128728 261122 128780 261128
rect 128740 259978 128768 261122
rect 129292 259978 129320 263094
rect 132316 263016 132368 263022
rect 132316 262958 132368 262964
rect 131764 262880 131816 262886
rect 131764 262822 131816 262828
rect 129832 262608 129884 262614
rect 129832 262550 129884 262556
rect 129844 261594 129872 262550
rect 131120 262404 131172 262410
rect 131120 262346 131172 262352
rect 129832 261588 129884 261594
rect 129832 261530 129884 261536
rect 129844 259978 129872 261530
rect 131132 261458 131160 262346
rect 131120 261452 131172 261458
rect 131120 261394 131172 261400
rect 130384 260908 130436 260914
rect 130384 260850 130436 260856
rect 130396 259978 130424 260850
rect 131132 259978 131160 261394
rect 131776 259978 131804 262822
rect 132040 260024 132092 260030
rect 122852 259950 123004 259978
rect 123220 259950 123556 259978
rect 124324 259950 124660 259978
rect 125612 259950 125764 259978
rect 125980 259950 126316 259978
rect 126532 259950 126868 259978
rect 127084 259950 127420 259978
rect 127636 259950 127972 259978
rect 128740 259950 129076 259978
rect 129292 259950 129628 259978
rect 129844 259950 130180 259978
rect 130396 259950 130732 259978
rect 131132 259950 131284 259978
rect 131776 259950 131836 259978
rect 132040 259966 132092 259972
rect 132052 259842 132080 259966
rect 132328 259842 132356 262958
rect 133156 262750 133184 271866
rect 134248 263968 134300 263974
rect 134248 263910 134300 263916
rect 133144 262744 133196 262750
rect 133144 262686 133196 262692
rect 133156 261202 133184 262686
rect 133156 261174 133368 261202
rect 133236 261112 133288 261118
rect 133236 261054 133288 261060
rect 133248 260438 133276 261054
rect 133236 260432 133288 260438
rect 133236 260374 133288 260380
rect 133248 259978 133276 260374
rect 132940 259950 133276 259978
rect 133340 259978 133368 261174
rect 133970 261080 134026 261089
rect 133970 261015 134026 261024
rect 133984 259978 134012 261015
rect 134260 259978 134288 263910
rect 134536 262818 134564 324294
rect 134616 298172 134668 298178
rect 134616 298114 134668 298120
rect 134628 263974 134656 298114
rect 134616 263968 134668 263974
rect 134616 263910 134668 263916
rect 134524 262812 134576 262818
rect 134524 262754 134576 262760
rect 134800 262812 134852 262818
rect 134800 262754 134852 262760
rect 134812 259978 134840 262754
rect 135272 260234 135300 351902
rect 135904 311908 135956 311914
rect 135904 311850 135956 311856
rect 135916 265305 135944 311850
rect 137284 286340 137336 286346
rect 137284 286282 137336 286288
rect 137296 267734 137324 286282
rect 137204 267706 137324 267734
rect 135902 265296 135958 265305
rect 135902 265231 135958 265240
rect 135260 260228 135312 260234
rect 135260 260170 135312 260176
rect 135272 260114 135300 260170
rect 135088 260098 135300 260114
rect 135076 260092 135300 260098
rect 135128 260086 135300 260092
rect 135076 260034 135128 260040
rect 135916 259978 135944 265231
rect 137204 263770 137232 267706
rect 137836 267028 137888 267034
rect 137836 266970 137888 266976
rect 137848 263906 137876 266970
rect 137836 263900 137888 263906
rect 137836 263842 137888 263848
rect 137192 263764 137244 263770
rect 137192 263706 137244 263712
rect 136226 260228 136278 260234
rect 136226 260170 136278 260176
rect 133340 259950 133492 259978
rect 133984 259964 134044 259978
rect 133984 259950 134058 259964
rect 134260 259950 134596 259978
rect 134812 259950 135148 259978
rect 135700 259950 135944 259978
rect 136238 259964 136266 260170
rect 137204 259978 137232 263706
rect 137468 263560 137520 263566
rect 137468 263502 137520 263508
rect 137480 260953 137508 263502
rect 137466 260944 137522 260953
rect 137466 260879 137522 260888
rect 136804 259950 137232 259978
rect 132052 259814 132388 259842
rect 134030 259706 134058 259950
rect 137480 259842 137508 260879
rect 137356 259814 137508 259842
rect 137848 259842 137876 263842
rect 138676 262857 138704 430578
rect 138756 418192 138808 418198
rect 138756 418134 138808 418140
rect 138768 265198 138796 418134
rect 139412 267734 139440 484366
rect 139676 470620 139728 470626
rect 139676 470562 139728 470568
rect 139412 267706 139532 267734
rect 138756 265192 138808 265198
rect 138756 265134 138808 265140
rect 138662 262848 138718 262857
rect 138662 262783 138718 262792
rect 138676 259978 138704 262783
rect 138460 259950 138704 259978
rect 138768 259978 138796 265134
rect 139400 264240 139452 264246
rect 139400 264182 139452 264188
rect 139412 263838 139440 264182
rect 139400 263832 139452 263838
rect 139400 263774 139452 263780
rect 139412 259978 139440 263774
rect 139504 260234 139532 267706
rect 139492 260228 139544 260234
rect 139492 260170 139544 260176
rect 139688 260166 139716 470562
rect 140780 280832 140832 280838
rect 140780 280774 140832 280780
rect 140090 260228 140142 260234
rect 140090 260170 140142 260176
rect 139676 260160 139728 260166
rect 139676 260102 139728 260108
rect 138768 259950 139012 259978
rect 139412 259950 139564 259978
rect 140102 259964 140130 260170
rect 140642 260160 140694 260166
rect 140792 260137 140820 280774
rect 141424 265736 141476 265742
rect 141424 265678 141476 265684
rect 141436 263702 141464 265678
rect 141148 263696 141200 263702
rect 141148 263638 141200 263644
rect 141424 263696 141476 263702
rect 141424 263638 141476 263644
rect 140642 260102 140694 260108
rect 140778 260128 140834 260137
rect 140654 259964 140682 260102
rect 140778 260063 140834 260072
rect 141160 259978 141188 263638
rect 141422 259992 141478 260001
rect 141160 259950 141220 259978
rect 141478 259950 141772 259978
rect 142172 259962 142200 590650
rect 142804 563100 142856 563106
rect 142804 563042 142856 563048
rect 142816 267734 142844 563042
rect 142896 524476 142948 524482
rect 142896 524418 142948 524424
rect 142632 267706 142844 267734
rect 142632 263945 142660 267706
rect 142618 263936 142674 263945
rect 142618 263871 142674 263880
rect 142250 262576 142306 262585
rect 142250 262511 142306 262520
rect 142264 259978 142292 262511
rect 142632 259978 142660 263871
rect 142908 262585 142936 524418
rect 142894 262576 142950 262585
rect 142894 262511 142950 262520
rect 143552 260234 143580 616830
rect 144184 576904 144236 576910
rect 144184 576846 144236 576852
rect 144196 265130 144224 576846
rect 145564 287700 145616 287706
rect 145564 287642 145616 287648
rect 143632 265124 143684 265130
rect 143632 265066 143684 265072
rect 144184 265124 144236 265130
rect 144184 265066 144236 265072
rect 143540 260228 143592 260234
rect 143540 260170 143592 260176
rect 142160 259956 142212 259962
rect 141422 259927 141478 259936
rect 142264 259950 142324 259978
rect 142632 259950 142876 259978
rect 143092 259962 143428 259978
rect 143080 259956 143428 259962
rect 142160 259898 142212 259904
rect 143132 259950 143428 259956
rect 143080 259898 143132 259904
rect 143552 259894 143580 260170
rect 143644 259978 143672 265066
rect 145576 265062 145604 287642
rect 145656 282192 145708 282198
rect 145656 282134 145708 282140
rect 145564 265056 145616 265062
rect 145564 264998 145616 265004
rect 145010 263120 145066 263129
rect 145010 263055 145066 263064
rect 145024 262313 145052 263055
rect 145010 262304 145066 262313
rect 145010 262239 145066 262248
rect 144506 260228 144558 260234
rect 144506 260170 144558 260176
rect 143644 259950 143980 259978
rect 144518 259964 144546 260170
rect 145024 259978 145052 262239
rect 145576 259978 145604 264998
rect 145668 263129 145696 282134
rect 146208 268456 146260 268462
rect 146208 268398 146260 268404
rect 146220 263809 146248 268398
rect 146206 263800 146262 263809
rect 146206 263735 146262 263744
rect 145654 263120 145710 263129
rect 145654 263055 145710 263064
rect 146220 260250 146248 263735
rect 146956 262449 146984 696934
rect 147036 683188 147088 683194
rect 147036 683130 147088 683136
rect 147048 265033 147076 683130
rect 147680 283620 147732 283626
rect 147680 283562 147732 283568
rect 147034 265024 147090 265033
rect 147034 264959 147090 264968
rect 146942 262440 146998 262449
rect 146942 262375 146998 262384
rect 146174 260222 146248 260250
rect 145024 259950 145084 259978
rect 145576 259950 145636 259978
rect 146174 259964 146202 260222
rect 146956 259978 146984 262375
rect 146740 259950 146984 259978
rect 147048 259978 147076 264959
rect 147692 260273 147720 283562
rect 147772 269816 147824 269822
rect 147772 269758 147824 269764
rect 147678 260264 147734 260273
rect 147678 260199 147734 260208
rect 147784 259978 147812 269758
rect 148336 267734 148364 700266
rect 149060 660340 149112 660346
rect 149060 660282 149112 660288
rect 148336 267706 148548 267734
rect 148520 265169 148548 267706
rect 148506 265160 148562 265169
rect 148506 265095 148562 265104
rect 148368 260264 148424 260273
rect 148368 260199 148424 260208
rect 147048 259950 147292 259978
rect 147784 259950 147844 259978
rect 143540 259888 143592 259894
rect 137848 259814 137908 259842
rect 143540 259830 143592 259836
rect 147678 259856 147734 259865
rect 147784 259842 147812 259950
rect 147734 259814 147812 259842
rect 147678 259791 147734 259800
rect 148138 259720 148194 259729
rect 123772 259690 124108 259706
rect 134030 259692 134380 259706
rect 123760 259684 124108 259690
rect 123812 259678 124108 259684
rect 134044 259690 134380 259692
rect 134044 259684 134392 259690
rect 134044 259678 134340 259684
rect 123760 259626 123812 259632
rect 148382 259706 148410 260199
rect 148520 259978 148548 265095
rect 148520 259950 148948 259978
rect 149072 259758 149100 660282
rect 150440 284980 150492 284986
rect 150440 284922 150492 284928
rect 149152 271176 149204 271182
rect 149152 271118 149204 271124
rect 149164 259978 149192 271118
rect 149164 259950 149500 259978
rect 148194 259692 148410 259706
rect 149060 259752 149112 259758
rect 149060 259694 149112 259700
rect 148194 259678 148396 259692
rect 148138 259655 148194 259664
rect 134340 259626 134392 259632
rect 149256 259593 149284 259950
rect 150452 259826 150480 284922
rect 151818 274680 151874 274689
rect 151818 274615 151874 274624
rect 151084 273964 151136 273970
rect 151084 273906 151136 273912
rect 151096 263673 151124 273906
rect 151832 267734 151860 274615
rect 151832 267706 152412 267734
rect 152188 264988 152240 264994
rect 152188 264930 152240 264936
rect 151082 263664 151138 263673
rect 151082 263599 151138 263608
rect 150530 262712 150586 262721
rect 150530 262647 150586 262656
rect 150544 259978 150572 262647
rect 151096 259978 151124 263599
rect 152200 259978 152228 264930
rect 152384 259978 152412 267706
rect 152476 264994 152504 700334
rect 152464 264988 152516 264994
rect 152464 264930 152516 264936
rect 153212 262818 153240 702406
rect 157984 700868 158036 700874
rect 157984 700810 158036 700816
rect 155960 700800 156012 700806
rect 155960 700742 156012 700748
rect 154580 700664 154632 700670
rect 154580 700606 154632 700612
rect 153844 700460 153896 700466
rect 153844 700402 153896 700408
rect 153292 276072 153344 276078
rect 153292 276014 153344 276020
rect 153304 267734 153332 276014
rect 153304 267706 153792 267734
rect 153200 262812 153252 262818
rect 153200 262754 153252 262760
rect 153292 262540 153344 262546
rect 153292 262482 153344 262488
rect 153304 259978 153332 262482
rect 153658 262440 153714 262449
rect 153658 262375 153714 262384
rect 153672 259978 153700 262375
rect 153764 260114 153792 267706
rect 153856 262546 153884 700402
rect 153844 262540 153896 262546
rect 153844 262482 153896 262488
rect 153764 260086 154068 260114
rect 154040 259978 154068 260086
rect 154592 259978 154620 700606
rect 155868 262608 155920 262614
rect 155868 262550 155920 262556
rect 155880 259978 155908 262550
rect 155972 260234 156000 700742
rect 156052 277432 156104 277438
rect 156052 277374 156104 277380
rect 155960 260228 156012 260234
rect 155960 260170 156012 260176
rect 150544 259950 150604 259978
rect 151096 259950 151156 259978
rect 152200 259950 152260 259978
rect 152384 259950 152812 259978
rect 153304 259950 153364 259978
rect 153672 259950 153916 259978
rect 154040 259950 154468 259978
rect 154592 259950 155264 259978
rect 155572 259950 155908 259978
rect 156064 259978 156092 277374
rect 157892 263696 157944 263702
rect 157892 263638 157944 263644
rect 157156 262540 157208 262546
rect 157156 262482 157208 262488
rect 156650 260228 156702 260234
rect 156650 260170 156702 260176
rect 156662 259978 156690 260170
rect 157168 259978 157196 262482
rect 157904 259978 157932 263638
rect 157996 262682 158024 700810
rect 160744 700732 160796 700738
rect 160744 700674 160796 700680
rect 158628 447840 158680 447846
rect 158628 447782 158680 447788
rect 158640 263702 158668 447782
rect 160100 279472 160152 279478
rect 160100 279414 160152 279420
rect 158812 269884 158864 269890
rect 158812 269826 158864 269832
rect 158628 263696 158680 263702
rect 158628 263638 158680 263644
rect 158720 262812 158772 262818
rect 158720 262754 158772 262760
rect 157984 262676 158036 262682
rect 157984 262618 158036 262624
rect 156064 259950 156124 259978
rect 156662 259964 157012 259978
rect 156676 259950 157012 259964
rect 157168 259950 157228 259978
rect 157780 259950 157932 259978
rect 157996 259978 158024 262618
rect 158732 261662 158760 262754
rect 158824 262721 158852 269826
rect 159088 263628 159140 263634
rect 159088 263570 159140 263576
rect 158810 262712 158866 262721
rect 158810 262647 158866 262656
rect 158720 261656 158772 261662
rect 158720 261598 158772 261604
rect 158732 259978 158760 261598
rect 159100 259978 159128 263570
rect 159914 262712 159970 262721
rect 159914 262647 159970 262656
rect 159928 259978 159956 262647
rect 160112 260001 160140 279414
rect 160756 267734 160784 700674
rect 162216 700596 162268 700602
rect 162216 700538 162268 700544
rect 162124 700528 162176 700534
rect 162124 700470 162176 700476
rect 161480 683256 161532 683262
rect 161480 683198 161532 683204
rect 160756 267706 160876 267734
rect 160848 265062 160876 267706
rect 160836 265056 160888 265062
rect 160836 264998 160888 265004
rect 160098 259992 160154 260001
rect 157996 259950 158332 259978
rect 158732 259950 158884 259978
rect 159100 259950 159436 259978
rect 159928 259950 159988 259978
rect 151372 259826 151708 259842
rect 150440 259820 150492 259826
rect 150440 259762 150492 259768
rect 151360 259820 151708 259826
rect 151412 259814 151708 259820
rect 151360 259762 151412 259768
rect 149704 259752 149756 259758
rect 149756 259700 150052 259706
rect 149704 259694 150052 259700
rect 149716 259678 150052 259694
rect 155236 259593 155264 259950
rect 156984 259758 157012 259950
rect 160848 259978 160876 264998
rect 161492 260817 161520 683198
rect 162136 267734 162164 700470
rect 162044 267706 162164 267734
rect 162044 262585 162072 267706
rect 162228 265198 162256 700538
rect 163504 670744 163556 670750
rect 163504 670686 163556 670692
rect 162216 265192 162268 265198
rect 162216 265134 162268 265140
rect 162030 262576 162086 262585
rect 162030 262511 162086 262520
rect 161478 260808 161534 260817
rect 161478 260743 161534 260752
rect 160540 259950 160876 259978
rect 160926 259992 160982 260001
rect 160098 259927 160154 259936
rect 162044 259978 162072 262511
rect 162228 260250 162256 265134
rect 163516 265033 163544 670686
rect 163596 656940 163648 656946
rect 163596 656882 163648 656888
rect 163502 265024 163558 265033
rect 163502 264959 163558 264968
rect 163412 263288 163464 263294
rect 163412 263230 163464 263236
rect 163424 262750 163452 263230
rect 163412 262744 163464 262750
rect 163412 262686 163464 262692
rect 162674 260808 162730 260817
rect 162674 260743 162730 260752
rect 160982 259964 161092 259978
rect 160982 259950 161106 259964
rect 161644 259950 162072 259978
rect 162182 260222 162256 260250
rect 162182 259964 162210 260222
rect 160926 259927 160982 259936
rect 156972 259752 157024 259758
rect 156972 259694 157024 259700
rect 161078 259706 161106 259950
rect 162582 259856 162638 259865
rect 162688 259842 162716 260743
rect 163424 259978 163452 262686
rect 163300 259950 163452 259978
rect 163516 259978 163544 264959
rect 163608 263294 163636 656882
rect 164240 632120 164292 632126
rect 164240 632062 164292 632068
rect 163596 263288 163648 263294
rect 163596 263230 163648 263236
rect 164252 260302 164280 632062
rect 164884 618316 164936 618322
rect 164884 618258 164936 618264
rect 164896 265878 164924 618258
rect 164976 605872 165028 605878
rect 164976 605814 165028 605820
rect 164884 265872 164936 265878
rect 164884 265814 164936 265820
rect 164988 262818 165016 605814
rect 165620 579692 165672 579698
rect 165620 579634 165672 579640
rect 165160 265872 165212 265878
rect 165160 265814 165212 265820
rect 165172 264994 165200 265814
rect 165160 264988 165212 264994
rect 165160 264930 165212 264936
rect 164976 262812 165028 262818
rect 164976 262754 165028 262760
rect 164240 260296 164292 260302
rect 164988 260250 165016 262754
rect 164240 260238 164292 260244
rect 164252 259978 164280 260238
rect 164942 260222 165016 260250
rect 163516 259950 163852 259978
rect 164252 259950 164404 259978
rect 164942 259964 164970 260222
rect 165172 259978 165200 264930
rect 165632 259978 165660 579634
rect 167644 565888 167696 565894
rect 167644 565830 167696 565836
rect 166264 553444 166316 553450
rect 166264 553386 166316 553392
rect 166276 265470 166304 553386
rect 167000 527196 167052 527202
rect 167000 527138 167052 527144
rect 166264 265464 166316 265470
rect 166264 265406 166316 265412
rect 166276 259978 166304 265406
rect 167012 260166 167040 527138
rect 167276 501016 167328 501022
rect 167276 500958 167328 500964
rect 167288 260234 167316 500958
rect 167656 267734 167684 565830
rect 169772 447846 169800 702406
rect 202800 700806 202828 703520
rect 202788 700800 202840 700806
rect 202788 700742 202840 700748
rect 185584 670744 185636 670750
rect 185584 670686 185636 670692
rect 184204 643136 184256 643142
rect 184204 643078 184256 643084
rect 178684 536852 178736 536858
rect 178684 536794 178736 536800
rect 170404 462392 170456 462398
rect 170404 462334 170456 462340
rect 169760 447840 169812 447846
rect 169760 447782 169812 447788
rect 169760 422340 169812 422346
rect 169760 422282 169812 422288
rect 169024 274032 169076 274038
rect 169024 273974 169076 273980
rect 167564 267706 167684 267734
rect 167564 265169 167592 267706
rect 169036 265305 169064 273974
rect 169116 265668 169168 265674
rect 169116 265610 169168 265616
rect 169022 265296 169078 265305
rect 169022 265231 169078 265240
rect 167550 265160 167606 265169
rect 167550 265095 167606 265104
rect 167276 260228 167328 260234
rect 167276 260170 167328 260176
rect 167000 260160 167052 260166
rect 167000 260102 167052 260108
rect 167564 259978 167592 265095
rect 168242 260228 168294 260234
rect 168242 260170 168294 260176
rect 167690 260160 167742 260166
rect 167690 260102 167742 260108
rect 165172 259950 165508 259978
rect 165632 259950 166212 259978
rect 166276 259950 166612 259978
rect 167164 259950 167592 259978
rect 167702 259964 167730 260102
rect 168254 259978 168282 260170
rect 169036 259978 169064 265231
rect 168254 259964 168420 259978
rect 168268 259962 168420 259964
rect 168268 259956 168432 259962
rect 168268 259950 168380 259956
rect 166184 259894 166212 259950
rect 168820 259950 169064 259978
rect 169128 259978 169156 265610
rect 169772 260234 169800 422282
rect 170416 265266 170444 462334
rect 170496 448588 170548 448594
rect 170496 448530 170548 448536
rect 170404 265260 170456 265266
rect 170404 265202 170456 265208
rect 170508 265130 170536 448530
rect 171784 409896 171836 409902
rect 171784 409838 171836 409844
rect 171796 265402 171824 409838
rect 171876 397520 171928 397526
rect 171876 397462 171928 397468
rect 171784 265396 171836 265402
rect 171784 265338 171836 265344
rect 170680 265260 170732 265266
rect 170680 265202 170732 265208
rect 170220 265124 170272 265130
rect 170220 265066 170272 265072
rect 170496 265124 170548 265130
rect 170496 265066 170548 265072
rect 169760 260228 169812 260234
rect 169760 260170 169812 260176
rect 169346 260092 169398 260098
rect 169346 260034 169398 260040
rect 169358 259978 169386 260034
rect 170232 259978 170260 265066
rect 170692 259978 170720 265202
rect 171692 263424 171744 263430
rect 171692 263366 171744 263372
rect 171704 263158 171732 263366
rect 171692 263152 171744 263158
rect 171692 263094 171744 263100
rect 171002 260228 171054 260234
rect 171002 260170 171054 260176
rect 169128 259964 169386 259978
rect 169128 259950 169372 259964
rect 169924 259950 170260 259978
rect 170476 259950 170720 259978
rect 168380 259898 168432 259904
rect 166172 259888 166224 259894
rect 162638 259814 162748 259842
rect 166172 259830 166224 259836
rect 171014 259842 171042 260170
rect 171704 259978 171732 263094
rect 171580 259950 171732 259978
rect 171796 259978 171824 265338
rect 171888 263430 171916 397462
rect 173900 318844 173952 318850
rect 173900 318786 173952 318792
rect 173164 289128 173216 289134
rect 173164 289070 173216 289076
rect 172520 271244 172572 271250
rect 172520 271186 172572 271192
rect 171876 263424 171928 263430
rect 171876 263366 171928 263372
rect 172532 260234 172560 271186
rect 172704 268388 172756 268394
rect 172704 268330 172756 268336
rect 172716 263770 172744 268330
rect 173176 267734 173204 289070
rect 173176 267706 173480 267734
rect 173452 265334 173480 267706
rect 173440 265328 173492 265334
rect 173440 265270 173492 265276
rect 172704 263764 172756 263770
rect 172704 263706 172756 263712
rect 172716 260250 172744 263706
rect 172520 260228 172572 260234
rect 172520 260170 172572 260176
rect 172670 260222 172744 260250
rect 173210 260228 173262 260234
rect 171796 259950 172132 259978
rect 172670 259964 172698 260222
rect 173210 260170 173262 260176
rect 173222 259978 173250 260170
rect 173452 259978 173480 265270
rect 173912 260506 173940 318786
rect 175924 305040 175976 305046
rect 175924 304982 175976 304988
rect 174544 292596 174596 292602
rect 174544 292538 174596 292544
rect 174556 265606 174584 292538
rect 175936 267734 175964 304982
rect 178696 280838 178724 536794
rect 181444 510672 181496 510678
rect 181444 510614 181496 510620
rect 180064 456816 180116 456822
rect 180064 456758 180116 456764
rect 178684 280832 178736 280838
rect 178684 280774 178736 280780
rect 175752 267706 175964 267734
rect 174544 265600 174596 265606
rect 174544 265542 174596 265548
rect 173900 260500 173952 260506
rect 173900 260442 173952 260448
rect 173912 259978 173940 260442
rect 174556 259978 174584 265542
rect 175752 263634 175780 267706
rect 175924 266416 175976 266422
rect 175924 266358 175976 266364
rect 175740 263628 175792 263634
rect 175740 263570 175792 263576
rect 175752 259978 175780 263570
rect 175832 260296 175884 260302
rect 175832 260238 175884 260244
rect 173222 259964 173388 259978
rect 173236 259950 173388 259964
rect 173452 259950 173788 259978
rect 173912 259950 174340 259978
rect 174556 259950 174892 259978
rect 175444 259950 175780 259978
rect 171014 259828 171180 259842
rect 171028 259826 171180 259828
rect 171028 259820 171192 259826
rect 171028 259814 171140 259820
rect 162582 259791 162638 259800
rect 171140 259762 171192 259768
rect 161202 259720 161258 259729
rect 161078 259692 161202 259706
rect 161092 259678 161202 259692
rect 161202 259655 161258 259664
rect 149242 259584 149298 259593
rect 124876 259554 125212 259570
rect 124864 259548 125212 259554
rect 124916 259542 125212 259548
rect 128372 259542 128524 259570
rect 124864 259490 124916 259496
rect 128372 259486 128400 259542
rect 149242 259519 149298 259528
rect 155222 259584 155278 259593
rect 173360 259554 173388 259950
rect 175844 259894 175872 260238
rect 175936 260234 175964 266358
rect 180076 264246 180104 456758
rect 181456 265742 181484 510614
rect 182824 378208 182876 378214
rect 182824 378150 182876 378156
rect 182836 286346 182864 378150
rect 182824 286340 182876 286346
rect 182824 286282 182876 286288
rect 184216 282198 184244 643078
rect 184204 282192 184256 282198
rect 184204 282134 184256 282140
rect 185596 268462 185624 670686
rect 203524 630692 203576 630698
rect 203524 630634 203576 630640
rect 199384 404388 199436 404394
rect 199384 404330 199436 404336
rect 189080 278044 189132 278050
rect 189080 277986 189132 277992
rect 189092 277438 189120 277986
rect 189080 277432 189132 277438
rect 189080 277374 189132 277380
rect 185584 268456 185636 268462
rect 185584 268398 185636 268404
rect 181444 265736 181496 265742
rect 181444 265678 181496 265684
rect 180064 264240 180116 264246
rect 180064 264182 180116 264188
rect 188252 263696 188304 263702
rect 188252 263638 188304 263644
rect 178408 263084 178460 263090
rect 178408 263026 178460 263032
rect 180156 263084 180208 263090
rect 180156 263026 180208 263032
rect 176752 262472 176804 262478
rect 176752 262414 176804 262420
rect 176764 261526 176792 262414
rect 176752 261520 176804 261526
rect 176752 261462 176804 261468
rect 176200 261180 176252 261186
rect 176200 261122 176252 261128
rect 176212 260982 176240 261122
rect 176200 260976 176252 260982
rect 176200 260918 176252 260924
rect 175924 260228 175976 260234
rect 175924 260170 175976 260176
rect 175936 259978 175964 260170
rect 176212 259978 176240 260918
rect 176764 259978 176792 261462
rect 177304 261316 177356 261322
rect 177304 261258 177356 261264
rect 177316 260370 177344 261258
rect 178420 261254 178448 263026
rect 179236 262472 179288 262478
rect 179236 262414 179288 262420
rect 178408 261248 178460 261254
rect 178408 261190 178460 261196
rect 177304 260364 177356 260370
rect 177304 260306 177356 260312
rect 177316 259978 177344 260306
rect 178420 259978 178448 261190
rect 179248 259978 179276 262414
rect 180168 259978 180196 263026
rect 187698 262984 187754 262993
rect 187698 262919 187754 262928
rect 187712 262449 187740 262919
rect 187698 262440 187754 262449
rect 182916 262404 182968 262410
rect 187698 262375 187754 262384
rect 187974 262440 188030 262449
rect 187974 262375 188030 262384
rect 182916 262346 182968 262352
rect 181260 262336 181312 262342
rect 181260 262278 181312 262284
rect 180524 261044 180576 261050
rect 180524 260986 180576 260992
rect 180536 259978 180564 260986
rect 180800 260568 180852 260574
rect 180800 260510 180852 260516
rect 180812 260166 180840 260510
rect 180800 260160 180852 260166
rect 180800 260102 180852 260108
rect 181272 259978 181300 262278
rect 181812 261384 181864 261390
rect 181812 261326 181864 261332
rect 181824 259978 181852 261326
rect 181996 260908 182048 260914
rect 181996 260850 182048 260856
rect 175936 259950 175996 259978
rect 176212 259950 176548 259978
rect 176764 259950 177100 259978
rect 177316 259950 177652 259978
rect 178420 259950 178756 259978
rect 179248 259950 179308 259978
rect 179860 259950 180196 259978
rect 180412 259950 180564 259978
rect 180964 259950 181300 259978
rect 181516 259950 181852 259978
rect 182008 259978 182036 260850
rect 182928 259978 182956 262346
rect 184572 262268 184624 262274
rect 184572 262210 184624 262216
rect 184020 261112 184072 261118
rect 184020 261054 184072 261060
rect 183468 260024 183520 260030
rect 182008 259950 182068 259978
rect 182620 259950 182956 259978
rect 183296 259972 183468 259978
rect 184032 259978 184060 261054
rect 184584 259978 184612 262210
rect 184756 260976 184808 260982
rect 184756 260918 184808 260924
rect 183296 259966 183520 259972
rect 183296 259962 183508 259966
rect 183284 259956 183508 259962
rect 183336 259950 183508 259956
rect 183724 259950 184060 259978
rect 184276 259950 184612 259978
rect 184768 259978 184796 260918
rect 185584 260500 185636 260506
rect 185584 260442 185636 260448
rect 185596 260302 185624 260442
rect 185584 260296 185636 260302
rect 185584 260238 185636 260244
rect 184768 259950 184828 259978
rect 183284 259898 183336 259904
rect 175832 259888 175884 259894
rect 183468 259888 183520 259894
rect 175832 259830 175884 259836
rect 183172 259836 183468 259842
rect 183172 259830 183520 259836
rect 183172 259814 183508 259830
rect 185768 259752 185820 259758
rect 185768 259694 185820 259700
rect 178040 259616 178092 259622
rect 185674 259584 185730 259593
rect 178092 259564 178204 259570
rect 178040 259558 178204 259564
rect 155222 259519 155278 259528
rect 173348 259548 173400 259554
rect 178052 259542 178204 259558
rect 185380 259542 185674 259570
rect 185674 259519 185730 259528
rect 173348 259490 173400 259496
rect 185780 259486 185808 259694
rect 187700 259684 187752 259690
rect 187700 259626 187752 259632
rect 128360 259480 128412 259486
rect 128360 259422 128412 259428
rect 185768 259480 185820 259486
rect 185768 259422 185820 259428
rect 187712 259418 187740 259626
rect 187700 259412 187752 259418
rect 187700 259354 187752 259360
rect 126244 200728 126296 200734
rect 132224 200728 132276 200734
rect 126244 200670 126296 200676
rect 127714 200696 127770 200705
rect 121368 200388 121420 200394
rect 121368 200330 121420 200336
rect 121276 198892 121328 198898
rect 121276 198834 121328 198840
rect 121092 197260 121144 197266
rect 121092 197202 121144 197208
rect 121000 143336 121052 143342
rect 121000 143278 121052 143284
rect 120998 143168 121054 143177
rect 120908 143132 120960 143138
rect 120998 143103 121054 143112
rect 120908 143074 120960 143080
rect 121012 142254 121040 143103
rect 121000 142248 121052 142254
rect 121000 142190 121052 142196
rect 120816 140752 120868 140758
rect 120816 140694 120868 140700
rect 120724 78124 120776 78130
rect 120724 78066 120776 78072
rect 120630 74624 120686 74633
rect 120630 74559 120686 74568
rect 120828 70038 120856 140694
rect 120998 138544 121054 138553
rect 120998 138479 121054 138488
rect 121012 138038 121040 138479
rect 121000 138032 121052 138038
rect 121000 137974 121052 137980
rect 121104 75138 121132 197202
rect 121182 196752 121238 196761
rect 121182 196687 121238 196696
rect 121092 75132 121144 75138
rect 121092 75074 121144 75080
rect 121196 74118 121224 196687
rect 121184 74112 121236 74118
rect 121184 74054 121236 74060
rect 121288 73098 121316 198834
rect 121380 73166 121408 200330
rect 125140 199912 125192 199918
rect 125140 199854 125192 199860
rect 122380 198484 122432 198490
rect 122380 198426 122432 198432
rect 122288 198348 122340 198354
rect 122288 198290 122340 198296
rect 122196 194200 122248 194206
rect 122196 194142 122248 194148
rect 121828 190460 121880 190466
rect 121828 190402 121880 190408
rect 121736 140616 121788 140622
rect 121736 140558 121788 140564
rect 121748 140078 121776 140558
rect 121736 140072 121788 140078
rect 121736 140014 121788 140020
rect 121734 138136 121790 138145
rect 121734 138071 121790 138080
rect 121748 132569 121776 138071
rect 121840 136649 121868 190402
rect 122104 148776 122156 148782
rect 122104 148718 122156 148724
rect 122010 148064 122066 148073
rect 122010 147999 122066 148008
rect 121920 140616 121972 140622
rect 121920 140558 121972 140564
rect 121826 136640 121882 136649
rect 121826 136575 121882 136584
rect 121734 132560 121790 132569
rect 121734 132495 121790 132504
rect 121826 132424 121882 132433
rect 121826 132359 121882 132368
rect 121840 122913 121868 132359
rect 121826 122904 121882 122913
rect 121826 122839 121882 122848
rect 121826 122768 121882 122777
rect 121826 122703 121882 122712
rect 121840 113257 121868 122703
rect 121826 113248 121882 113257
rect 121826 113183 121882 113192
rect 121826 113112 121882 113121
rect 121826 113047 121882 113056
rect 121840 103601 121868 113047
rect 121826 103592 121882 103601
rect 121826 103527 121882 103536
rect 121826 103456 121882 103465
rect 121826 103391 121882 103400
rect 121840 93945 121868 103391
rect 121826 93936 121882 93945
rect 121826 93871 121882 93880
rect 121828 81116 121880 81122
rect 121828 81058 121880 81064
rect 121840 80646 121868 81058
rect 121828 80640 121880 80646
rect 121828 80582 121880 80588
rect 121368 73160 121420 73166
rect 121368 73102 121420 73108
rect 121276 73092 121328 73098
rect 121276 73034 121328 73040
rect 121460 72412 121512 72418
rect 121460 72354 121512 72360
rect 120816 70032 120868 70038
rect 120816 69974 120868 69980
rect 120446 55040 120502 55049
rect 120446 54975 120502 54984
rect 120460 54505 120488 54975
rect 120446 54496 120502 54505
rect 120446 54431 120502 54440
rect 120724 3392 120776 3398
rect 120724 3334 120776 3340
rect 119908 3182 120212 3210
rect 118792 3052 118844 3058
rect 118792 2994 118844 3000
rect 118804 480 118832 2994
rect 119908 480 119936 3182
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120736 354 120764 3334
rect 121472 3058 121500 72354
rect 121932 71738 121960 140558
rect 122024 73642 122052 147999
rect 122012 73636 122064 73642
rect 122012 73578 122064 73584
rect 121920 71732 121972 71738
rect 121920 71674 121972 71680
rect 122116 71194 122144 148718
rect 122208 78538 122236 194142
rect 122300 81054 122328 198290
rect 122288 81048 122340 81054
rect 122392 81025 122420 198426
rect 125048 198416 125100 198422
rect 125048 198358 125100 198364
rect 124864 197940 124916 197946
rect 124864 197882 124916 197888
rect 123484 195900 123536 195906
rect 123484 195842 123536 195848
rect 123392 195424 123444 195430
rect 123392 195366 123444 195372
rect 123404 195090 123432 195366
rect 123392 195084 123444 195090
rect 123392 195026 123444 195032
rect 122472 192976 122524 192982
rect 122472 192918 122524 192924
rect 122288 80990 122340 80996
rect 122378 81016 122434 81025
rect 122378 80951 122434 80960
rect 122196 78532 122248 78538
rect 122196 78474 122248 78480
rect 122104 71188 122156 71194
rect 122104 71130 122156 71136
rect 122484 67114 122512 192918
rect 122564 191480 122616 191486
rect 122564 191422 122616 191428
rect 122576 151814 122604 191422
rect 122576 151786 122696 151814
rect 122564 149048 122616 149054
rect 122564 148990 122616 148996
rect 122576 147801 122604 148990
rect 122562 147792 122618 147801
rect 122562 147727 122618 147736
rect 122668 144090 122696 151786
rect 122746 151600 122802 151609
rect 122746 151535 122802 151544
rect 122760 146713 122788 151535
rect 123496 147674 123524 195842
rect 123576 195424 123628 195430
rect 123576 195366 123628 195372
rect 123588 195226 123616 195366
rect 123576 195220 123628 195226
rect 123576 195162 123628 195168
rect 123574 194576 123630 194585
rect 123574 194511 123630 194520
rect 123312 147646 123524 147674
rect 122746 146704 122802 146713
rect 122746 146639 122802 146648
rect 122656 144084 122708 144090
rect 122656 144026 122708 144032
rect 123116 142384 123168 142390
rect 123116 142326 123168 142332
rect 123128 139369 123156 142326
rect 123208 141364 123260 141370
rect 123208 141306 123260 141312
rect 123220 139890 123248 141306
rect 123312 140962 123340 147646
rect 123588 142905 123616 194511
rect 123944 192704 123996 192710
rect 123944 192646 123996 192652
rect 123852 191412 123904 191418
rect 123852 191354 123904 191360
rect 123574 142896 123630 142905
rect 123574 142831 123630 142840
rect 123484 142044 123536 142050
rect 123484 141986 123536 141992
rect 123390 141944 123446 141953
rect 123390 141879 123446 141888
rect 123404 140962 123432 141879
rect 123496 141710 123524 141986
rect 123484 141704 123536 141710
rect 123484 141646 123536 141652
rect 123300 140956 123352 140962
rect 123300 140898 123352 140904
rect 123392 140956 123444 140962
rect 123392 140898 123444 140904
rect 123220 139862 123556 139890
rect 123390 139768 123446 139777
rect 123390 139703 123446 139712
rect 123404 139602 123432 139703
rect 123392 139596 123444 139602
rect 123392 139538 123444 139544
rect 123864 139369 123892 191354
rect 123956 142390 123984 192646
rect 124772 150476 124824 150482
rect 124772 150418 124824 150424
rect 123944 142384 123996 142390
rect 123944 142326 123996 142332
rect 123942 142216 123998 142225
rect 123942 142151 123998 142160
rect 123956 139890 123984 142151
rect 124586 141944 124642 141953
rect 124586 141879 124642 141888
rect 124600 141137 124628 141879
rect 124586 141128 124642 141137
rect 124586 141063 124642 141072
rect 124496 140208 124548 140214
rect 124496 140150 124548 140156
rect 123956 139862 124108 139890
rect 124508 139641 124536 140150
rect 124600 139890 124628 141063
rect 124784 139890 124812 150418
rect 124876 140321 124904 197882
rect 124956 197804 125008 197810
rect 124956 197746 125008 197752
rect 124968 141030 124996 197746
rect 124956 141024 125008 141030
rect 124956 140966 125008 140972
rect 125060 140622 125088 198358
rect 125152 150482 125180 199854
rect 125140 150476 125192 150482
rect 125140 150418 125192 150424
rect 125140 148980 125192 148986
rect 125140 148922 125192 148928
rect 125152 141953 125180 148922
rect 126256 147674 126284 200670
rect 132224 200670 132276 200676
rect 177764 200728 177816 200734
rect 177764 200670 177816 200676
rect 178868 200728 178920 200734
rect 178868 200670 178920 200676
rect 179972 200728 180024 200734
rect 179972 200670 180024 200676
rect 180248 200728 180300 200734
rect 180248 200670 180300 200676
rect 127714 200631 127770 200640
rect 129004 200660 129056 200666
rect 127624 200252 127676 200258
rect 127624 200194 127676 200200
rect 127532 199844 127584 199850
rect 127532 199786 127584 199792
rect 126336 198824 126388 198830
rect 126336 198766 126388 198772
rect 126164 147646 126284 147674
rect 125232 143608 125284 143614
rect 125232 143550 125284 143556
rect 125244 143313 125272 143550
rect 125230 143304 125286 143313
rect 125230 143239 125286 143248
rect 126060 142384 126112 142390
rect 126060 142326 126112 142332
rect 125600 142112 125652 142118
rect 125598 142080 125600 142089
rect 125652 142080 125654 142089
rect 125598 142015 125654 142024
rect 125600 141976 125652 141982
rect 125138 141944 125194 141953
rect 125600 141918 125652 141924
rect 125138 141879 125194 141888
rect 125048 140616 125100 140622
rect 125048 140558 125100 140564
rect 125508 140344 125560 140350
rect 124862 140312 124918 140321
rect 125508 140286 125560 140292
rect 124862 140247 124918 140256
rect 124600 139862 124660 139890
rect 124784 139862 125212 139890
rect 125520 139641 125548 140286
rect 125612 139890 125640 141918
rect 126072 140078 126100 142326
rect 126164 140554 126192 147646
rect 126244 143608 126296 143614
rect 126244 143550 126296 143556
rect 126152 140548 126204 140554
rect 126152 140490 126204 140496
rect 126060 140072 126112 140078
rect 126060 140014 126112 140020
rect 126256 139890 126284 143550
rect 126348 140418 126376 198766
rect 126428 198756 126480 198762
rect 126428 198698 126480 198704
rect 126440 142390 126468 198698
rect 126520 198552 126572 198558
rect 126520 198494 126572 198500
rect 126428 142384 126480 142390
rect 126428 142326 126480 142332
rect 126532 142202 126560 198494
rect 127544 198286 127572 199786
rect 127532 198280 127584 198286
rect 127532 198222 127584 198228
rect 126704 196512 126756 196518
rect 126704 196454 126756 196460
rect 126612 196376 126664 196382
rect 126612 196318 126664 196324
rect 126440 142174 126560 142202
rect 126440 140690 126468 142174
rect 126520 142044 126572 142050
rect 126520 141986 126572 141992
rect 126532 141273 126560 141986
rect 126518 141264 126574 141273
rect 126518 141199 126574 141208
rect 126428 140684 126480 140690
rect 126428 140626 126480 140632
rect 126336 140412 126388 140418
rect 126336 140354 126388 140360
rect 126532 139890 126560 141199
rect 126624 140758 126652 196318
rect 126612 140752 126664 140758
rect 126612 140694 126664 140700
rect 126716 140486 126744 196454
rect 126980 145920 127032 145926
rect 126980 145862 127032 145868
rect 126992 142361 127020 145862
rect 127532 142452 127584 142458
rect 127532 142394 127584 142400
rect 126978 142352 127034 142361
rect 126978 142287 127034 142296
rect 127072 141908 127124 141914
rect 127072 141850 127124 141856
rect 127084 140865 127112 141850
rect 127070 140856 127126 140865
rect 127070 140791 127126 140800
rect 126704 140480 126756 140486
rect 126704 140422 126756 140428
rect 127084 139890 127112 140791
rect 125612 139862 125916 139890
rect 126256 139862 126316 139890
rect 126532 139862 126868 139890
rect 127084 139862 127420 139890
rect 124494 139632 124550 139641
rect 124494 139567 124550 139576
rect 125506 139632 125562 139641
rect 125506 139567 125562 139576
rect 125888 139466 125916 139862
rect 127544 139641 127572 142394
rect 127636 140010 127664 200194
rect 127728 140593 127756 200631
rect 129004 200602 129056 200608
rect 128544 200592 128596 200598
rect 128544 200534 128596 200540
rect 128360 199912 128412 199918
rect 128360 199854 128412 199860
rect 127898 199064 127954 199073
rect 127898 198999 127954 199008
rect 127808 194336 127860 194342
rect 127808 194278 127860 194284
rect 127820 142458 127848 194278
rect 127808 142452 127860 142458
rect 127808 142394 127860 142400
rect 127806 142352 127862 142361
rect 127806 142287 127862 142296
rect 127714 140584 127770 140593
rect 127714 140519 127770 140528
rect 127624 140004 127676 140010
rect 127624 139946 127676 139952
rect 127820 139890 127848 142287
rect 127912 140729 127940 198999
rect 128082 198928 128138 198937
rect 128082 198863 128138 198872
rect 127992 194268 128044 194274
rect 127992 194210 128044 194216
rect 128004 141302 128032 194210
rect 127992 141296 128044 141302
rect 127992 141238 128044 141244
rect 127898 140720 127954 140729
rect 127898 140655 127954 140664
rect 128096 140457 128124 198863
rect 128176 195220 128228 195226
rect 128176 195162 128228 195168
rect 128188 144022 128216 195162
rect 128372 193905 128400 199854
rect 128452 195628 128504 195634
rect 128452 195570 128504 195576
rect 128464 195022 128492 195570
rect 128452 195016 128504 195022
rect 128452 194958 128504 194964
rect 128358 193896 128414 193905
rect 128358 193831 128414 193840
rect 128556 192914 128584 200534
rect 129016 199782 129044 200602
rect 132236 200598 132264 200670
rect 131948 200592 132000 200598
rect 131486 200560 131542 200569
rect 132224 200592 132276 200598
rect 131948 200534 132000 200540
rect 132130 200560 132186 200569
rect 131486 200495 131542 200504
rect 131580 200524 131632 200530
rect 130292 200320 130344 200326
rect 130292 200262 130344 200268
rect 130106 200016 130162 200025
rect 130106 199951 130162 199960
rect 129004 199776 129056 199782
rect 129004 199718 129056 199724
rect 130016 198960 130068 198966
rect 130016 198902 130068 198908
rect 129280 198688 129332 198694
rect 129280 198630 129332 198636
rect 129004 198620 129056 198626
rect 129004 198562 129056 198568
rect 128544 192908 128596 192914
rect 128544 192850 128596 192856
rect 128360 148912 128412 148918
rect 128360 148854 128412 148860
rect 128372 147694 128400 148854
rect 128360 147688 128412 147694
rect 128360 147630 128412 147636
rect 128636 147688 128688 147694
rect 128636 147630 128688 147636
rect 128176 144016 128228 144022
rect 128176 143958 128228 143964
rect 128452 143540 128504 143546
rect 128452 143482 128504 143488
rect 128464 141001 128492 143482
rect 128450 140992 128506 141001
rect 128450 140927 128506 140936
rect 128082 140448 128138 140457
rect 128082 140383 128138 140392
rect 127820 139862 127972 139890
rect 128464 139754 128492 140927
rect 128648 139890 128676 147630
rect 129016 140282 129044 198562
rect 129188 197668 129240 197674
rect 129188 197610 129240 197616
rect 129200 142154 129228 197610
rect 129108 142126 129228 142154
rect 129108 140457 129136 142126
rect 129292 141930 129320 198630
rect 129924 196444 129976 196450
rect 129924 196386 129976 196392
rect 129936 193050 129964 196386
rect 130028 193118 130056 198902
rect 130120 194449 130148 199951
rect 130304 197334 130332 200262
rect 130476 200184 130528 200190
rect 130476 200126 130528 200132
rect 130384 200048 130436 200054
rect 130384 199990 130436 199996
rect 130396 199646 130424 199990
rect 130488 199714 130516 200126
rect 131500 200122 131528 200495
rect 131580 200466 131632 200472
rect 131592 200161 131620 200466
rect 131578 200152 131634 200161
rect 131488 200116 131540 200122
rect 131578 200087 131634 200096
rect 131488 200058 131540 200064
rect 131856 200048 131908 200054
rect 131856 199990 131908 199996
rect 130476 199708 130528 199714
rect 130476 199650 130528 199656
rect 130568 199708 130620 199714
rect 130568 199650 130620 199656
rect 130384 199640 130436 199646
rect 130384 199582 130436 199588
rect 130292 197328 130344 197334
rect 130292 197270 130344 197276
rect 130580 195265 130608 199650
rect 131762 199608 131818 199617
rect 131762 199543 131818 199552
rect 131578 199472 131634 199481
rect 131578 199407 131634 199416
rect 131592 199102 131620 199407
rect 131580 199096 131632 199102
rect 131580 199038 131632 199044
rect 131776 199034 131804 199543
rect 131764 199028 131816 199034
rect 131764 198970 131816 198976
rect 131868 198801 131896 199990
rect 131960 199889 131988 200534
rect 132224 200534 132276 200540
rect 132130 200495 132186 200504
rect 132040 200388 132092 200394
rect 132040 200330 132092 200336
rect 132052 200190 132080 200330
rect 132040 200184 132092 200190
rect 132040 200126 132092 200132
rect 131946 199880 132002 199889
rect 131946 199815 132002 199824
rect 132144 199560 132172 200495
rect 132224 200456 132276 200462
rect 132224 200398 132276 200404
rect 132236 200258 132264 200398
rect 177776 200394 177804 200670
rect 178684 200660 178736 200666
rect 178684 200602 178736 200608
rect 177856 200592 177908 200598
rect 177856 200534 177908 200540
rect 177764 200388 177816 200394
rect 177764 200330 177816 200336
rect 132224 200252 132276 200258
rect 177652 200246 177804 200274
rect 132224 200194 132276 200200
rect 132328 200110 132388 200138
rect 132224 199980 132276 199986
rect 132224 199922 132276 199928
rect 132236 199617 132264 199922
rect 132328 199714 132356 200110
rect 132466 199900 132494 200124
rect 132420 199872 132494 199900
rect 132316 199708 132368 199714
rect 132316 199650 132368 199656
rect 131960 199532 132172 199560
rect 132222 199608 132278 199617
rect 132222 199543 132278 199552
rect 132316 199572 132368 199578
rect 131854 198792 131910 198801
rect 131854 198727 131910 198736
rect 131856 197328 131908 197334
rect 131856 197270 131908 197276
rect 131762 197024 131818 197033
rect 131762 196959 131818 196968
rect 131028 196240 131080 196246
rect 131028 196182 131080 196188
rect 130566 195256 130622 195265
rect 130566 195191 130622 195200
rect 130568 194540 130620 194546
rect 130568 194482 130620 194488
rect 130384 194472 130436 194478
rect 130106 194440 130162 194449
rect 130384 194414 130436 194420
rect 130106 194375 130162 194384
rect 130016 193112 130068 193118
rect 130016 193054 130068 193060
rect 129924 193044 129976 193050
rect 129924 192986 129976 192992
rect 130292 191684 130344 191690
rect 130292 191626 130344 191632
rect 130304 191282 130332 191626
rect 130292 191276 130344 191282
rect 130292 191218 130344 191224
rect 130292 190324 130344 190330
rect 130292 190266 130344 190272
rect 130304 189990 130332 190266
rect 130292 189984 130344 189990
rect 130292 189926 130344 189932
rect 130108 189916 130160 189922
rect 130108 189858 130160 189864
rect 130120 189718 130148 189858
rect 130108 189712 130160 189718
rect 130108 189654 130160 189660
rect 129830 146296 129886 146305
rect 129830 146231 129886 146240
rect 129740 146124 129792 146130
rect 129740 146066 129792 146072
rect 129752 143274 129780 146066
rect 129740 143268 129792 143274
rect 129740 143210 129792 143216
rect 129844 142186 129872 146231
rect 130292 145988 130344 145994
rect 130292 145930 130344 145936
rect 130200 144220 130252 144226
rect 130200 144162 130252 144168
rect 129832 142180 129884 142186
rect 129832 142122 129884 142128
rect 129200 141902 129320 141930
rect 129094 140448 129150 140457
rect 129094 140383 129150 140392
rect 129004 140276 129056 140282
rect 129004 140218 129056 140224
rect 128648 139862 129076 139890
rect 128464 139726 128524 139754
rect 127530 139632 127586 139641
rect 127530 139567 127586 139576
rect 125876 139460 125928 139466
rect 125876 139402 125928 139408
rect 129200 139369 129228 141902
rect 129280 141840 129332 141846
rect 129280 141782 129332 141788
rect 129292 139890 129320 141782
rect 130212 140162 130240 144162
rect 130166 140134 130240 140162
rect 129292 139862 129628 139890
rect 130166 139876 130194 140134
rect 130304 139890 130332 145930
rect 130396 143410 130424 194414
rect 130580 193882 130608 194482
rect 130936 194404 130988 194410
rect 130936 194346 130988 194352
rect 130488 193854 130608 193882
rect 130488 144158 130516 193854
rect 130752 193792 130804 193798
rect 130752 193734 130804 193740
rect 130568 193724 130620 193730
rect 130568 193666 130620 193672
rect 130580 144838 130608 193666
rect 130660 190324 130712 190330
rect 130660 190266 130712 190272
rect 130672 146849 130700 190266
rect 130764 147422 130792 193734
rect 130844 193656 130896 193662
rect 130844 193598 130896 193604
rect 130752 147416 130804 147422
rect 130752 147358 130804 147364
rect 130856 147354 130884 193598
rect 130948 190330 130976 194346
rect 131040 192545 131068 196182
rect 131026 192536 131082 192545
rect 131026 192471 131082 192480
rect 131028 191616 131080 191622
rect 131028 191558 131080 191564
rect 131040 191350 131068 191558
rect 131028 191344 131080 191350
rect 131028 191286 131080 191292
rect 130936 190324 130988 190330
rect 130936 190266 130988 190272
rect 130844 147348 130896 147354
rect 130844 147290 130896 147296
rect 130658 146840 130714 146849
rect 130658 146775 130714 146784
rect 131776 146198 131804 196959
rect 131868 147393 131896 197270
rect 131854 147384 131910 147393
rect 131854 147319 131910 147328
rect 131764 146192 131816 146198
rect 131764 146134 131816 146140
rect 131304 146056 131356 146062
rect 131304 145998 131356 146004
rect 131118 145480 131174 145489
rect 131118 145415 131174 145424
rect 130568 144832 130620 144838
rect 130568 144774 130620 144780
rect 130476 144152 130528 144158
rect 130476 144094 130528 144100
rect 131132 143410 131160 145415
rect 131212 144288 131264 144294
rect 131212 144230 131264 144236
rect 130384 143404 130436 143410
rect 130384 143346 130436 143352
rect 131120 143404 131172 143410
rect 131120 143346 131172 143352
rect 131224 139890 131252 144230
rect 131316 140758 131344 145998
rect 131488 143472 131540 143478
rect 131488 143414 131540 143420
rect 131304 140752 131356 140758
rect 131304 140694 131356 140700
rect 131500 139890 131528 143414
rect 130304 139862 130732 139890
rect 131224 139862 131284 139890
rect 131500 139862 131836 139890
rect 129476 139641 129504 139862
rect 129462 139632 129518 139641
rect 129462 139567 129518 139576
rect 131960 139369 131988 199532
rect 132316 199514 132368 199520
rect 132224 199504 132276 199510
rect 132130 199472 132186 199481
rect 132328 199481 132356 199514
rect 132224 199446 132276 199452
rect 132314 199472 132370 199481
rect 132130 199407 132186 199416
rect 132040 199028 132092 199034
rect 132040 198970 132092 198976
rect 132052 197985 132080 198970
rect 132144 198966 132172 199407
rect 132132 198960 132184 198966
rect 132132 198902 132184 198908
rect 132236 198914 132264 199446
rect 132314 199407 132370 199416
rect 132236 198886 132356 198914
rect 132328 198734 132356 198886
rect 132236 198706 132356 198734
rect 132038 197976 132094 197985
rect 132038 197911 132094 197920
rect 132132 195152 132184 195158
rect 132132 195094 132184 195100
rect 132040 194812 132092 194818
rect 132040 194754 132092 194760
rect 132052 147286 132080 194754
rect 132144 147490 132172 195094
rect 132236 191834 132264 198706
rect 132420 198257 132448 199872
rect 132558 199832 132586 200124
rect 132650 199918 132678 200124
rect 132638 199912 132690 199918
rect 132638 199854 132690 199860
rect 132512 199804 132586 199832
rect 132512 198393 132540 199804
rect 132742 199628 132770 200124
rect 132834 199764 132862 200124
rect 132926 199918 132954 200124
rect 132914 199912 132966 199918
rect 133018 199889 133046 200124
rect 132914 199854 132966 199860
rect 133004 199880 133060 199889
rect 133004 199815 133060 199824
rect 132960 199776 133012 199782
rect 132834 199736 132908 199764
rect 132696 199600 132770 199628
rect 132696 198734 132724 199600
rect 132880 199560 132908 199736
rect 132958 199744 132960 199753
rect 133110 199764 133138 200124
rect 133012 199744 133014 199753
rect 132958 199679 133014 199688
rect 133064 199736 133138 199764
rect 132604 198706 132724 198734
rect 132788 199532 132908 199560
rect 132498 198384 132554 198393
rect 132498 198319 132554 198328
rect 132406 198248 132462 198257
rect 132406 198183 132462 198192
rect 132604 191834 132632 198706
rect 132236 191806 132356 191834
rect 132224 191548 132276 191554
rect 132224 191490 132276 191496
rect 132236 147529 132264 191490
rect 132328 190194 132356 191806
rect 132512 191806 132632 191834
rect 132512 191690 132540 191806
rect 132592 191752 132644 191758
rect 132592 191694 132644 191700
rect 132500 191684 132552 191690
rect 132500 191626 132552 191632
rect 132316 190188 132368 190194
rect 132316 190130 132368 190136
rect 132604 151298 132632 191694
rect 132788 187134 132816 199532
rect 132868 199436 132920 199442
rect 132868 199378 132920 199384
rect 132960 199436 133012 199442
rect 132960 199378 133012 199384
rect 132880 198966 132908 199378
rect 132868 198960 132920 198966
rect 132868 198902 132920 198908
rect 132868 196920 132920 196926
rect 132868 196862 132920 196868
rect 132880 196314 132908 196862
rect 132868 196308 132920 196314
rect 132868 196250 132920 196256
rect 132972 191593 133000 199378
rect 132958 191584 133014 191593
rect 132958 191519 133014 191528
rect 132776 187128 132828 187134
rect 132776 187070 132828 187076
rect 133064 186314 133092 199736
rect 133202 199696 133230 200124
rect 133156 199668 133230 199696
rect 133156 197996 133184 199668
rect 133294 199628 133322 200124
rect 133248 199600 133322 199628
rect 133248 198121 133276 199600
rect 133386 199560 133414 200124
rect 133340 199532 133414 199560
rect 133234 198112 133290 198121
rect 133234 198047 133290 198056
rect 133156 197968 133276 197996
rect 133144 196784 133196 196790
rect 133144 196726 133196 196732
rect 133156 196178 133184 196726
rect 133144 196172 133196 196178
rect 133144 196114 133196 196120
rect 133248 187066 133276 197968
rect 133340 189961 133368 199532
rect 133478 199492 133506 200124
rect 133570 199764 133598 200124
rect 133662 199923 133690 200124
rect 133648 199914 133704 199923
rect 133754 199918 133782 200124
rect 133648 199849 133704 199858
rect 133742 199912 133794 199918
rect 133742 199854 133794 199860
rect 133570 199736 133644 199764
rect 133432 199464 133506 199492
rect 133432 191758 133460 199464
rect 133512 199096 133564 199102
rect 133512 199038 133564 199044
rect 133524 198665 133552 199038
rect 133510 198656 133566 198665
rect 133510 198591 133566 198600
rect 133512 197396 133564 197402
rect 133512 197338 133564 197344
rect 133524 196586 133552 197338
rect 133512 196580 133564 196586
rect 133512 196522 133564 196528
rect 133420 191752 133472 191758
rect 133420 191694 133472 191700
rect 133326 189952 133382 189961
rect 133326 189887 133382 189896
rect 133616 187202 133644 199736
rect 133846 199730 133874 200124
rect 133938 199918 133966 200124
rect 134030 199918 134058 200124
rect 133926 199912 133978 199918
rect 133926 199854 133978 199860
rect 134018 199912 134070 199918
rect 134018 199854 134070 199860
rect 134122 199764 134150 200124
rect 134214 199918 134242 200124
rect 134306 199918 134334 200124
rect 134202 199912 134254 199918
rect 134202 199854 134254 199860
rect 134294 199912 134346 199918
rect 134294 199854 134346 199860
rect 133984 199736 134150 199764
rect 134398 199764 134426 200124
rect 134490 199918 134518 200124
rect 134582 199918 134610 200124
rect 134674 199918 134702 200124
rect 134478 199912 134530 199918
rect 134478 199854 134530 199860
rect 134570 199912 134622 199918
rect 134570 199854 134622 199860
rect 134662 199912 134714 199918
rect 134766 199889 134794 200124
rect 134858 199918 134886 200124
rect 134950 199918 134978 200124
rect 134846 199912 134898 199918
rect 134662 199854 134714 199860
rect 134752 199880 134808 199889
rect 134846 199854 134898 199860
rect 134938 199912 134990 199918
rect 134938 199854 134990 199860
rect 134752 199815 134808 199824
rect 134892 199776 134944 199782
rect 134398 199736 134472 199764
rect 133984 199730 134012 199736
rect 133708 199702 133874 199730
rect 133938 199702 134012 199730
rect 134444 199730 134472 199736
rect 134248 199708 134300 199714
rect 133708 190454 133736 199702
rect 133788 199640 133840 199646
rect 133938 199628 133966 199702
rect 134444 199702 134656 199730
rect 135042 199764 135070 200124
rect 135134 199918 135162 200124
rect 135122 199912 135174 199918
rect 135122 199854 135174 199860
rect 134892 199718 134944 199724
rect 134996 199736 135070 199764
rect 135226 199764 135254 200124
rect 135318 199918 135346 200124
rect 135306 199912 135358 199918
rect 135306 199854 135358 199860
rect 135226 199736 135300 199764
rect 134248 199650 134300 199656
rect 133788 199582 133840 199588
rect 133892 199600 133966 199628
rect 134064 199640 134116 199646
rect 133800 196353 133828 199582
rect 133892 199442 133920 199600
rect 134064 199582 134116 199588
rect 134156 199640 134208 199646
rect 134156 199582 134208 199588
rect 133972 199504 134024 199510
rect 133972 199446 134024 199452
rect 133880 199436 133932 199442
rect 133880 199378 133932 199384
rect 133786 196344 133842 196353
rect 133786 196279 133842 196288
rect 133984 191282 134012 199446
rect 134076 198082 134104 199582
rect 134064 198076 134116 198082
rect 134064 198018 134116 198024
rect 133972 191276 134024 191282
rect 133972 191218 134024 191224
rect 134064 191208 134116 191214
rect 134064 191150 134116 191156
rect 134168 191162 134196 199582
rect 134260 193214 134288 199650
rect 134524 199640 134576 199646
rect 134524 199582 134576 199588
rect 134628 199594 134656 199702
rect 134800 199708 134852 199714
rect 134800 199650 134852 199656
rect 134340 199572 134392 199578
rect 134340 199514 134392 199520
rect 134352 194041 134380 199514
rect 134432 199436 134484 199442
rect 134432 199378 134484 199384
rect 134338 194032 134394 194041
rect 134338 193967 134394 193976
rect 134444 193214 134472 199378
rect 134536 198665 134564 199582
rect 134628 199566 134702 199594
rect 134674 199560 134702 199566
rect 134674 199532 134748 199560
rect 134614 199472 134670 199481
rect 134614 199407 134616 199416
rect 134668 199407 134670 199416
rect 134616 199378 134668 199384
rect 134522 198656 134578 198665
rect 134522 198591 134578 198600
rect 134720 196246 134748 199532
rect 134708 196240 134760 196246
rect 134708 196182 134760 196188
rect 134260 193186 134380 193214
rect 134444 193186 134564 193214
rect 133708 190426 133828 190454
rect 133604 187196 133656 187202
rect 133604 187138 133656 187144
rect 133236 187060 133288 187066
rect 133236 187002 133288 187008
rect 133800 186314 133828 190426
rect 132972 186286 133092 186314
rect 133340 186286 133828 186314
rect 132684 154420 132736 154426
rect 132684 154362 132736 154368
rect 132592 151292 132644 151298
rect 132592 151234 132644 151240
rect 132222 147520 132278 147529
rect 132132 147484 132184 147490
rect 132222 147455 132278 147464
rect 132132 147426 132184 147432
rect 132040 147280 132092 147286
rect 132040 147222 132092 147228
rect 132040 140752 132092 140758
rect 132040 140694 132092 140700
rect 132052 139890 132080 140694
rect 132696 139890 132724 154362
rect 132972 148374 133000 186286
rect 133340 154086 133368 186286
rect 133328 154080 133380 154086
rect 133328 154022 133380 154028
rect 134076 153882 134104 191150
rect 134168 191134 134288 191162
rect 134156 191072 134208 191078
rect 134156 191014 134208 191020
rect 134168 154154 134196 191014
rect 134260 186314 134288 191134
rect 134352 186998 134380 193186
rect 134536 191214 134564 193186
rect 134524 191208 134576 191214
rect 134524 191150 134576 191156
rect 134340 186992 134392 186998
rect 134340 186934 134392 186940
rect 134260 186286 134380 186314
rect 134156 154148 134208 154154
rect 134156 154090 134208 154096
rect 134352 154018 134380 186286
rect 134812 180794 134840 199650
rect 134904 194313 134932 199718
rect 134890 194304 134946 194313
rect 134890 194239 134946 194248
rect 134996 187270 135024 199736
rect 135168 199640 135220 199646
rect 135168 199582 135220 199588
rect 135076 199300 135128 199306
rect 135076 199242 135128 199248
rect 135088 199102 135116 199242
rect 135076 199096 135128 199102
rect 135076 199038 135128 199044
rect 135180 191078 135208 199582
rect 135272 199578 135300 199736
rect 135410 199696 135438 200124
rect 135502 199918 135530 200124
rect 135490 199912 135542 199918
rect 135594 199889 135622 200124
rect 135686 199918 135714 200124
rect 135674 199912 135726 199918
rect 135490 199854 135542 199860
rect 135580 199880 135636 199889
rect 135674 199854 135726 199860
rect 135580 199815 135636 199824
rect 135778 199764 135806 200124
rect 135732 199736 135806 199764
rect 135732 199696 135760 199736
rect 135410 199668 135576 199696
rect 135260 199572 135312 199578
rect 135260 199514 135312 199520
rect 135352 199572 135404 199578
rect 135352 199514 135404 199520
rect 135444 199572 135496 199578
rect 135444 199514 135496 199520
rect 135258 199472 135314 199481
rect 135258 199407 135314 199416
rect 135272 199209 135300 199407
rect 135258 199200 135314 199209
rect 135258 199135 135314 199144
rect 135258 196208 135314 196217
rect 135258 196143 135314 196152
rect 135272 191622 135300 196143
rect 135364 195945 135392 199514
rect 135350 195936 135406 195945
rect 135350 195871 135406 195880
rect 135456 195673 135484 199514
rect 135548 196081 135576 199668
rect 135640 199668 135760 199696
rect 135534 196072 135590 196081
rect 135534 196007 135590 196016
rect 135442 195664 135498 195673
rect 135442 195599 135498 195608
rect 135640 191834 135668 199668
rect 135870 199628 135898 200124
rect 135962 199696 135990 200124
rect 136054 199918 136082 200124
rect 136042 199912 136094 199918
rect 136042 199854 136094 199860
rect 136146 199764 136174 200124
rect 136238 199918 136266 200124
rect 136330 199918 136358 200124
rect 136422 199923 136450 200124
rect 136226 199912 136278 199918
rect 136226 199854 136278 199860
rect 136318 199912 136370 199918
rect 136318 199854 136370 199860
rect 136408 199914 136464 199923
rect 136408 199849 136464 199858
rect 136514 199764 136542 200124
rect 136146 199736 136220 199764
rect 135962 199668 136036 199696
rect 135870 199600 135944 199628
rect 135720 199572 135772 199578
rect 135772 199532 135852 199560
rect 135720 199514 135772 199520
rect 135720 199300 135772 199306
rect 135720 199242 135772 199248
rect 135732 199102 135760 199242
rect 135720 199096 135772 199102
rect 135720 199038 135772 199044
rect 135640 191806 135760 191834
rect 135260 191616 135312 191622
rect 135260 191558 135312 191564
rect 135732 191298 135760 191806
rect 135640 191270 135760 191298
rect 135168 191072 135220 191078
rect 135168 191014 135220 191020
rect 135536 191072 135588 191078
rect 135536 191014 135588 191020
rect 134984 187264 135036 187270
rect 134984 187206 135036 187212
rect 134444 180766 134840 180794
rect 134340 154012 134392 154018
rect 134340 153954 134392 153960
rect 134444 153950 134472 180766
rect 134432 153944 134484 153950
rect 134432 153886 134484 153892
rect 134064 153876 134116 153882
rect 134064 153818 134116 153824
rect 135548 151162 135576 191014
rect 135640 190126 135668 191270
rect 135720 191208 135772 191214
rect 135720 191150 135772 191156
rect 135628 190120 135680 190126
rect 135628 190062 135680 190068
rect 135536 151156 135588 151162
rect 135536 151098 135588 151104
rect 135732 148889 135760 191150
rect 135824 149802 135852 199532
rect 135916 199209 135944 199600
rect 136008 199594 136036 199668
rect 136008 199566 136128 199594
rect 135996 199504 136048 199510
rect 135996 199446 136048 199452
rect 135902 199200 135958 199209
rect 135902 199135 135958 199144
rect 135904 199096 135956 199102
rect 135904 199038 135956 199044
rect 135916 198966 135944 199038
rect 135904 198960 135956 198966
rect 135904 198902 135956 198908
rect 136008 198218 136036 199446
rect 135996 198212 136048 198218
rect 135996 198154 136048 198160
rect 136100 195974 136128 199566
rect 135916 195946 136128 195974
rect 135812 149796 135864 149802
rect 135812 149738 135864 149744
rect 135916 149734 135944 195946
rect 136192 191834 136220 199736
rect 136468 199736 136542 199764
rect 136272 199640 136324 199646
rect 136272 199582 136324 199588
rect 136100 191806 136220 191834
rect 136100 189786 136128 191806
rect 136284 191214 136312 199582
rect 136362 199200 136418 199209
rect 136362 199135 136418 199144
rect 136272 191208 136324 191214
rect 136272 191150 136324 191156
rect 136376 190262 136404 199135
rect 136468 191078 136496 199736
rect 136606 199696 136634 200124
rect 136698 199918 136726 200124
rect 136686 199912 136738 199918
rect 136686 199854 136738 199860
rect 136790 199764 136818 200124
rect 136882 199923 136910 200124
rect 136868 199914 136924 199923
rect 136868 199849 136924 199858
rect 136974 199764 137002 200124
rect 137066 199918 137094 200124
rect 137158 199923 137186 200124
rect 137054 199912 137106 199918
rect 137054 199854 137106 199860
rect 137144 199914 137200 199923
rect 137250 199918 137278 200124
rect 137342 199918 137370 200124
rect 137144 199849 137200 199858
rect 137238 199912 137290 199918
rect 137238 199854 137290 199860
rect 137330 199912 137382 199918
rect 137330 199854 137382 199860
rect 136790 199736 136864 199764
rect 136560 199668 136634 199696
rect 136560 196897 136588 199668
rect 136732 199640 136784 199646
rect 136732 199582 136784 199588
rect 136640 199572 136692 199578
rect 136640 199514 136692 199520
rect 136546 196888 136602 196897
rect 136546 196823 136602 196832
rect 136652 196722 136680 199514
rect 136744 197169 136772 199582
rect 136730 197160 136786 197169
rect 136730 197095 136786 197104
rect 136836 196897 136864 199736
rect 136928 199736 137002 199764
rect 137284 199776 137336 199782
rect 136822 196888 136878 196897
rect 136822 196823 136878 196832
rect 136640 196716 136692 196722
rect 136640 196658 136692 196664
rect 136456 191072 136508 191078
rect 136456 191014 136508 191020
rect 136364 190256 136416 190262
rect 136364 190198 136416 190204
rect 136928 189854 136956 199736
rect 137434 199764 137462 200124
rect 137526 199923 137554 200124
rect 137512 199914 137568 199923
rect 137618 199918 137646 200124
rect 137710 199918 137738 200124
rect 137802 199918 137830 200124
rect 137894 199918 137922 200124
rect 137512 199849 137568 199858
rect 137606 199912 137658 199918
rect 137606 199854 137658 199860
rect 137698 199912 137750 199918
rect 137698 199854 137750 199860
rect 137790 199912 137842 199918
rect 137790 199854 137842 199860
rect 137882 199912 137934 199918
rect 137882 199854 137934 199860
rect 137284 199718 137336 199724
rect 137388 199736 137462 199764
rect 137652 199776 137704 199782
rect 137100 199708 137152 199714
rect 137100 199650 137152 199656
rect 137008 199436 137060 199442
rect 137008 199378 137060 199384
rect 137020 198966 137048 199378
rect 137008 198960 137060 198966
rect 137008 198902 137060 198908
rect 137112 191834 137140 199650
rect 137192 199436 137244 199442
rect 137192 199378 137244 199384
rect 137204 198801 137232 199378
rect 137190 198792 137246 198801
rect 137190 198727 137246 198736
rect 137296 197305 137324 199718
rect 137282 197296 137338 197305
rect 137282 197231 137338 197240
rect 137388 197198 137416 199736
rect 137652 199718 137704 199724
rect 137744 199776 137796 199782
rect 137986 199764 138014 200124
rect 138078 199918 138106 200124
rect 138170 199918 138198 200124
rect 138262 199918 138290 200124
rect 138354 199923 138382 200124
rect 138066 199912 138118 199918
rect 138066 199854 138118 199860
rect 138158 199912 138210 199918
rect 138158 199854 138210 199860
rect 138250 199912 138302 199918
rect 138250 199854 138302 199860
rect 138340 199914 138396 199923
rect 138446 199918 138474 200124
rect 138538 199923 138566 200124
rect 138340 199849 138396 199858
rect 138434 199912 138486 199918
rect 138434 199854 138486 199860
rect 138524 199914 138580 199923
rect 138630 199918 138658 200124
rect 138524 199849 138580 199858
rect 138618 199912 138670 199918
rect 138618 199854 138670 199860
rect 137744 199718 137796 199724
rect 137940 199736 138014 199764
rect 138112 199776 138164 199782
rect 137468 199640 137520 199646
rect 137468 199582 137520 199588
rect 137560 199640 137612 199646
rect 137560 199582 137612 199588
rect 137480 197198 137508 199582
rect 137376 197192 137428 197198
rect 137376 197134 137428 197140
rect 137468 197192 137520 197198
rect 137468 197134 137520 197140
rect 137284 196920 137336 196926
rect 137284 196862 137336 196868
rect 137466 196888 137522 196897
rect 137112 191806 137232 191834
rect 137100 191208 137152 191214
rect 137100 191150 137152 191156
rect 136916 189848 136968 189854
rect 136916 189790 136968 189796
rect 136088 189780 136140 189786
rect 136088 189722 136140 189728
rect 135904 149728 135956 149734
rect 135904 149670 135956 149676
rect 136178 149016 136234 149025
rect 136178 148951 136234 148960
rect 135718 148880 135774 148889
rect 135718 148815 135774 148824
rect 132960 148368 133012 148374
rect 132960 148310 133012 148316
rect 136192 147694 136220 148951
rect 136180 147688 136232 147694
rect 136180 147630 136232 147636
rect 137112 147257 137140 191150
rect 137204 151366 137232 191806
rect 137296 189922 137324 196862
rect 137466 196823 137522 196832
rect 137284 189916 137336 189922
rect 137284 189858 137336 189864
rect 137480 189718 137508 196823
rect 137572 191214 137600 199582
rect 137664 195498 137692 199718
rect 137652 195492 137704 195498
rect 137652 195434 137704 195440
rect 137560 191208 137612 191214
rect 137560 191150 137612 191156
rect 137756 189990 137784 199718
rect 137836 199708 137888 199714
rect 137836 199650 137888 199656
rect 137744 189984 137796 189990
rect 137744 189926 137796 189932
rect 137468 189712 137520 189718
rect 137468 189654 137520 189660
rect 137848 180794 137876 199650
rect 137940 195090 137968 199736
rect 138112 199718 138164 199724
rect 138204 199776 138256 199782
rect 138204 199718 138256 199724
rect 138388 199776 138440 199782
rect 138722 199764 138750 200124
rect 138814 199923 138842 200124
rect 138800 199914 138856 199923
rect 138800 199849 138856 199858
rect 138906 199764 138934 200124
rect 138998 199918 139026 200124
rect 138986 199912 139038 199918
rect 138986 199854 139038 199860
rect 139090 199764 139118 200124
rect 138388 199718 138440 199724
rect 138676 199736 138750 199764
rect 138860 199736 138934 199764
rect 139044 199736 139118 199764
rect 138020 199504 138072 199510
rect 138020 199446 138072 199452
rect 137928 195084 137980 195090
rect 137928 195026 137980 195032
rect 138032 192574 138060 199446
rect 138124 198529 138152 199718
rect 138110 198520 138166 198529
rect 138110 198455 138166 198464
rect 138112 197192 138164 197198
rect 138112 197134 138164 197140
rect 138020 192568 138072 192574
rect 138020 192510 138072 192516
rect 138124 191834 138152 197134
rect 138216 196704 138244 199718
rect 138294 199200 138350 199209
rect 138294 199135 138350 199144
rect 138308 199034 138336 199135
rect 138296 199028 138348 199034
rect 138296 198970 138348 198976
rect 138400 196926 138428 199718
rect 138572 199708 138624 199714
rect 138572 199650 138624 199656
rect 138388 196920 138440 196926
rect 138388 196862 138440 196868
rect 138584 196840 138612 199650
rect 138676 196897 138704 199736
rect 138756 199504 138808 199510
rect 138756 199446 138808 199452
rect 138492 196812 138612 196840
rect 138662 196888 138718 196897
rect 138662 196823 138718 196832
rect 138216 196676 138428 196704
rect 138296 195492 138348 195498
rect 138296 195434 138348 195440
rect 138124 191806 138244 191834
rect 137480 180766 137876 180794
rect 137480 151473 137508 180766
rect 138216 151502 138244 191806
rect 138204 151496 138256 151502
rect 137466 151464 137522 151473
rect 138204 151438 138256 151444
rect 137466 151399 137522 151408
rect 137192 151360 137244 151366
rect 137192 151302 137244 151308
rect 138308 151094 138336 195434
rect 138296 151088 138348 151094
rect 138296 151030 138348 151036
rect 137098 147248 137154 147257
rect 137098 147183 137154 147192
rect 135810 146160 135866 146169
rect 135810 146095 135866 146104
rect 133880 144900 133932 144906
rect 133880 144842 133932 144848
rect 133144 143200 133196 143206
rect 133144 143142 133196 143148
rect 133156 139890 133184 143142
rect 133892 139890 133920 144842
rect 135444 144696 135496 144702
rect 135444 144638 135496 144644
rect 134800 143336 134852 143342
rect 134800 143278 134852 143284
rect 134248 142180 134300 142186
rect 134248 142122 134300 142128
rect 134260 139890 134288 142122
rect 134812 139890 134840 143278
rect 135456 139890 135484 144638
rect 135824 139890 135852 146095
rect 138112 144764 138164 144770
rect 138112 144706 138164 144712
rect 137560 143404 137612 143410
rect 137560 143346 137612 143352
rect 137008 143268 137060 143274
rect 137008 143210 137060 143216
rect 136640 141704 136692 141710
rect 136640 141646 136692 141652
rect 136652 139890 136680 141646
rect 137020 139890 137048 143210
rect 137572 139890 137600 143346
rect 138124 139890 138152 144706
rect 138400 140350 138428 196676
rect 138492 196042 138520 196812
rect 138572 196716 138624 196722
rect 138572 196658 138624 196664
rect 138480 196036 138532 196042
rect 138480 195978 138532 195984
rect 138480 193044 138532 193050
rect 138480 192986 138532 192992
rect 138492 151745 138520 192986
rect 138584 187241 138612 196658
rect 138664 196036 138716 196042
rect 138664 195978 138716 195984
rect 138676 190398 138704 195978
rect 138768 194177 138796 199446
rect 138860 196722 138888 199736
rect 138940 199640 138992 199646
rect 138940 199582 138992 199588
rect 138848 196716 138900 196722
rect 138848 196658 138900 196664
rect 138952 195974 138980 199582
rect 139044 199510 139072 199736
rect 139182 199696 139210 200124
rect 139274 199923 139302 200124
rect 139260 199914 139316 199923
rect 139366 199918 139394 200124
rect 139458 199918 139486 200124
rect 139550 199923 139578 200124
rect 139260 199849 139316 199858
rect 139354 199912 139406 199918
rect 139354 199854 139406 199860
rect 139446 199912 139498 199918
rect 139446 199854 139498 199860
rect 139536 199914 139592 199923
rect 139642 199918 139670 200124
rect 139734 199918 139762 200124
rect 139536 199849 139592 199858
rect 139630 199912 139682 199918
rect 139630 199854 139682 199860
rect 139722 199912 139774 199918
rect 139722 199854 139774 199860
rect 139826 199850 139854 200124
rect 139918 199923 139946 200124
rect 139904 199914 139960 199923
rect 139814 199844 139866 199850
rect 139904 199849 139960 199858
rect 140010 199850 140038 200124
rect 140102 199923 140130 200124
rect 140088 199914 140144 199923
rect 139814 199786 139866 199792
rect 139998 199844 140050 199850
rect 140088 199849 140144 199858
rect 139998 199786 140050 199792
rect 139398 199744 139454 199753
rect 139182 199668 139256 199696
rect 140042 199744 140098 199753
rect 139398 199679 139454 199688
rect 139492 199708 139544 199714
rect 139032 199504 139084 199510
rect 139032 199446 139084 199452
rect 139124 199504 139176 199510
rect 139124 199446 139176 199452
rect 138952 195946 139072 195974
rect 139044 195498 139072 195946
rect 139032 195492 139084 195498
rect 139032 195434 139084 195440
rect 138754 194168 138810 194177
rect 138754 194103 138810 194112
rect 139136 194070 139164 199446
rect 139228 194818 139256 199668
rect 139412 199424 139440 199679
rect 139492 199650 139544 199656
rect 139860 199708 139912 199714
rect 139860 199650 139912 199656
rect 139952 199708 140004 199714
rect 140194 199714 140222 200124
rect 140286 199918 140314 200124
rect 140274 199912 140326 199918
rect 140274 199854 140326 199860
rect 140042 199679 140098 199688
rect 140182 199708 140234 199714
rect 139952 199650 140004 199656
rect 139320 199396 139440 199424
rect 139216 194812 139268 194818
rect 139216 194754 139268 194760
rect 139124 194064 139176 194070
rect 139124 194006 139176 194012
rect 139320 193050 139348 199396
rect 139398 199200 139454 199209
rect 139398 199135 139454 199144
rect 139412 198966 139440 199135
rect 139400 198960 139452 198966
rect 139400 198902 139452 198908
rect 139504 197334 139532 199650
rect 139768 199572 139820 199578
rect 139768 199514 139820 199520
rect 139492 197328 139544 197334
rect 139492 197270 139544 197276
rect 139584 197328 139636 197334
rect 139780 197305 139808 199514
rect 139584 197270 139636 197276
rect 139766 197296 139822 197305
rect 139308 193044 139360 193050
rect 139308 192986 139360 192992
rect 139596 191554 139624 197270
rect 139766 197231 139822 197240
rect 139768 197192 139820 197198
rect 139768 197134 139820 197140
rect 139676 196920 139728 196926
rect 139676 196862 139728 196868
rect 139584 191548 139636 191554
rect 139584 191490 139636 191496
rect 138664 190392 138716 190398
rect 138664 190334 138716 190340
rect 138570 187232 138626 187241
rect 138570 187167 138626 187176
rect 138478 151736 138534 151745
rect 138478 151671 138534 151680
rect 139688 151230 139716 196862
rect 139676 151224 139728 151230
rect 139676 151166 139728 151172
rect 139780 146962 139808 197134
rect 139872 196874 139900 199650
rect 139964 197334 139992 199650
rect 139952 197328 140004 197334
rect 139952 197270 140004 197276
rect 140056 197198 140084 199679
rect 140378 199696 140406 200124
rect 140470 199918 140498 200124
rect 140562 199918 140590 200124
rect 140458 199912 140510 199918
rect 140458 199854 140510 199860
rect 140550 199912 140602 199918
rect 140654 199889 140682 200124
rect 140550 199854 140602 199860
rect 140640 199880 140696 199889
rect 140640 199815 140696 199824
rect 140746 199764 140774 200124
rect 140838 199918 140866 200124
rect 140930 199923 140958 200124
rect 140826 199912 140878 199918
rect 140826 199854 140878 199860
rect 140916 199914 140972 199923
rect 141022 199918 141050 200124
rect 141114 199918 141142 200124
rect 141206 199923 141234 200124
rect 140916 199849 140972 199858
rect 141010 199912 141062 199918
rect 141010 199854 141062 199860
rect 141102 199912 141154 199918
rect 141102 199854 141154 199860
rect 141192 199914 141248 199923
rect 141298 199918 141326 200124
rect 141390 199918 141418 200124
rect 141192 199849 141248 199858
rect 141286 199912 141338 199918
rect 141286 199854 141338 199860
rect 141378 199912 141430 199918
rect 141378 199854 141430 199860
rect 141482 199782 141510 200124
rect 141574 199923 141602 200124
rect 141560 199914 141616 199923
rect 141560 199849 141616 199858
rect 140182 199650 140234 199656
rect 140332 199668 140406 199696
rect 140502 199744 140558 199753
rect 140502 199679 140558 199688
rect 140700 199736 140774 199764
rect 140872 199776 140924 199782
rect 140136 199572 140188 199578
rect 140136 199514 140188 199520
rect 140148 198734 140176 199514
rect 140148 198706 140268 198734
rect 140044 197192 140096 197198
rect 140044 197134 140096 197140
rect 139872 196846 140084 196874
rect 139860 196784 139912 196790
rect 139860 196726 139912 196732
rect 139688 146934 139808 146962
rect 138662 144664 138718 144673
rect 138662 144599 138718 144608
rect 138388 140344 138440 140350
rect 138388 140286 138440 140292
rect 138676 139890 138704 144599
rect 139400 141636 139452 141642
rect 139400 141578 139452 141584
rect 139412 139890 139440 141578
rect 139688 140214 139716 146934
rect 139768 143132 139820 143138
rect 139768 143074 139820 143080
rect 139676 140208 139728 140214
rect 139676 140150 139728 140156
rect 139780 139890 139808 143074
rect 139872 140321 139900 196726
rect 139952 196716 140004 196722
rect 139952 196658 140004 196664
rect 139964 187105 139992 196658
rect 139950 187096 140006 187105
rect 139950 187031 140006 187040
rect 140056 141681 140084 196846
rect 140240 195809 140268 198706
rect 140332 196790 140360 199668
rect 140412 199572 140464 199578
rect 140412 199514 140464 199520
rect 140320 196784 140372 196790
rect 140320 196726 140372 196732
rect 140424 196722 140452 199514
rect 140516 196926 140544 199679
rect 140596 199640 140648 199646
rect 140596 199582 140648 199588
rect 140504 196920 140556 196926
rect 140504 196862 140556 196868
rect 140412 196716 140464 196722
rect 140412 196658 140464 196664
rect 140608 196450 140636 199582
rect 140596 196444 140648 196450
rect 140596 196386 140648 196392
rect 140700 195974 140728 199736
rect 141148 199776 141200 199782
rect 140872 199718 140924 199724
rect 140962 199744 141018 199753
rect 140780 199640 140832 199646
rect 140780 199582 140832 199588
rect 140792 198014 140820 199582
rect 140884 198257 140912 199718
rect 141148 199718 141200 199724
rect 141470 199776 141522 199782
rect 141666 199764 141694 200124
rect 141758 199918 141786 200124
rect 141850 199918 141878 200124
rect 141746 199912 141798 199918
rect 141746 199854 141798 199860
rect 141838 199912 141890 199918
rect 141838 199854 141890 199860
rect 141942 199764 141970 200124
rect 142034 199918 142062 200124
rect 142022 199912 142074 199918
rect 142022 199854 142074 199860
rect 141666 199736 141740 199764
rect 141470 199718 141522 199724
rect 140962 199679 141018 199688
rect 140976 198734 141004 199679
rect 141160 199481 141188 199718
rect 141516 199640 141568 199646
rect 141516 199582 141568 199588
rect 141240 199572 141292 199578
rect 141240 199514 141292 199520
rect 141146 199472 141202 199481
rect 141146 199407 141202 199416
rect 141252 198801 141280 199514
rect 141332 199504 141384 199510
rect 141332 199446 141384 199452
rect 141424 199504 141476 199510
rect 141424 199446 141476 199452
rect 141238 198792 141294 198801
rect 140976 198706 141188 198734
rect 141238 198727 141294 198736
rect 140870 198248 140926 198257
rect 140870 198183 140926 198192
rect 141056 198212 141108 198218
rect 141056 198154 141108 198160
rect 140962 198112 141018 198121
rect 140962 198047 141018 198056
rect 140780 198008 140832 198014
rect 140780 197950 140832 197956
rect 140872 196648 140924 196654
rect 140872 196590 140924 196596
rect 140700 195946 140820 195974
rect 140226 195800 140282 195809
rect 140226 195735 140282 195744
rect 140792 194138 140820 195946
rect 140780 194132 140832 194138
rect 140780 194074 140832 194080
rect 140884 149841 140912 196590
rect 140976 151434 141004 198047
rect 141068 151609 141096 198154
rect 141160 151706 141188 198706
rect 141344 197402 141372 199446
rect 141436 198966 141464 199446
rect 141424 198960 141476 198966
rect 141424 198902 141476 198908
rect 141422 198792 141478 198801
rect 141422 198727 141478 198736
rect 141332 197396 141384 197402
rect 141332 197338 141384 197344
rect 141240 197328 141292 197334
rect 141240 197270 141292 197276
rect 141252 191486 141280 197270
rect 141436 196722 141464 198727
rect 141528 198218 141556 199582
rect 141606 199472 141662 199481
rect 141606 199407 141662 199416
rect 141516 198212 141568 198218
rect 141516 198154 141568 198160
rect 141424 196716 141476 196722
rect 141424 196658 141476 196664
rect 141620 196110 141648 199407
rect 141608 196104 141660 196110
rect 141608 196046 141660 196052
rect 141712 193594 141740 199736
rect 141896 199736 141970 199764
rect 141896 199696 141924 199736
rect 141804 199668 141924 199696
rect 142022 199708 142074 199714
rect 141804 199617 141832 199668
rect 142022 199650 142074 199656
rect 141790 199608 141846 199617
rect 142034 199560 142062 199650
rect 142126 199594 142154 200124
rect 142218 199696 142246 200124
rect 142310 199764 142338 200124
rect 142402 199918 142430 200124
rect 142390 199912 142442 199918
rect 142390 199854 142442 199860
rect 142310 199736 142384 199764
rect 142218 199668 142292 199696
rect 142126 199566 142200 199594
rect 141790 199543 141846 199552
rect 141942 199532 142062 199560
rect 141792 199504 141844 199510
rect 141942 199492 141970 199532
rect 141942 199464 142016 199492
rect 141792 199446 141844 199452
rect 141804 196654 141832 199446
rect 141882 198792 141938 198801
rect 141882 198727 141938 198736
rect 141896 197334 141924 198727
rect 141884 197328 141936 197334
rect 141884 197270 141936 197276
rect 141884 197192 141936 197198
rect 141884 197134 141936 197140
rect 141792 196648 141844 196654
rect 141792 196590 141844 196596
rect 141896 195537 141924 197134
rect 141882 195528 141938 195537
rect 141882 195463 141938 195472
rect 141700 193588 141752 193594
rect 141700 193530 141752 193536
rect 141240 191480 141292 191486
rect 141240 191422 141292 191428
rect 141988 180794 142016 199464
rect 142172 198898 142200 199566
rect 142160 198892 142212 198898
rect 142160 198834 142212 198840
rect 142066 198792 142122 198801
rect 142066 198727 142122 198736
rect 142080 197062 142108 198727
rect 142068 197056 142120 197062
rect 142068 196998 142120 197004
rect 142264 194313 142292 199668
rect 142356 197198 142384 199736
rect 142494 199696 142522 200124
rect 142448 199668 142522 199696
rect 142344 197192 142396 197198
rect 142344 197134 142396 197140
rect 142448 196058 142476 199668
rect 142586 199628 142614 200124
rect 142678 199923 142706 200124
rect 142664 199914 142720 199923
rect 142664 199849 142720 199858
rect 142770 199730 142798 200124
rect 142540 199600 142614 199628
rect 142724 199702 142798 199730
rect 142540 197878 142568 199600
rect 142618 199472 142674 199481
rect 142618 199407 142674 199416
rect 142632 198966 142660 199407
rect 142620 198960 142672 198966
rect 142620 198902 142672 198908
rect 142528 197872 142580 197878
rect 142528 197814 142580 197820
rect 142448 196030 142568 196058
rect 142434 195936 142490 195945
rect 142434 195871 142490 195880
rect 142250 194304 142306 194313
rect 142250 194239 142306 194248
rect 141804 180766 142016 180794
rect 141240 154284 141292 154290
rect 141240 154226 141292 154232
rect 141148 151700 141200 151706
rect 141148 151642 141200 151648
rect 141054 151600 141110 151609
rect 141054 151535 141110 151544
rect 140964 151428 141016 151434
rect 140964 151370 141016 151376
rect 140870 149832 140926 149841
rect 140870 149767 140926 149776
rect 140320 141772 140372 141778
rect 140320 141714 140372 141720
rect 140042 141672 140098 141681
rect 140042 141607 140098 141616
rect 139858 140312 139914 140321
rect 139858 140247 139914 140256
rect 140332 139890 140360 141714
rect 141252 140162 141280 154226
rect 141804 149870 141832 180766
rect 142448 151570 142476 195871
rect 142436 151564 142488 151570
rect 142436 151506 142488 151512
rect 141792 149864 141844 149870
rect 141792 149806 141844 149812
rect 142540 148850 142568 196030
rect 142528 148844 142580 148850
rect 142528 148786 142580 148792
rect 142724 148714 142752 199702
rect 142862 199594 142890 200124
rect 142954 199850 142982 200124
rect 142942 199844 142994 199850
rect 142942 199786 142994 199792
rect 143046 199753 143074 200124
rect 143138 199923 143166 200124
rect 143124 199914 143180 199923
rect 143230 199918 143258 200124
rect 143124 199849 143180 199858
rect 143218 199912 143270 199918
rect 143218 199854 143270 199860
rect 143322 199764 143350 200124
rect 143414 199923 143442 200124
rect 143400 199914 143456 199923
rect 143400 199849 143456 199858
rect 143032 199744 143088 199753
rect 143276 199736 143350 199764
rect 143276 199696 143304 199736
rect 143506 199696 143534 200124
rect 143598 199714 143626 200124
rect 143690 199730 143718 200124
rect 143782 199850 143810 200124
rect 143874 199850 143902 200124
rect 143966 199850 143994 200124
rect 144058 199923 144086 200124
rect 144044 199914 144100 199923
rect 143770 199844 143822 199850
rect 143770 199786 143822 199792
rect 143862 199844 143914 199850
rect 143862 199786 143914 199792
rect 143954 199844 144006 199850
rect 144044 199849 144100 199858
rect 144150 199850 144178 200124
rect 144242 199923 144270 200124
rect 144228 199914 144284 199923
rect 143954 199786 144006 199792
rect 144138 199844 144190 199850
rect 144228 199849 144284 199858
rect 144138 199786 144190 199792
rect 144334 199730 144362 200124
rect 144426 199764 144454 200124
rect 144518 199918 144546 200124
rect 144610 199918 144638 200124
rect 144702 199918 144730 200124
rect 144794 199918 144822 200124
rect 144506 199912 144558 199918
rect 144506 199854 144558 199860
rect 144598 199912 144650 199918
rect 144598 199854 144650 199860
rect 144690 199912 144742 199918
rect 144690 199854 144742 199860
rect 144782 199912 144834 199918
rect 144782 199854 144834 199860
rect 144886 199764 144914 200124
rect 144978 199918 145006 200124
rect 145070 199918 145098 200124
rect 145162 199923 145190 200124
rect 144966 199912 145018 199918
rect 144966 199854 145018 199860
rect 145058 199912 145110 199918
rect 145058 199854 145110 199860
rect 145148 199914 145204 199923
rect 145148 199849 145204 199858
rect 145012 199776 145064 199782
rect 144426 199736 144500 199764
rect 144886 199736 144960 199764
rect 143032 199679 143088 199688
rect 143184 199668 143304 199696
rect 143460 199668 143534 199696
rect 143586 199708 143638 199714
rect 143184 199628 143212 199668
rect 142816 199566 142890 199594
rect 143092 199600 143212 199628
rect 143354 199608 143410 199617
rect 142988 199572 143040 199578
rect 142816 195430 142844 199566
rect 142988 199514 143040 199520
rect 143000 199424 143028 199514
rect 143092 199481 143120 199600
rect 143264 199572 143316 199578
rect 143354 199543 143410 199552
rect 143264 199514 143316 199520
rect 142908 199396 143028 199424
rect 143078 199472 143134 199481
rect 143078 199407 143134 199416
rect 142804 195424 142856 195430
rect 142804 195366 142856 195372
rect 142908 194954 142936 199396
rect 142988 198960 143040 198966
rect 142988 198902 143040 198908
rect 143000 196654 143028 198902
rect 143172 198892 143224 198898
rect 143172 198834 143224 198840
rect 143078 198792 143134 198801
rect 143078 198727 143134 198736
rect 142988 196648 143040 196654
rect 142988 196590 143040 196596
rect 142896 194948 142948 194954
rect 142896 194890 142948 194896
rect 143092 192642 143120 198727
rect 143184 196897 143212 198834
rect 143276 196994 143304 199514
rect 143368 198150 143396 199543
rect 143356 198144 143408 198150
rect 143356 198086 143408 198092
rect 143460 197010 143488 199668
rect 143690 199702 143764 199730
rect 143586 199650 143638 199656
rect 143540 199572 143592 199578
rect 143540 199514 143592 199520
rect 143632 199572 143684 199578
rect 143632 199514 143684 199520
rect 143264 196988 143316 196994
rect 143264 196930 143316 196936
rect 143368 196982 143488 197010
rect 143170 196888 143226 196897
rect 143170 196823 143226 196832
rect 143172 196648 143224 196654
rect 143172 196590 143224 196596
rect 143080 192636 143132 192642
rect 143080 192578 143132 192584
rect 143184 191834 143212 196590
rect 143368 195294 143396 196982
rect 143448 196920 143500 196926
rect 143448 196862 143500 196868
rect 143356 195288 143408 195294
rect 143356 195230 143408 195236
rect 143000 191806 143212 191834
rect 143000 151638 143028 191806
rect 143460 191146 143488 196862
rect 143552 194206 143580 199514
rect 143644 197674 143672 199514
rect 143632 197668 143684 197674
rect 143632 197610 143684 197616
rect 143736 196840 143764 199702
rect 143908 199708 143960 199714
rect 143908 199650 143960 199656
rect 144092 199708 144144 199714
rect 144092 199650 144144 199656
rect 144288 199702 144362 199730
rect 143816 199504 143868 199510
rect 143814 199472 143816 199481
rect 143868 199472 143870 199481
rect 143814 199407 143870 199416
rect 143920 199356 143948 199650
rect 143998 199608 144054 199617
rect 143998 199543 144054 199552
rect 143828 199328 143948 199356
rect 143828 196926 143856 199328
rect 143908 198960 143960 198966
rect 143908 198902 143960 198908
rect 143816 196920 143868 196926
rect 143816 196862 143868 196868
rect 143644 196812 143764 196840
rect 143540 194200 143592 194206
rect 143540 194142 143592 194148
rect 143644 193712 143672 196812
rect 143724 196716 143776 196722
rect 143724 196658 143776 196664
rect 143552 193684 143672 193712
rect 143552 192506 143580 193684
rect 143632 193588 143684 193594
rect 143632 193530 143684 193536
rect 143540 192500 143592 192506
rect 143540 192442 143592 192448
rect 143448 191140 143500 191146
rect 143448 191082 143500 191088
rect 143540 154352 143592 154358
rect 143540 154294 143592 154300
rect 142988 151632 143040 151638
rect 142988 151574 143040 151580
rect 142712 148708 142764 148714
rect 142712 148650 142764 148656
rect 143552 146962 143580 154294
rect 143644 147082 143672 193530
rect 143736 147218 143764 196658
rect 143814 196480 143870 196489
rect 143814 196415 143870 196424
rect 143724 147212 143776 147218
rect 143724 147154 143776 147160
rect 143632 147076 143684 147082
rect 143632 147018 143684 147024
rect 143828 147014 143856 196415
rect 143920 196246 143948 198902
rect 143908 196240 143960 196246
rect 143908 196182 143960 196188
rect 144012 196178 144040 199543
rect 144104 198694 144132 199650
rect 144182 199608 144238 199617
rect 144182 199543 144238 199552
rect 144092 198688 144144 198694
rect 144092 198630 144144 198636
rect 144092 196240 144144 196246
rect 144092 196182 144144 196188
rect 144000 196172 144052 196178
rect 144000 196114 144052 196120
rect 143908 196104 143960 196110
rect 143908 196046 143960 196052
rect 143920 147150 143948 196046
rect 144104 193730 144132 196182
rect 144092 193724 144144 193730
rect 144092 193666 144144 193672
rect 144196 192778 144224 199543
rect 144288 199442 144316 199702
rect 144368 199640 144420 199646
rect 144368 199582 144420 199588
rect 144276 199436 144328 199442
rect 144276 199378 144328 199384
rect 144380 192846 144408 199582
rect 144472 197810 144500 199736
rect 144552 199708 144604 199714
rect 144552 199650 144604 199656
rect 144644 199708 144696 199714
rect 144644 199650 144696 199656
rect 144736 199708 144788 199714
rect 144736 199650 144788 199656
rect 144460 197804 144512 197810
rect 144460 197746 144512 197752
rect 144564 196314 144592 199650
rect 144656 197878 144684 199650
rect 144644 197872 144696 197878
rect 144644 197814 144696 197820
rect 144552 196308 144604 196314
rect 144552 196250 144604 196256
rect 144642 194440 144698 194449
rect 144642 194375 144698 194384
rect 144656 194342 144684 194375
rect 144644 194336 144696 194342
rect 144644 194278 144696 194284
rect 144368 192840 144420 192846
rect 144368 192782 144420 192788
rect 144184 192772 144236 192778
rect 144184 192714 144236 192720
rect 144748 190058 144776 199650
rect 144828 199640 144880 199646
rect 144828 199582 144880 199588
rect 144840 199102 144868 199582
rect 144828 199096 144880 199102
rect 144828 199038 144880 199044
rect 144932 196314 144960 199736
rect 145254 199764 145282 200124
rect 145346 199782 145374 200124
rect 145012 199718 145064 199724
rect 145102 199744 145158 199753
rect 144920 196308 144972 196314
rect 144920 196250 144972 196256
rect 144920 196172 144972 196178
rect 144920 196114 144972 196120
rect 144932 194546 144960 196114
rect 144920 194540 144972 194546
rect 144920 194482 144972 194488
rect 145024 193866 145052 199718
rect 145102 199679 145158 199688
rect 145208 199736 145282 199764
rect 145334 199776 145386 199782
rect 145116 199374 145144 199679
rect 145208 199374 145236 199736
rect 145334 199718 145386 199724
rect 145288 199572 145340 199578
rect 145438 199560 145466 200124
rect 145530 199923 145558 200124
rect 145516 199914 145572 199923
rect 145516 199849 145572 199858
rect 145622 199764 145650 200124
rect 145714 199918 145742 200124
rect 145702 199912 145754 199918
rect 145702 199854 145754 199860
rect 145806 199764 145834 200124
rect 145898 199918 145926 200124
rect 145886 199912 145938 199918
rect 145886 199854 145938 199860
rect 145990 199764 146018 200124
rect 146082 199918 146110 200124
rect 146174 199918 146202 200124
rect 146266 199918 146294 200124
rect 146070 199912 146122 199918
rect 146070 199854 146122 199860
rect 146162 199912 146214 199918
rect 146162 199854 146214 199860
rect 146254 199912 146306 199918
rect 146254 199854 146306 199860
rect 145288 199514 145340 199520
rect 145392 199532 145466 199560
rect 145576 199736 145650 199764
rect 145760 199736 145834 199764
rect 145944 199736 146018 199764
rect 146208 199776 146260 199782
rect 145104 199368 145156 199374
rect 145104 199310 145156 199316
rect 145196 199368 145248 199374
rect 145196 199310 145248 199316
rect 145300 198098 145328 199514
rect 145392 199238 145420 199532
rect 145470 199472 145526 199481
rect 145470 199407 145526 199416
rect 145380 199232 145432 199238
rect 145380 199174 145432 199180
rect 145484 198098 145512 199407
rect 145208 198070 145328 198098
rect 145392 198070 145512 198098
rect 145102 196888 145158 196897
rect 145102 196823 145158 196832
rect 145012 193860 145064 193866
rect 145012 193802 145064 193808
rect 145116 193662 145144 196823
rect 145208 195974 145236 198070
rect 145288 198008 145340 198014
rect 145288 197950 145340 197956
rect 145196 195968 145248 195974
rect 145196 195910 145248 195916
rect 145104 193656 145156 193662
rect 145104 193598 145156 193604
rect 144736 190052 144788 190058
rect 144736 189994 144788 190000
rect 145196 148436 145248 148442
rect 145196 148378 145248 148384
rect 143908 147144 143960 147150
rect 143908 147086 143960 147092
rect 143816 147008 143868 147014
rect 143552 146934 143764 146962
rect 143816 146950 143868 146956
rect 143632 145852 143684 145858
rect 143632 145794 143684 145800
rect 142526 144392 142582 144401
rect 142526 144327 142582 144336
rect 141424 143064 141476 143070
rect 141424 143006 141476 143012
rect 141206 140134 141280 140162
rect 132052 139862 132388 139890
rect 132696 139862 132940 139890
rect 133156 139862 133492 139890
rect 133892 139862 134044 139890
rect 134260 139862 134596 139890
rect 134812 139862 135148 139890
rect 135456 139862 135700 139890
rect 135824 139862 136252 139890
rect 136652 139862 136804 139890
rect 137020 139862 137356 139890
rect 137572 139862 137908 139890
rect 138124 139862 138460 139890
rect 138676 139862 139012 139890
rect 139412 139862 139564 139890
rect 139780 139862 140116 139890
rect 140332 139862 140668 139890
rect 141206 139876 141234 140134
rect 141436 139890 141464 143006
rect 142252 140956 142304 140962
rect 142252 140898 142304 140904
rect 142264 139890 142292 140898
rect 142540 139890 142568 144327
rect 143078 143032 143134 143041
rect 143078 142967 143134 142976
rect 143092 139890 143120 142967
rect 143644 139890 143672 145794
rect 143736 142154 143764 146934
rect 145012 145648 145064 145654
rect 145012 145590 145064 145596
rect 144920 142996 144972 143002
rect 144920 142938 144972 142944
rect 143736 142126 144224 142154
rect 144196 139890 144224 142126
rect 144932 139890 144960 142938
rect 145024 140758 145052 145590
rect 145012 140752 145064 140758
rect 145012 140694 145064 140700
rect 145208 139890 145236 148378
rect 145300 146946 145328 197950
rect 145392 195974 145420 198070
rect 145472 196036 145524 196042
rect 145472 195978 145524 195984
rect 145380 195968 145432 195974
rect 145380 195910 145432 195916
rect 145484 148646 145512 195978
rect 145576 194002 145604 199736
rect 145656 199436 145708 199442
rect 145656 199378 145708 199384
rect 145564 193996 145616 194002
rect 145564 193938 145616 193944
rect 145668 193934 145696 199378
rect 145656 193928 145708 193934
rect 145656 193870 145708 193876
rect 145760 191834 145788 199736
rect 145838 199608 145894 199617
rect 145838 199543 145894 199552
rect 145852 197266 145880 199543
rect 145944 199170 145972 199736
rect 146208 199718 146260 199724
rect 146024 199640 146076 199646
rect 146024 199582 146076 199588
rect 145932 199164 145984 199170
rect 145932 199106 145984 199112
rect 145840 197260 145892 197266
rect 145840 197202 145892 197208
rect 145840 196308 145892 196314
rect 145840 196250 145892 196256
rect 145576 191806 145788 191834
rect 145472 148640 145524 148646
rect 145472 148582 145524 148588
rect 145576 148578 145604 191806
rect 145852 180794 145880 196250
rect 146036 196042 146064 199582
rect 146116 199436 146168 199442
rect 146116 199378 146168 199384
rect 146128 196858 146156 199378
rect 146220 199306 146248 199718
rect 146358 199628 146386 200124
rect 146450 199918 146478 200124
rect 146542 199923 146570 200124
rect 146438 199912 146490 199918
rect 146438 199854 146490 199860
rect 146528 199914 146584 199923
rect 146528 199849 146584 199858
rect 146484 199776 146536 199782
rect 146484 199718 146536 199724
rect 146358 199600 146432 199628
rect 146300 199504 146352 199510
rect 146300 199446 146352 199452
rect 146208 199300 146260 199306
rect 146208 199242 146260 199248
rect 146312 198966 146340 199446
rect 146300 198960 146352 198966
rect 146300 198902 146352 198908
rect 146208 198008 146260 198014
rect 146208 197950 146260 197956
rect 146116 196852 146168 196858
rect 146116 196794 146168 196800
rect 146024 196036 146076 196042
rect 146024 195978 146076 195984
rect 145760 180766 145880 180794
rect 145564 148572 145616 148578
rect 145564 148514 145616 148520
rect 145288 146940 145340 146946
rect 145288 146882 145340 146888
rect 145760 144362 145788 180766
rect 146220 146946 146248 197950
rect 146404 196058 146432 199600
rect 146496 196178 146524 199718
rect 146634 199696 146662 200124
rect 146726 199923 146754 200124
rect 146712 199914 146768 199923
rect 146818 199918 146846 200124
rect 146910 199923 146938 200124
rect 146712 199849 146768 199858
rect 146806 199912 146858 199918
rect 146806 199854 146858 199860
rect 146896 199914 146952 199923
rect 147002 199918 147030 200124
rect 146896 199849 146952 199858
rect 146990 199912 147042 199918
rect 146990 199854 147042 199860
rect 147094 199764 147122 200124
rect 146588 199668 146662 199696
rect 146850 199744 146906 199753
rect 146850 199679 146906 199688
rect 147048 199736 147122 199764
rect 146588 196518 146616 199668
rect 146760 199640 146812 199646
rect 146760 199582 146812 199588
rect 146576 196512 146628 196518
rect 146576 196454 146628 196460
rect 146484 196172 146536 196178
rect 146484 196114 146536 196120
rect 146404 196030 146708 196058
rect 146576 195968 146628 195974
rect 146576 195910 146628 195916
rect 146392 154216 146444 154222
rect 146392 154158 146444 154164
rect 146404 151814 146432 154158
rect 146404 151786 146524 151814
rect 146208 146940 146260 146946
rect 146208 146882 146260 146888
rect 145748 144356 145800 144362
rect 145748 144298 145800 144304
rect 146392 142248 146444 142254
rect 146392 142190 146444 142196
rect 145840 140752 145892 140758
rect 145840 140694 145892 140700
rect 145852 139890 145880 140694
rect 146404 139890 146432 142190
rect 146496 142154 146524 151786
rect 146588 145790 146616 195910
rect 146680 148510 146708 196030
rect 146772 194478 146800 199582
rect 146864 198354 146892 199679
rect 147048 199209 147076 199736
rect 147186 199696 147214 200124
rect 147278 199923 147306 200124
rect 147264 199914 147320 199923
rect 147264 199849 147320 199858
rect 147370 199764 147398 200124
rect 147462 199923 147490 200124
rect 147448 199914 147504 199923
rect 147554 199918 147582 200124
rect 147646 199923 147674 200124
rect 147448 199849 147504 199858
rect 147542 199912 147594 199918
rect 147542 199854 147594 199860
rect 147632 199914 147688 199923
rect 147632 199849 147688 199858
rect 147496 199776 147548 199782
rect 147370 199736 147444 199764
rect 147140 199668 147214 199696
rect 147034 199200 147090 199209
rect 147034 199135 147090 199144
rect 147140 198490 147168 199668
rect 147312 199640 147364 199646
rect 147312 199582 147364 199588
rect 147128 198484 147180 198490
rect 147128 198426 147180 198432
rect 146852 198348 146904 198354
rect 146852 198290 146904 198296
rect 147220 196648 147272 196654
rect 147220 196590 147272 196596
rect 146760 194472 146812 194478
rect 146760 194414 146812 194420
rect 147232 192982 147260 196590
rect 147324 195566 147352 199582
rect 147416 196625 147444 199736
rect 147496 199718 147548 199724
rect 147738 199730 147766 200124
rect 147830 199850 147858 200124
rect 147922 199923 147950 200124
rect 147908 199914 147964 199923
rect 147818 199844 147870 199850
rect 147908 199849 147964 199858
rect 147818 199786 147870 199792
rect 147908 199778 147964 199787
rect 147402 196616 147458 196625
rect 147402 196551 147458 196560
rect 147312 195560 147364 195566
rect 147312 195502 147364 195508
rect 147508 193798 147536 199718
rect 147588 199708 147640 199714
rect 147738 199702 147812 199730
rect 148014 199764 148042 200124
rect 147964 199736 148042 199764
rect 147908 199713 147964 199722
rect 147588 199650 147640 199656
rect 147600 194410 147628 199650
rect 147678 199608 147734 199617
rect 147678 199543 147734 199552
rect 147784 199560 147812 199702
rect 148106 199696 148134 200124
rect 148014 199668 148134 199696
rect 147692 199034 147720 199543
rect 147784 199532 147904 199560
rect 147770 199472 147826 199481
rect 147770 199407 147826 199416
rect 147680 199028 147732 199034
rect 147680 198970 147732 198976
rect 147784 198558 147812 199407
rect 147876 198830 147904 199532
rect 148014 199492 148042 199668
rect 148198 199628 148226 200124
rect 148152 199600 148226 199628
rect 148014 199464 148088 199492
rect 147864 198824 147916 198830
rect 147864 198766 147916 198772
rect 147772 198552 147824 198558
rect 147772 198494 147824 198500
rect 147862 198112 147918 198121
rect 147862 198047 147918 198056
rect 147876 195702 147904 198047
rect 147864 195696 147916 195702
rect 147864 195638 147916 195644
rect 147588 194404 147640 194410
rect 147588 194346 147640 194352
rect 148060 194274 148088 199464
rect 148152 195770 148180 199600
rect 148290 199560 148318 200124
rect 148382 199714 148410 200124
rect 148474 199850 148502 200124
rect 148566 199923 148594 200124
rect 148552 199914 148608 199923
rect 148462 199844 148514 199850
rect 148552 199849 148608 199858
rect 148658 199850 148686 200124
rect 148750 199923 148778 200124
rect 148736 199914 148792 199923
rect 148462 199786 148514 199792
rect 148646 199844 148698 199850
rect 148736 199849 148792 199858
rect 148646 199786 148698 199792
rect 148842 199764 148870 200124
rect 148690 199744 148746 199753
rect 148370 199708 148422 199714
rect 148370 199650 148422 199656
rect 148600 199708 148652 199714
rect 148690 199679 148746 199688
rect 148796 199736 148870 199764
rect 148600 199650 148652 199656
rect 148244 199532 148318 199560
rect 148506 199608 148562 199617
rect 148506 199543 148562 199552
rect 148140 195764 148192 195770
rect 148140 195706 148192 195712
rect 148048 194268 148100 194274
rect 148048 194210 148100 194216
rect 147496 193792 147548 193798
rect 147496 193734 147548 193740
rect 147220 192976 147272 192982
rect 147220 192918 147272 192924
rect 148244 191834 148272 199532
rect 148324 199436 148376 199442
rect 148324 199378 148376 199384
rect 148336 196382 148364 199378
rect 148416 199368 148468 199374
rect 148416 199310 148468 199316
rect 148428 198150 148456 199310
rect 148416 198144 148468 198150
rect 148416 198086 148468 198092
rect 148324 196376 148376 196382
rect 148324 196318 148376 196324
rect 148152 191806 148272 191834
rect 146668 148504 146720 148510
rect 146668 148446 146720 148452
rect 146576 145784 146628 145790
rect 146576 145726 146628 145732
rect 147770 145616 147826 145625
rect 147770 145551 147826 145560
rect 147678 144528 147734 144537
rect 147678 144463 147734 144472
rect 147692 143546 147720 144463
rect 147680 143540 147732 143546
rect 147680 143482 147732 143488
rect 146496 142126 146892 142154
rect 146864 139890 146892 142126
rect 147784 139890 147812 145551
rect 148048 142928 148100 142934
rect 148048 142870 148100 142876
rect 148060 139890 148088 142870
rect 148152 140078 148180 191806
rect 148520 180794 148548 199543
rect 148612 195022 148640 199650
rect 148704 196722 148732 199679
rect 148692 196716 148744 196722
rect 148692 196658 148744 196664
rect 148600 195016 148652 195022
rect 148600 194958 148652 194964
rect 148796 180794 148824 199736
rect 148934 199696 148962 200124
rect 148888 199668 148962 199696
rect 148888 194585 148916 199668
rect 149026 199628 149054 200124
rect 149118 199918 149146 200124
rect 149210 199918 149238 200124
rect 149106 199912 149158 199918
rect 149106 199854 149158 199860
rect 149198 199912 149250 199918
rect 149198 199854 149250 199860
rect 149302 199764 149330 200124
rect 149394 199923 149422 200124
rect 149380 199914 149436 199923
rect 149486 199918 149514 200124
rect 149578 199923 149606 200124
rect 149380 199849 149436 199858
rect 149474 199912 149526 199918
rect 149474 199854 149526 199860
rect 149564 199914 149620 199923
rect 149564 199849 149620 199858
rect 149670 199850 149698 200124
rect 149658 199844 149710 199850
rect 149658 199786 149710 199792
rect 149256 199736 149330 199764
rect 149152 199708 149204 199714
rect 149152 199650 149204 199656
rect 148980 199600 149054 199628
rect 148980 195838 149008 199600
rect 149060 199504 149112 199510
rect 149060 199446 149112 199452
rect 149072 198762 149100 199446
rect 149060 198756 149112 198762
rect 149060 198698 149112 198704
rect 149164 195906 149192 199650
rect 149256 197878 149284 199736
rect 149612 199640 149664 199646
rect 149334 199608 149390 199617
rect 149518 199608 149574 199617
rect 149334 199543 149390 199552
rect 149428 199572 149480 199578
rect 149348 198626 149376 199543
rect 149762 199628 149790 200124
rect 149854 199918 149882 200124
rect 149842 199912 149894 199918
rect 149842 199854 149894 199860
rect 149946 199730 149974 200124
rect 150038 199918 150066 200124
rect 150130 199923 150158 200124
rect 150026 199912 150078 199918
rect 150026 199854 150078 199860
rect 150116 199914 150172 199923
rect 150222 199918 150250 200124
rect 150116 199849 150172 199858
rect 150210 199912 150262 199918
rect 150210 199854 150262 199860
rect 150314 199850 150342 200124
rect 150406 199889 150434 200124
rect 150498 199918 150526 200124
rect 150590 199918 150618 200124
rect 150682 199918 150710 200124
rect 150774 199923 150802 200124
rect 150486 199912 150538 199918
rect 150392 199880 150448 199889
rect 150302 199844 150354 199850
rect 150486 199854 150538 199860
rect 150578 199912 150630 199918
rect 150578 199854 150630 199860
rect 150670 199912 150722 199918
rect 150670 199854 150722 199860
rect 150760 199914 150816 199923
rect 150760 199849 150816 199858
rect 150866 199850 150894 200124
rect 150958 199918 150986 200124
rect 151050 199918 151078 200124
rect 150946 199912 150998 199918
rect 150946 199854 150998 199860
rect 151038 199912 151090 199918
rect 151038 199854 151090 199860
rect 150392 199815 150448 199824
rect 150854 199844 150906 199850
rect 150302 199786 150354 199792
rect 150854 199786 150906 199792
rect 149900 199702 149974 199730
rect 150440 199776 150492 199782
rect 150440 199718 150492 199724
rect 150532 199776 150584 199782
rect 151142 199764 151170 200124
rect 151234 199918 151262 200124
rect 151326 199918 151354 200124
rect 151418 199918 151446 200124
rect 151222 199912 151274 199918
rect 151222 199854 151274 199860
rect 151314 199912 151366 199918
rect 151314 199854 151366 199860
rect 151406 199912 151458 199918
rect 151510 199889 151538 200124
rect 151406 199854 151458 199860
rect 151496 199880 151552 199889
rect 151496 199815 151552 199824
rect 151452 199776 151504 199782
rect 150532 199718 150584 199724
rect 150622 199744 150678 199753
rect 150256 199708 150308 199714
rect 149762 199600 149836 199628
rect 149612 199582 149664 199588
rect 149518 199543 149574 199552
rect 149428 199514 149480 199520
rect 149336 198620 149388 198626
rect 149336 198562 149388 198568
rect 149440 198422 149468 199514
rect 149532 199306 149560 199543
rect 149520 199300 149572 199306
rect 149520 199242 149572 199248
rect 149428 198416 149480 198422
rect 149428 198358 149480 198364
rect 149336 198076 149388 198082
rect 149336 198018 149388 198024
rect 149244 197872 149296 197878
rect 149244 197814 149296 197820
rect 149348 196704 149376 198018
rect 149624 197946 149652 199582
rect 149702 199472 149758 199481
rect 149702 199407 149758 199416
rect 149612 197940 149664 197946
rect 149612 197882 149664 197888
rect 149256 196676 149376 196704
rect 149152 195900 149204 195906
rect 149152 195842 149204 195848
rect 148968 195832 149020 195838
rect 148968 195774 149020 195780
rect 148874 194576 148930 194585
rect 148874 194511 148930 194520
rect 148244 180766 148548 180794
rect 148612 180766 148824 180794
rect 148244 145722 148272 180766
rect 148612 148345 148640 180766
rect 149256 148617 149284 196676
rect 149336 196580 149388 196586
rect 149336 196522 149388 196528
rect 149348 187134 149376 196522
rect 149716 195673 149744 199407
rect 149808 197606 149836 199600
rect 149900 198082 149928 199702
rect 150256 199650 150308 199656
rect 150164 199640 150216 199646
rect 149978 199608 150034 199617
rect 150164 199582 150216 199588
rect 149978 199543 150034 199552
rect 150072 199572 150124 199578
rect 149888 198076 149940 198082
rect 149888 198018 149940 198024
rect 149888 197940 149940 197946
rect 149888 197882 149940 197888
rect 149796 197600 149848 197606
rect 149796 197542 149848 197548
rect 149796 197464 149848 197470
rect 149796 197406 149848 197412
rect 149702 195664 149758 195673
rect 149702 195599 149758 195608
rect 149704 193588 149756 193594
rect 149704 193530 149756 193536
rect 149336 187128 149388 187134
rect 149336 187070 149388 187076
rect 149716 148782 149744 193530
rect 149808 149054 149836 197406
rect 149900 191834 149928 197882
rect 149992 197810 150020 199543
rect 150072 199514 150124 199520
rect 149980 197804 150032 197810
rect 149980 197746 150032 197752
rect 150084 197690 150112 199514
rect 149992 197662 150112 197690
rect 149992 195430 150020 197662
rect 150072 197600 150124 197606
rect 150072 197542 150124 197548
rect 149980 195424 150032 195430
rect 149980 195366 150032 195372
rect 149900 191806 150020 191834
rect 149888 191004 149940 191010
rect 149888 190946 149940 190952
rect 149796 149048 149848 149054
rect 149796 148990 149848 148996
rect 149704 148776 149756 148782
rect 149704 148718 149756 148724
rect 149242 148608 149298 148617
rect 149242 148543 149298 148552
rect 148598 148336 148654 148345
rect 148598 148271 148654 148280
rect 149058 145888 149114 145897
rect 149058 145823 149114 145832
rect 148232 145716 148284 145722
rect 148232 145658 148284 145664
rect 148598 144120 148654 144129
rect 148598 144055 148654 144064
rect 148140 140072 148192 140078
rect 148140 140014 148192 140020
rect 148612 139890 148640 144055
rect 149072 139890 149100 145823
rect 149704 142860 149756 142866
rect 149704 142802 149756 142808
rect 149716 139890 149744 142802
rect 149900 141438 149928 190946
rect 149992 190466 150020 191806
rect 149980 190460 150032 190466
rect 149980 190402 150032 190408
rect 150084 144634 150112 197542
rect 150176 191010 150204 199582
rect 150268 196586 150296 199650
rect 150256 196580 150308 196586
rect 150256 196522 150308 196528
rect 150452 193594 150480 199718
rect 150440 193588 150492 193594
rect 150440 193530 150492 193536
rect 150544 192778 150572 199718
rect 151142 199736 151308 199764
rect 150622 199679 150678 199688
rect 150716 199708 150768 199714
rect 150636 199374 150664 199679
rect 150716 199650 150768 199656
rect 150808 199708 150860 199714
rect 151280 199696 151308 199736
rect 151602 199764 151630 200124
rect 151694 199918 151722 200124
rect 151682 199912 151734 199918
rect 151682 199854 151734 199860
rect 151452 199718 151504 199724
rect 151556 199736 151630 199764
rect 151786 199764 151814 200124
rect 151878 199918 151906 200124
rect 151970 199923 151998 200124
rect 151866 199912 151918 199918
rect 151866 199854 151918 199860
rect 151956 199914 152012 199923
rect 152062 199918 152090 200124
rect 152154 199918 152182 200124
rect 152246 199918 152274 200124
rect 151956 199849 152012 199858
rect 152050 199912 152102 199918
rect 152050 199854 152102 199860
rect 152142 199912 152194 199918
rect 152142 199854 152194 199860
rect 152234 199912 152286 199918
rect 152234 199854 152286 199860
rect 152338 199764 152366 200124
rect 152430 199850 152458 200124
rect 152418 199844 152470 199850
rect 152418 199786 152470 199792
rect 151786 199736 151860 199764
rect 151280 199668 151400 199696
rect 150808 199650 150860 199656
rect 150624 199368 150676 199374
rect 150624 199310 150676 199316
rect 150728 199034 150756 199650
rect 150716 199028 150768 199034
rect 150716 198970 150768 198976
rect 150624 193180 150676 193186
rect 150624 193122 150676 193128
rect 150532 192772 150584 192778
rect 150532 192714 150584 192720
rect 150164 191004 150216 191010
rect 150164 190946 150216 190952
rect 150636 151162 150664 193122
rect 150820 186998 150848 199650
rect 151084 199640 151136 199646
rect 151084 199582 151136 199588
rect 151176 199640 151228 199646
rect 151176 199582 151228 199588
rect 151096 199345 151124 199582
rect 151082 199336 151138 199345
rect 151082 199271 151138 199280
rect 151084 197804 151136 197810
rect 151084 197746 151136 197752
rect 150992 195764 151044 195770
rect 150992 195706 151044 195712
rect 150808 186992 150860 186998
rect 150808 186934 150860 186940
rect 150624 151156 150676 151162
rect 150624 151098 150676 151104
rect 150072 144628 150124 144634
rect 150072 144570 150124 144576
rect 150808 143540 150860 143546
rect 150808 143482 150860 143488
rect 150532 142180 150584 142186
rect 150532 142122 150584 142128
rect 149888 141432 149940 141438
rect 149888 141374 149940 141380
rect 150544 139890 150572 142122
rect 150820 139890 150848 143482
rect 151004 140146 151032 195706
rect 151096 187066 151124 197746
rect 151188 196897 151216 199582
rect 151268 199572 151320 199578
rect 151268 199514 151320 199520
rect 151174 196888 151230 196897
rect 151174 196823 151230 196832
rect 151084 187060 151136 187066
rect 151084 187002 151136 187008
rect 151280 141438 151308 199514
rect 151372 196654 151400 199668
rect 151360 196648 151412 196654
rect 151464 196625 151492 199718
rect 151360 196590 151412 196596
rect 151450 196616 151506 196625
rect 151450 196551 151506 196560
rect 151556 193186 151584 199736
rect 151636 199640 151688 199646
rect 151636 199582 151688 199588
rect 151648 195770 151676 199582
rect 151728 198212 151780 198218
rect 151728 198154 151780 198160
rect 151636 195764 151688 195770
rect 151636 195706 151688 195712
rect 151544 193180 151596 193186
rect 151544 193122 151596 193128
rect 151740 148345 151768 198154
rect 151832 197130 151860 199736
rect 152292 199736 152366 199764
rect 151912 199708 151964 199714
rect 151912 199650 151964 199656
rect 152096 199708 152148 199714
rect 152096 199650 152148 199656
rect 152188 199708 152240 199714
rect 152188 199650 152240 199656
rect 151820 197124 151872 197130
rect 151820 197066 151872 197072
rect 151924 196874 151952 199650
rect 151924 196846 152044 196874
rect 151820 196648 151872 196654
rect 151820 196590 151872 196596
rect 151726 148336 151782 148345
rect 151726 148271 151782 148280
rect 151832 144566 151860 196590
rect 151912 196308 151964 196314
rect 151912 196250 151964 196256
rect 151924 148209 151952 196250
rect 152016 148481 152044 196846
rect 152108 158098 152136 199650
rect 152200 191146 152228 199650
rect 152292 198966 152320 199736
rect 152522 199696 152550 200124
rect 152614 199764 152642 200124
rect 152706 199918 152734 200124
rect 152798 199918 152826 200124
rect 152694 199912 152746 199918
rect 152694 199854 152746 199860
rect 152786 199912 152838 199918
rect 152786 199854 152838 199860
rect 152740 199776 152792 199782
rect 152614 199736 152688 199764
rect 152476 199668 152550 199696
rect 152372 199640 152424 199646
rect 152372 199582 152424 199588
rect 152280 198960 152332 198966
rect 152280 198902 152332 198908
rect 152384 196654 152412 199582
rect 152476 197033 152504 199668
rect 152660 199209 152688 199736
rect 152890 199764 152918 200124
rect 152982 199918 153010 200124
rect 153074 199918 153102 200124
rect 153166 199918 153194 200124
rect 153258 199923 153286 200124
rect 152970 199912 153022 199918
rect 152970 199854 153022 199860
rect 153062 199912 153114 199918
rect 153062 199854 153114 199860
rect 153154 199912 153206 199918
rect 153154 199854 153206 199860
rect 153244 199914 153300 199923
rect 153350 199918 153378 200124
rect 153442 199918 153470 200124
rect 153534 199923 153562 200124
rect 153244 199849 153300 199858
rect 153338 199912 153390 199918
rect 153338 199854 153390 199860
rect 153430 199912 153482 199918
rect 153430 199854 153482 199860
rect 153520 199914 153576 199923
rect 153626 199918 153654 200124
rect 153718 199918 153746 200124
rect 153810 199923 153838 200124
rect 153520 199849 153576 199858
rect 153614 199912 153666 199918
rect 153614 199854 153666 199860
rect 153706 199912 153758 199918
rect 153706 199854 153758 199860
rect 153796 199914 153852 199923
rect 153796 199849 153852 199858
rect 152740 199718 152792 199724
rect 152844 199736 152918 199764
rect 153016 199776 153068 199782
rect 152646 199200 152702 199209
rect 152646 199135 152702 199144
rect 152462 197024 152518 197033
rect 152462 196959 152518 196968
rect 152372 196648 152424 196654
rect 152372 196590 152424 196596
rect 152648 196648 152700 196654
rect 152648 196590 152700 196596
rect 152660 192250 152688 196590
rect 152752 192681 152780 199718
rect 152738 192672 152794 192681
rect 152738 192607 152794 192616
rect 152292 192222 152688 192250
rect 152188 191140 152240 191146
rect 152188 191082 152240 191088
rect 152292 191026 152320 192222
rect 152200 190998 152320 191026
rect 152096 158092 152148 158098
rect 152096 158034 152148 158040
rect 152200 158030 152228 190998
rect 152844 187202 152872 199736
rect 153016 199718 153068 199724
rect 153108 199776 153160 199782
rect 153108 199718 153160 199724
rect 153200 199776 153252 199782
rect 153200 199718 153252 199724
rect 153384 199776 153436 199782
rect 153384 199718 153436 199724
rect 153568 199776 153620 199782
rect 153568 199718 153620 199724
rect 152924 199640 152976 199646
rect 152924 199582 152976 199588
rect 152936 196654 152964 199582
rect 152924 196648 152976 196654
rect 152924 196590 152976 196596
rect 153028 196314 153056 199718
rect 153120 199617 153148 199718
rect 153106 199608 153162 199617
rect 153106 199543 153162 199552
rect 153212 196897 153240 199718
rect 153198 196888 153254 196897
rect 153198 196823 153254 196832
rect 153016 196308 153068 196314
rect 153016 196250 153068 196256
rect 153396 194342 153424 199718
rect 153476 199708 153528 199714
rect 153476 199650 153528 199656
rect 153488 199617 153516 199650
rect 153474 199608 153530 199617
rect 153474 199543 153530 199552
rect 153580 198744 153608 199718
rect 153902 199696 153930 200124
rect 153994 199918 154022 200124
rect 154086 199918 154114 200124
rect 154178 199918 154206 200124
rect 154270 199918 154298 200124
rect 153982 199912 154034 199918
rect 153982 199854 154034 199860
rect 154074 199912 154126 199918
rect 154074 199854 154126 199860
rect 154166 199912 154218 199918
rect 154166 199854 154218 199860
rect 154258 199912 154310 199918
rect 154258 199854 154310 199860
rect 154118 199744 154174 199753
rect 153856 199668 153930 199696
rect 154028 199708 154080 199714
rect 153660 199640 153712 199646
rect 153660 199582 153712 199588
rect 153672 198937 153700 199582
rect 153658 198928 153714 198937
rect 153658 198863 153714 198872
rect 153580 198716 153700 198744
rect 153474 198112 153530 198121
rect 153474 198047 153530 198056
rect 153488 195974 153516 198047
rect 153566 197976 153622 197985
rect 153566 197911 153622 197920
rect 153476 195968 153528 195974
rect 153476 195910 153528 195916
rect 153476 195832 153528 195838
rect 153476 195774 153528 195780
rect 153384 194336 153436 194342
rect 153384 194278 153436 194284
rect 153292 193996 153344 194002
rect 153292 193938 153344 193944
rect 152832 187196 152884 187202
rect 152832 187138 152884 187144
rect 152188 158024 152240 158030
rect 152188 157966 152240 157972
rect 152002 148472 152058 148481
rect 152002 148407 152058 148416
rect 151910 148200 151966 148209
rect 151910 148135 151966 148144
rect 151820 144560 151872 144566
rect 151820 144502 151872 144508
rect 152464 144492 152516 144498
rect 152464 144434 152516 144440
rect 151912 144424 151964 144430
rect 151912 144366 151964 144372
rect 151358 142760 151414 142769
rect 151358 142695 151414 142704
rect 151268 141432 151320 141438
rect 151268 141374 151320 141380
rect 150992 140140 151044 140146
rect 150992 140082 151044 140088
rect 151372 139890 151400 142695
rect 151924 139890 151952 144366
rect 152476 139890 152504 144434
rect 153304 141545 153332 193938
rect 153488 145761 153516 195774
rect 153580 148753 153608 197911
rect 153672 196058 153700 198716
rect 153672 196030 153792 196058
rect 153660 195968 153712 195974
rect 153764 195945 153792 196030
rect 153660 195910 153712 195916
rect 153750 195936 153806 195945
rect 153672 190454 153700 195910
rect 153750 195871 153806 195880
rect 153856 192545 153884 199668
rect 154362 199696 154390 200124
rect 154454 199918 154482 200124
rect 154546 199923 154574 200124
rect 154442 199912 154494 199918
rect 154442 199854 154494 199860
rect 154532 199914 154588 199923
rect 154532 199849 154588 199858
rect 154638 199850 154666 200124
rect 154730 199850 154758 200124
rect 154626 199844 154678 199850
rect 154626 199786 154678 199792
rect 154718 199844 154770 199850
rect 154718 199786 154770 199792
rect 154118 199679 154174 199688
rect 154028 199650 154080 199656
rect 153934 199608 153990 199617
rect 153934 199543 153990 199552
rect 153948 197470 153976 199543
rect 153936 197464 153988 197470
rect 153936 197406 153988 197412
rect 154040 194002 154068 199650
rect 154132 199578 154160 199679
rect 154316 199668 154390 199696
rect 154212 199640 154264 199646
rect 154212 199582 154264 199588
rect 154120 199572 154172 199578
rect 154120 199514 154172 199520
rect 154224 195401 154252 199582
rect 154316 195838 154344 199668
rect 154532 199642 154588 199651
rect 154822 199628 154850 200124
rect 154914 199923 154942 200124
rect 154900 199914 154956 199923
rect 154900 199849 154956 199858
rect 155006 199764 155034 200124
rect 155098 199918 155126 200124
rect 155086 199912 155138 199918
rect 155086 199854 155138 199860
rect 155190 199764 155218 200124
rect 155006 199736 155080 199764
rect 154396 199572 154448 199578
rect 154532 199577 154588 199586
rect 154776 199600 154850 199628
rect 154396 199514 154448 199520
rect 154304 195832 154356 195838
rect 154304 195774 154356 195780
rect 154302 195664 154358 195673
rect 154302 195599 154358 195608
rect 154210 195392 154266 195401
rect 154210 195327 154266 195336
rect 154028 193996 154080 194002
rect 154028 193938 154080 193944
rect 153842 192536 153898 192545
rect 153842 192471 153898 192480
rect 153672 190426 154068 190454
rect 153658 151328 153714 151337
rect 153658 151263 153714 151272
rect 153566 148744 153622 148753
rect 153566 148679 153622 148688
rect 153474 145752 153530 145761
rect 153474 145687 153530 145696
rect 153290 141536 153346 141545
rect 153290 141471 153346 141480
rect 153672 139890 153700 151263
rect 153752 141568 153804 141574
rect 153752 141510 153804 141516
rect 141436 139862 141772 139890
rect 142264 139862 142324 139890
rect 142540 139862 142876 139890
rect 143092 139862 143428 139890
rect 143644 139862 143980 139890
rect 144196 139862 144532 139890
rect 144932 139862 145084 139890
rect 145208 139862 145636 139890
rect 145852 139862 146188 139890
rect 146404 139862 146740 139890
rect 146864 139862 147292 139890
rect 147784 139862 147844 139890
rect 148060 139862 148396 139890
rect 148612 139862 148948 139890
rect 149072 139862 149500 139890
rect 149716 139862 150052 139890
rect 150544 139862 150604 139890
rect 150820 139862 151156 139890
rect 151372 139862 151708 139890
rect 151924 139862 152260 139890
rect 152476 139862 152812 139890
rect 153364 139862 153700 139890
rect 153764 139890 153792 141510
rect 154040 141409 154068 190426
rect 154316 143002 154344 195599
rect 154408 189786 154436 199514
rect 154672 199504 154724 199510
rect 154500 199481 154620 199492
rect 154500 199472 154634 199481
rect 154500 199464 154578 199472
rect 154500 195430 154528 199464
rect 154672 199446 154724 199452
rect 154578 199407 154634 199416
rect 154684 199356 154712 199446
rect 154592 199328 154712 199356
rect 154592 199102 154620 199328
rect 154580 199096 154632 199102
rect 154580 199038 154632 199044
rect 154776 198830 154804 199600
rect 154948 199572 155000 199578
rect 154948 199514 155000 199520
rect 154856 199504 154908 199510
rect 154856 199446 154908 199452
rect 154764 198824 154816 198830
rect 154764 198766 154816 198772
rect 154868 198694 154896 199446
rect 154856 198688 154908 198694
rect 154856 198630 154908 198636
rect 154672 196988 154724 196994
rect 154672 196930 154724 196936
rect 154580 195492 154632 195498
rect 154580 195434 154632 195440
rect 154488 195424 154540 195430
rect 154488 195366 154540 195372
rect 154592 191418 154620 195434
rect 154580 191412 154632 191418
rect 154580 191354 154632 191360
rect 154396 189780 154448 189786
rect 154396 189722 154448 189728
rect 154684 151094 154712 196930
rect 154764 196648 154816 196654
rect 154764 196590 154816 196596
rect 154776 187270 154804 196590
rect 154960 196586 154988 199514
rect 154948 196580 155000 196586
rect 154948 196522 155000 196528
rect 155052 195498 155080 199736
rect 155144 199736 155218 199764
rect 155040 195492 155092 195498
rect 155040 195434 155092 195440
rect 155144 195090 155172 199736
rect 155282 199696 155310 200124
rect 155374 199850 155402 200124
rect 155466 199923 155494 200124
rect 155452 199914 155508 199923
rect 155362 199844 155414 199850
rect 155452 199849 155508 199858
rect 155362 199786 155414 199792
rect 155236 199668 155310 199696
rect 155406 199744 155462 199753
rect 155558 199730 155586 200124
rect 155650 199850 155678 200124
rect 155742 199889 155770 200124
rect 155728 199880 155784 199889
rect 155638 199844 155690 199850
rect 155834 199850 155862 200124
rect 155926 199923 155954 200124
rect 155912 199914 155968 199923
rect 155728 199815 155784 199824
rect 155822 199844 155874 199850
rect 155912 199849 155968 199858
rect 156018 199850 156046 200124
rect 156110 199923 156138 200124
rect 156096 199914 156152 199923
rect 155638 199786 155690 199792
rect 155822 199786 155874 199792
rect 156006 199844 156058 199850
rect 156096 199849 156152 199858
rect 156202 199850 156230 200124
rect 156294 199850 156322 200124
rect 156006 199786 156058 199792
rect 156190 199844 156242 199850
rect 156190 199786 156242 199792
rect 156282 199844 156334 199850
rect 156282 199786 156334 199792
rect 155406 199679 155462 199688
rect 155512 199702 155586 199730
rect 155958 199744 156014 199753
rect 155684 199708 155736 199714
rect 155132 195084 155184 195090
rect 155132 195026 155184 195032
rect 155236 192506 155264 199668
rect 155316 199572 155368 199578
rect 155316 199514 155368 199520
rect 155328 196926 155356 199514
rect 155420 196994 155448 199679
rect 155408 196988 155460 196994
rect 155408 196930 155460 196936
rect 155316 196920 155368 196926
rect 155316 196862 155368 196868
rect 155512 196840 155540 199702
rect 155684 199650 155736 199656
rect 155868 199708 155920 199714
rect 156142 199744 156198 199753
rect 155958 199679 156014 199688
rect 156052 199708 156104 199714
rect 155868 199650 155920 199656
rect 155592 199640 155644 199646
rect 155590 199608 155592 199617
rect 155644 199608 155646 199617
rect 155590 199543 155646 199552
rect 155420 196812 155540 196840
rect 155224 192500 155276 192506
rect 155224 192442 155276 192448
rect 155420 189854 155448 196812
rect 155500 196716 155552 196722
rect 155500 196658 155552 196664
rect 155408 189848 155460 189854
rect 155408 189790 155460 189796
rect 154764 187264 154816 187270
rect 154764 187206 154816 187212
rect 154764 151224 154816 151230
rect 154764 151166 154816 151172
rect 154672 151088 154724 151094
rect 154672 151030 154724 151036
rect 154488 144492 154540 144498
rect 154488 144434 154540 144440
rect 154304 142996 154356 143002
rect 154304 142938 154356 142944
rect 154026 141400 154082 141409
rect 154026 141335 154082 141344
rect 154500 140162 154528 144434
rect 154454 140134 154528 140162
rect 153764 139862 153916 139890
rect 154454 139876 154482 140134
rect 154776 139890 154804 151166
rect 155512 142866 155540 196658
rect 155696 196654 155724 199650
rect 155774 199608 155830 199617
rect 155774 199543 155830 199552
rect 155788 198082 155816 199543
rect 155776 198076 155828 198082
rect 155776 198018 155828 198024
rect 155684 196648 155736 196654
rect 155684 196590 155736 196596
rect 155684 195084 155736 195090
rect 155684 195026 155736 195032
rect 155696 148374 155724 195026
rect 155880 192574 155908 199650
rect 155972 199073 156000 199679
rect 156386 199730 156414 200124
rect 156478 199753 156506 200124
rect 156570 199918 156598 200124
rect 156662 199923 156690 200124
rect 156558 199912 156610 199918
rect 156558 199854 156610 199860
rect 156648 199914 156704 199923
rect 156648 199849 156704 199858
rect 156142 199679 156198 199688
rect 156236 199708 156288 199714
rect 156052 199650 156104 199656
rect 155958 199064 156014 199073
rect 155958 198999 156014 199008
rect 156064 197606 156092 199650
rect 156052 197600 156104 197606
rect 156052 197542 156104 197548
rect 156052 197396 156104 197402
rect 156052 197338 156104 197344
rect 155960 194948 156012 194954
rect 155960 194890 156012 194896
rect 155868 192568 155920 192574
rect 155868 192510 155920 192516
rect 155684 148368 155736 148374
rect 155684 148310 155736 148316
rect 155972 145858 156000 194890
rect 155960 145852 156012 145858
rect 155960 145794 156012 145800
rect 156064 145654 156092 197338
rect 156156 194410 156184 199679
rect 156236 199650 156288 199656
rect 156340 199702 156414 199730
rect 156464 199744 156520 199753
rect 156248 199442 156276 199650
rect 156236 199436 156288 199442
rect 156236 199378 156288 199384
rect 156236 198144 156288 198150
rect 156236 198086 156288 198092
rect 156248 195974 156276 198086
rect 156236 195968 156288 195974
rect 156236 195910 156288 195916
rect 156236 195832 156288 195838
rect 156236 195774 156288 195780
rect 156144 194404 156196 194410
rect 156144 194346 156196 194352
rect 156248 151502 156276 195774
rect 156340 189650 156368 199702
rect 156464 199679 156520 199688
rect 156602 199744 156658 199753
rect 156754 199730 156782 200124
rect 156846 199787 156874 200124
rect 156602 199679 156658 199688
rect 156708 199702 156782 199730
rect 156832 199778 156888 199787
rect 156938 199782 156966 200124
rect 156832 199713 156888 199722
rect 156926 199776 156978 199782
rect 157030 199764 157058 200124
rect 157122 199923 157150 200124
rect 157108 199914 157164 199923
rect 157108 199849 157164 199858
rect 157214 199787 157242 200124
rect 157306 199850 157334 200124
rect 157398 199850 157426 200124
rect 157490 199918 157518 200124
rect 157478 199912 157530 199918
rect 157478 199854 157530 199860
rect 157294 199844 157346 199850
rect 157200 199778 157256 199787
rect 157294 199786 157346 199792
rect 157386 199844 157438 199850
rect 157386 199786 157438 199792
rect 157030 199736 157104 199764
rect 156926 199718 156978 199724
rect 156512 199640 156564 199646
rect 156512 199582 156564 199588
rect 156418 199472 156474 199481
rect 156418 199407 156474 199416
rect 156432 199102 156460 199407
rect 156420 199096 156472 199102
rect 156420 199038 156472 199044
rect 156524 195838 156552 199582
rect 156616 197402 156644 199679
rect 156708 199102 156736 199702
rect 156880 199640 156932 199646
rect 156786 199608 156842 199617
rect 156880 199582 156932 199588
rect 156786 199543 156842 199552
rect 156696 199096 156748 199102
rect 156696 199038 156748 199044
rect 156604 197396 156656 197402
rect 156604 197338 156656 197344
rect 156604 196580 156656 196586
rect 156604 196522 156656 196528
rect 156512 195832 156564 195838
rect 156512 195774 156564 195780
rect 156616 191834 156644 196522
rect 156800 194954 156828 199543
rect 156788 194948 156840 194954
rect 156788 194890 156840 194896
rect 156892 192642 156920 199582
rect 157076 195498 157104 199736
rect 157582 199764 157610 200124
rect 157674 199918 157702 200124
rect 157766 199923 157794 200124
rect 157662 199912 157714 199918
rect 157662 199854 157714 199860
rect 157752 199914 157808 199923
rect 157752 199849 157808 199858
rect 157200 199713 157256 199722
rect 157536 199736 157610 199764
rect 157432 199708 157484 199714
rect 157432 199650 157484 199656
rect 157156 199640 157208 199646
rect 157156 199582 157208 199588
rect 157340 199640 157392 199646
rect 157340 199582 157392 199588
rect 157168 198937 157196 199582
rect 157248 199504 157300 199510
rect 157248 199446 157300 199452
rect 157260 199238 157288 199446
rect 157248 199232 157300 199238
rect 157248 199174 157300 199180
rect 157154 198928 157210 198937
rect 157154 198863 157210 198872
rect 157352 198762 157380 199582
rect 157340 198756 157392 198762
rect 157340 198698 157392 198704
rect 157444 197674 157472 199650
rect 157536 199617 157564 199736
rect 157858 199730 157886 200124
rect 157950 199782 157978 200124
rect 157708 199708 157760 199714
rect 157708 199650 157760 199656
rect 157812 199702 157886 199730
rect 157938 199776 157990 199782
rect 158042 199753 158070 200124
rect 158134 199918 158162 200124
rect 158122 199912 158174 199918
rect 158122 199854 158174 199860
rect 158122 199776 158174 199782
rect 157938 199718 157990 199724
rect 158028 199744 158084 199753
rect 157522 199608 157578 199617
rect 157522 199543 157578 199552
rect 157524 199504 157576 199510
rect 157524 199446 157576 199452
rect 157616 199504 157668 199510
rect 157616 199446 157668 199452
rect 157432 197668 157484 197674
rect 157432 197610 157484 197616
rect 157248 197260 157300 197266
rect 157248 197202 157300 197208
rect 157154 196888 157210 196897
rect 157154 196823 157210 196832
rect 157064 195492 157116 195498
rect 157064 195434 157116 195440
rect 156880 192636 156932 192642
rect 156880 192578 156932 192584
rect 156616 191806 156736 191834
rect 156708 190454 156736 191806
rect 156708 190426 156828 190454
rect 156328 189644 156380 189650
rect 156328 189586 156380 189592
rect 156236 151496 156288 151502
rect 156236 151438 156288 151444
rect 156236 147212 156288 147218
rect 156236 147154 156288 147160
rect 156052 145648 156104 145654
rect 156052 145590 156104 145596
rect 156142 144256 156198 144265
rect 156142 144191 156198 144200
rect 155500 142860 155552 142866
rect 155500 142802 155552 142808
rect 155868 142180 155920 142186
rect 155868 142122 155920 142128
rect 155880 139890 155908 142122
rect 156156 140162 156184 144191
rect 154776 139862 155020 139890
rect 155572 139862 155908 139890
rect 156110 140134 156184 140162
rect 156110 139876 156138 140134
rect 156248 139890 156276 147154
rect 156800 140078 156828 190426
rect 157168 148578 157196 196823
rect 157156 148572 157208 148578
rect 157156 148514 157208 148520
rect 157260 147014 157288 197202
rect 157536 196722 157564 199446
rect 157524 196716 157576 196722
rect 157524 196658 157576 196664
rect 157338 196616 157394 196625
rect 157338 196551 157394 196560
rect 157248 147008 157300 147014
rect 157248 146950 157300 146956
rect 157352 146962 157380 196551
rect 157432 195900 157484 195906
rect 157432 195842 157484 195848
rect 157444 148730 157472 195842
rect 157524 192976 157576 192982
rect 157524 192918 157576 192924
rect 157536 148918 157564 192918
rect 157628 151570 157656 199446
rect 157720 198626 157748 199650
rect 157812 199306 157840 199702
rect 158226 199764 158254 200124
rect 158174 199736 158254 199764
rect 158122 199718 158174 199724
rect 158028 199679 158084 199688
rect 158318 199628 158346 200124
rect 158410 199764 158438 200124
rect 158502 199918 158530 200124
rect 158490 199912 158542 199918
rect 158490 199854 158542 199860
rect 158594 199850 158622 200124
rect 158686 199918 158714 200124
rect 158674 199912 158726 199918
rect 158674 199854 158726 199860
rect 158582 199844 158634 199850
rect 158582 199786 158634 199792
rect 158778 199764 158806 200124
rect 158410 199753 158484 199764
rect 158410 199744 158498 199753
rect 158410 199736 158442 199744
rect 158686 199736 158806 199764
rect 158686 199696 158714 199736
rect 158442 199679 158498 199688
rect 158640 199668 158714 199696
rect 157982 199608 158038 199617
rect 157892 199572 157944 199578
rect 158272 199600 158346 199628
rect 158444 199640 158496 199646
rect 157982 199543 158038 199552
rect 158076 199572 158128 199578
rect 157892 199514 157944 199520
rect 157800 199300 157852 199306
rect 157800 199242 157852 199248
rect 157798 199064 157854 199073
rect 157798 198999 157800 199008
rect 157852 198999 157854 199008
rect 157800 198970 157852 198976
rect 157708 198620 157760 198626
rect 157708 198562 157760 198568
rect 157708 196716 157760 196722
rect 157708 196658 157760 196664
rect 157720 152794 157748 196658
rect 157904 196625 157932 199514
rect 157890 196616 157946 196625
rect 157890 196551 157946 196560
rect 157996 196314 158024 199543
rect 158076 199514 158128 199520
rect 157984 196308 158036 196314
rect 157984 196250 158036 196256
rect 157800 196240 157852 196246
rect 157800 196182 157852 196188
rect 157812 152862 157840 196182
rect 157984 195968 158036 195974
rect 157984 195910 158036 195916
rect 157996 190454 158024 195910
rect 158088 195906 158116 199514
rect 158076 195900 158128 195906
rect 158076 195842 158128 195848
rect 158272 193214 158300 199600
rect 158444 199582 158496 199588
rect 158536 199640 158588 199646
rect 158536 199582 158588 199588
rect 158456 196246 158484 199582
rect 158444 196240 158496 196246
rect 158444 196182 158496 196188
rect 158548 196081 158576 199582
rect 158640 198257 158668 199668
rect 158870 199560 158898 200124
rect 158962 199730 158990 200124
rect 159054 199850 159082 200124
rect 159042 199844 159094 199850
rect 159042 199786 159094 199792
rect 159146 199764 159174 200124
rect 159238 199918 159266 200124
rect 159330 199918 159358 200124
rect 159422 199918 159450 200124
rect 159514 199923 159542 200124
rect 159226 199912 159278 199918
rect 159226 199854 159278 199860
rect 159318 199912 159370 199918
rect 159318 199854 159370 199860
rect 159410 199912 159462 199918
rect 159410 199854 159462 199860
rect 159500 199914 159556 199923
rect 159606 199918 159634 200124
rect 159698 199918 159726 200124
rect 159500 199849 159556 199858
rect 159594 199912 159646 199918
rect 159594 199854 159646 199860
rect 159686 199912 159738 199918
rect 159686 199854 159738 199860
rect 159272 199776 159324 199782
rect 159146 199736 159220 199764
rect 158962 199702 159036 199730
rect 159008 199617 159036 199702
rect 159088 199640 159140 199646
rect 158824 199532 158898 199560
rect 158994 199608 159050 199617
rect 159088 199582 159140 199588
rect 158994 199543 159050 199552
rect 158720 199300 158772 199306
rect 158720 199242 158772 199248
rect 158626 198248 158682 198257
rect 158626 198183 158682 198192
rect 158534 196072 158590 196081
rect 158534 196007 158590 196016
rect 158732 195362 158760 199242
rect 158824 195566 158852 199532
rect 158994 199472 159050 199481
rect 158994 199407 159050 199416
rect 159008 197266 159036 199407
rect 158996 197260 159048 197266
rect 158996 197202 159048 197208
rect 159100 197112 159128 199582
rect 158916 197084 159128 197112
rect 158812 195560 158864 195566
rect 158812 195502 158864 195508
rect 158810 195392 158866 195401
rect 158720 195356 158772 195362
rect 158810 195327 158866 195336
rect 158720 195298 158772 195304
rect 158272 193186 158392 193214
rect 158364 192982 158392 193186
rect 158352 192976 158404 192982
rect 158352 192918 158404 192924
rect 158628 192092 158680 192098
rect 158628 192034 158680 192040
rect 157996 190426 158116 190454
rect 157800 152856 157852 152862
rect 157800 152798 157852 152804
rect 157708 152788 157760 152794
rect 157708 152730 157760 152736
rect 157616 151564 157668 151570
rect 157616 151506 157668 151512
rect 157524 148912 157576 148918
rect 157524 148854 157576 148860
rect 157444 148702 157564 148730
rect 157352 146934 157472 146962
rect 157340 142180 157392 142186
rect 157340 142122 157392 142128
rect 157352 142089 157380 142122
rect 157338 142080 157394 142089
rect 157338 142015 157394 142024
rect 157154 141400 157210 141409
rect 157154 141335 157210 141344
rect 156788 140072 156840 140078
rect 156788 140014 156840 140020
rect 156248 139862 156676 139890
rect 157168 139754 157196 141335
rect 157444 140146 157472 146934
rect 157536 146062 157564 148702
rect 157890 148608 157946 148617
rect 157890 148543 157946 148552
rect 157524 146056 157576 146062
rect 157524 145998 157576 146004
rect 157800 144424 157852 144430
rect 157800 144366 157852 144372
rect 157812 140162 157840 144366
rect 157432 140140 157484 140146
rect 157432 140082 157484 140088
rect 157766 140134 157840 140162
rect 157766 139876 157794 140134
rect 157904 139890 157932 148543
rect 158088 141506 158116 190426
rect 158640 148442 158668 192034
rect 158824 148986 158852 195327
rect 158916 152998 158944 197084
rect 159088 196988 159140 196994
rect 159088 196930 159140 196936
rect 158996 195900 159048 195906
rect 158996 195842 159048 195848
rect 158904 152992 158956 152998
rect 158904 152934 158956 152940
rect 159008 152930 159036 195842
rect 159100 187406 159128 196930
rect 159192 189922 159220 199736
rect 159272 199718 159324 199724
rect 159790 199730 159818 200124
rect 159882 199923 159910 200124
rect 159868 199914 159924 199923
rect 159868 199849 159924 199858
rect 159974 199764 160002 200124
rect 160066 199850 160094 200124
rect 160158 199918 160186 200124
rect 160146 199912 160198 199918
rect 160146 199854 160198 199860
rect 160054 199844 160106 199850
rect 160054 199786 160106 199792
rect 159928 199736 160002 199764
rect 159284 195906 159312 199718
rect 159364 199708 159416 199714
rect 159364 199650 159416 199656
rect 159640 199708 159692 199714
rect 159790 199702 159864 199730
rect 159640 199650 159692 199656
rect 159272 195900 159324 195906
rect 159272 195842 159324 195848
rect 159376 195294 159404 199650
rect 159548 199640 159600 199646
rect 159548 199582 159600 199588
rect 159456 199572 159508 199578
rect 159456 199514 159508 199520
rect 159468 198014 159496 199514
rect 159560 199374 159588 199582
rect 159548 199368 159600 199374
rect 159548 199310 159600 199316
rect 159546 198520 159602 198529
rect 159546 198455 159548 198464
rect 159600 198455 159602 198464
rect 159548 198426 159600 198432
rect 159456 198008 159508 198014
rect 159456 197950 159508 197956
rect 159548 196308 159600 196314
rect 159548 196250 159600 196256
rect 159364 195288 159416 195294
rect 159364 195230 159416 195236
rect 159560 191834 159588 196250
rect 159652 193214 159680 199650
rect 159732 199640 159784 199646
rect 159732 199582 159784 199588
rect 159744 198422 159772 199582
rect 159732 198416 159784 198422
rect 159732 198358 159784 198364
rect 159836 198218 159864 199702
rect 159824 198212 159876 198218
rect 159824 198154 159876 198160
rect 159928 196994 159956 199736
rect 160250 199696 160278 200124
rect 160342 199923 160370 200124
rect 160328 199914 160384 199923
rect 160328 199849 160384 199858
rect 160434 199730 160462 200124
rect 160526 199923 160554 200124
rect 160512 199914 160568 199923
rect 160618 199918 160646 200124
rect 160710 199918 160738 200124
rect 160802 199923 160830 200124
rect 160512 199849 160568 199858
rect 160606 199912 160658 199918
rect 160606 199854 160658 199860
rect 160698 199912 160750 199918
rect 160698 199854 160750 199860
rect 160788 199914 160844 199923
rect 160788 199849 160844 199858
rect 160894 199850 160922 200124
rect 160986 199850 161014 200124
rect 160882 199844 160934 199850
rect 160882 199786 160934 199792
rect 160974 199844 161026 199850
rect 160974 199786 161026 199792
rect 160020 199668 160278 199696
rect 160388 199702 160462 199730
rect 160834 199744 160890 199753
rect 160560 199708 160612 199714
rect 160020 197198 160048 199668
rect 160282 199608 160338 199617
rect 160192 199572 160244 199578
rect 160112 199532 160192 199560
rect 160008 197192 160060 197198
rect 160008 197134 160060 197140
rect 159916 196988 159968 196994
rect 159916 196930 159968 196936
rect 160112 193214 160140 199532
rect 160282 199543 160338 199552
rect 160192 199514 160244 199520
rect 160192 199436 160244 199442
rect 160192 199378 160244 199384
rect 160204 198966 160232 199378
rect 160192 198960 160244 198966
rect 160192 198902 160244 198908
rect 160296 197810 160324 199543
rect 160284 197804 160336 197810
rect 160284 197746 160336 197752
rect 160388 196976 160416 199702
rect 161078 199730 161106 200124
rect 161170 199918 161198 200124
rect 161262 199918 161290 200124
rect 161354 199923 161382 200124
rect 161158 199912 161210 199918
rect 161158 199854 161210 199860
rect 161250 199912 161302 199918
rect 161250 199854 161302 199860
rect 161340 199914 161396 199923
rect 161446 199918 161474 200124
rect 161538 199918 161566 200124
rect 161630 199923 161658 200124
rect 161340 199849 161396 199858
rect 161434 199912 161486 199918
rect 161434 199854 161486 199860
rect 161526 199912 161578 199918
rect 161526 199854 161578 199860
rect 161616 199914 161672 199923
rect 161722 199918 161750 200124
rect 161814 199918 161842 200124
rect 161906 199918 161934 200124
rect 161616 199849 161672 199858
rect 161710 199912 161762 199918
rect 161710 199854 161762 199860
rect 161802 199912 161854 199918
rect 161802 199854 161854 199860
rect 161894 199912 161946 199918
rect 161894 199854 161946 199860
rect 161204 199776 161256 199782
rect 161202 199744 161204 199753
rect 161478 199778 161534 199787
rect 161256 199744 161258 199753
rect 160834 199679 160890 199688
rect 160928 199708 160980 199714
rect 160560 199650 160612 199656
rect 160466 199608 160522 199617
rect 160466 199543 160522 199552
rect 159652 193186 159956 193214
rect 159560 191806 159680 191834
rect 159652 190454 159680 191806
rect 159652 190426 159772 190454
rect 159180 189916 159232 189922
rect 159180 189858 159232 189864
rect 159088 187400 159140 187406
rect 159088 187342 159140 187348
rect 159744 158166 159772 190426
rect 159732 158160 159784 158166
rect 159732 158102 159784 158108
rect 158996 152924 159048 152930
rect 158996 152866 159048 152872
rect 158812 148980 158864 148986
rect 158812 148922 158864 148928
rect 158628 148436 158680 148442
rect 158628 148378 158680 148384
rect 159928 145994 159956 193186
rect 160020 193186 160140 193214
rect 160204 196948 160416 196976
rect 160020 187474 160048 193186
rect 160008 187468 160060 187474
rect 160008 187410 160060 187416
rect 159916 145988 159968 145994
rect 159916 145930 159968 145936
rect 160204 145790 160232 196948
rect 160376 196852 160428 196858
rect 160376 196794 160428 196800
rect 160284 196716 160336 196722
rect 160284 196658 160336 196664
rect 160296 149054 160324 196658
rect 160388 153202 160416 196794
rect 160480 189582 160508 199543
rect 160572 196858 160600 199650
rect 160744 199640 160796 199646
rect 160744 199582 160796 199588
rect 160652 199572 160704 199578
rect 160652 199514 160704 199520
rect 160664 197305 160692 199514
rect 160756 197742 160784 199582
rect 160744 197736 160796 197742
rect 160744 197678 160796 197684
rect 160650 197296 160706 197305
rect 160848 197266 160876 199679
rect 161078 199702 161152 199730
rect 160928 199650 160980 199656
rect 160650 197231 160706 197240
rect 160836 197260 160888 197266
rect 160836 197202 160888 197208
rect 160652 197192 160704 197198
rect 160652 197134 160704 197140
rect 160560 196852 160612 196858
rect 160560 196794 160612 196800
rect 160664 196704 160692 197134
rect 160940 196722 160968 199650
rect 161018 199608 161074 199617
rect 161018 199543 161074 199552
rect 160572 196676 160692 196704
rect 160928 196716 160980 196722
rect 160572 190194 160600 196676
rect 160928 196658 160980 196664
rect 161032 193214 161060 199543
rect 161124 196761 161152 199702
rect 161202 199679 161258 199688
rect 161388 199708 161440 199714
rect 161478 199713 161534 199722
rect 161664 199776 161716 199782
rect 161664 199718 161716 199724
rect 161756 199776 161808 199782
rect 161756 199718 161808 199724
rect 161388 199650 161440 199656
rect 161204 199572 161256 199578
rect 161400 199560 161428 199650
rect 161480 199640 161532 199646
rect 161480 199582 161532 199588
rect 161572 199640 161624 199646
rect 161572 199582 161624 199588
rect 161204 199514 161256 199520
rect 161308 199532 161428 199560
rect 161110 196752 161166 196761
rect 161110 196687 161166 196696
rect 161216 196636 161244 199514
rect 160664 193186 161060 193214
rect 161124 196608 161244 196636
rect 160664 192098 160692 193186
rect 160652 192092 160704 192098
rect 160652 192034 160704 192040
rect 161124 190454 161152 196608
rect 161202 196480 161258 196489
rect 161202 196415 161258 196424
rect 161216 191214 161244 196415
rect 161308 195906 161336 199532
rect 161388 199436 161440 199442
rect 161388 199378 161440 199384
rect 161400 196722 161428 199378
rect 161388 196716 161440 196722
rect 161388 196658 161440 196664
rect 161296 195900 161348 195906
rect 161296 195842 161348 195848
rect 161492 195401 161520 199582
rect 161584 199481 161612 199582
rect 161570 199472 161626 199481
rect 161570 199407 161626 199416
rect 161676 199322 161704 199718
rect 161584 199294 161704 199322
rect 161584 197946 161612 199294
rect 161664 199232 161716 199238
rect 161664 199174 161716 199180
rect 161676 199102 161704 199174
rect 161664 199096 161716 199102
rect 161664 199038 161716 199044
rect 161572 197940 161624 197946
rect 161572 197882 161624 197888
rect 161768 196178 161796 199718
rect 161848 199708 161900 199714
rect 161998 199696 162026 200124
rect 162090 199923 162118 200124
rect 162076 199914 162132 199923
rect 162182 199918 162210 200124
rect 162274 199923 162302 200124
rect 162076 199849 162132 199858
rect 162170 199912 162222 199918
rect 162170 199854 162222 199860
rect 162260 199914 162316 199923
rect 162366 199918 162394 200124
rect 162458 199918 162486 200124
rect 162550 199918 162578 200124
rect 162642 199918 162670 200124
rect 162260 199849 162316 199858
rect 162354 199912 162406 199918
rect 162354 199854 162406 199860
rect 162446 199912 162498 199918
rect 162446 199854 162498 199860
rect 162538 199912 162590 199918
rect 162538 199854 162590 199860
rect 162630 199912 162682 199918
rect 162630 199854 162682 199860
rect 162308 199776 162360 199782
rect 162214 199744 162270 199753
rect 161848 199650 161900 199656
rect 161952 199668 162026 199696
rect 162124 199708 162176 199714
rect 161756 196172 161808 196178
rect 161756 196114 161808 196120
rect 161754 196072 161810 196081
rect 161754 196007 161810 196016
rect 161664 195968 161716 195974
rect 161664 195910 161716 195916
rect 161570 195800 161626 195809
rect 161570 195735 161626 195744
rect 161478 195392 161534 195401
rect 161478 195327 161534 195336
rect 161204 191208 161256 191214
rect 161204 191150 161256 191156
rect 161124 190426 161336 190454
rect 160560 190188 160612 190194
rect 160560 190130 160612 190136
rect 160468 189576 160520 189582
rect 160468 189518 160520 189524
rect 160376 153196 160428 153202
rect 160376 153138 160428 153144
rect 160284 149048 160336 149054
rect 160284 148990 160336 148996
rect 161308 145926 161336 190426
rect 161584 148850 161612 195735
rect 161676 153134 161704 195910
rect 161664 153128 161716 153134
rect 161664 153070 161716 153076
rect 161768 153066 161796 196007
rect 161860 192710 161888 199650
rect 161952 196858 161980 199668
rect 162308 199718 162360 199724
rect 162400 199776 162452 199782
rect 162400 199718 162452 199724
rect 162214 199679 162270 199688
rect 162124 199650 162176 199656
rect 162032 199368 162084 199374
rect 162032 199310 162084 199316
rect 161940 196852 161992 196858
rect 161940 196794 161992 196800
rect 161940 196376 161992 196382
rect 161940 196318 161992 196324
rect 161848 192704 161900 192710
rect 161848 192646 161900 192652
rect 161848 192432 161900 192438
rect 161848 192374 161900 192380
rect 161860 187542 161888 192374
rect 161848 187536 161900 187542
rect 161848 187478 161900 187484
rect 161952 187338 161980 196318
rect 162044 195673 162072 199310
rect 162030 195664 162086 195673
rect 162030 195599 162086 195608
rect 162136 193118 162164 199650
rect 162228 196761 162256 199679
rect 162214 196752 162270 196761
rect 162214 196687 162270 196696
rect 162124 193112 162176 193118
rect 162124 193054 162176 193060
rect 161940 187332 161992 187338
rect 161940 187274 161992 187280
rect 161756 153060 161808 153066
rect 161756 153002 161808 153008
rect 161572 148844 161624 148850
rect 161572 148786 161624 148792
rect 161296 145920 161348 145926
rect 161296 145862 161348 145868
rect 160192 145784 160244 145790
rect 160192 145726 160244 145732
rect 162320 145722 162348 199718
rect 162412 199617 162440 199718
rect 162584 199708 162636 199714
rect 162734 199696 162762 200124
rect 162826 199764 162854 200124
rect 162918 199923 162946 200124
rect 162904 199914 162960 199923
rect 163010 199918 163038 200124
rect 162904 199849 162960 199858
rect 162998 199912 163050 199918
rect 162998 199854 163050 199860
rect 163102 199764 163130 200124
rect 162826 199736 162900 199764
rect 162584 199650 162636 199656
rect 162688 199668 162762 199696
rect 162398 199608 162454 199617
rect 162398 199543 162454 199552
rect 162400 199504 162452 199510
rect 162400 199446 162452 199452
rect 162412 199209 162440 199446
rect 162492 199368 162544 199374
rect 162492 199310 162544 199316
rect 162398 199200 162454 199209
rect 162398 199135 162454 199144
rect 162504 198694 162532 199310
rect 162492 198688 162544 198694
rect 162492 198630 162544 198636
rect 162490 197840 162546 197849
rect 162490 197775 162546 197784
rect 162398 196888 162454 196897
rect 162398 196823 162454 196832
rect 162412 192438 162440 196823
rect 162504 195634 162532 197775
rect 162492 195628 162544 195634
rect 162492 195570 162544 195576
rect 162596 195537 162624 199650
rect 162688 196382 162716 199668
rect 162872 199458 162900 199736
rect 163056 199736 163130 199764
rect 162950 199608 163006 199617
rect 162950 199543 163006 199552
rect 162780 199430 162900 199458
rect 162780 197198 162808 199430
rect 162768 197192 162820 197198
rect 162768 197134 162820 197140
rect 162768 196716 162820 196722
rect 162768 196658 162820 196664
rect 162676 196376 162728 196382
rect 162676 196318 162728 196324
rect 162582 195528 162638 195537
rect 162582 195463 162638 195472
rect 162676 193112 162728 193118
rect 162676 193054 162728 193060
rect 162400 192432 162452 192438
rect 162400 192374 162452 192380
rect 162688 191486 162716 193054
rect 162676 191480 162728 191486
rect 162676 191422 162728 191428
rect 162780 151434 162808 196658
rect 162964 196450 162992 199543
rect 163056 198286 163084 199736
rect 163194 199628 163222 200124
rect 163286 199918 163314 200124
rect 163378 199918 163406 200124
rect 163470 199923 163498 200124
rect 163274 199912 163326 199918
rect 163274 199854 163326 199860
rect 163366 199912 163418 199918
rect 163366 199854 163418 199860
rect 163456 199914 163512 199923
rect 163456 199849 163512 199858
rect 163274 199776 163326 199782
rect 163562 199764 163590 200124
rect 163654 199787 163682 200124
rect 163516 199753 163590 199764
rect 163274 199718 163326 199724
rect 163502 199744 163590 199753
rect 163286 199646 163314 199718
rect 163558 199736 163590 199744
rect 163640 199778 163696 199787
rect 163640 199713 163696 199722
rect 163502 199679 163558 199688
rect 163746 199696 163774 200124
rect 163838 199850 163866 200124
rect 163930 199918 163958 200124
rect 163918 199912 163970 199918
rect 163918 199854 163970 199860
rect 163826 199844 163878 199850
rect 163826 199786 163878 199792
rect 164022 199730 164050 200124
rect 164114 199923 164142 200124
rect 164100 199914 164156 199923
rect 164100 199849 164156 199858
rect 164206 199764 164234 200124
rect 164298 199918 164326 200124
rect 164390 199923 164418 200124
rect 164286 199912 164338 199918
rect 164286 199854 164338 199860
rect 164376 199914 164432 199923
rect 164376 199849 164432 199858
rect 164160 199736 164234 199764
rect 164332 199776 164384 199782
rect 163872 199708 163924 199714
rect 163746 199668 163820 199696
rect 163148 199600 163222 199628
rect 163274 199640 163326 199646
rect 163044 198280 163096 198286
rect 163044 198222 163096 198228
rect 162952 196444 163004 196450
rect 162952 196386 163004 196392
rect 163148 195514 163176 199600
rect 163274 199582 163326 199588
rect 163412 199640 163464 199646
rect 163412 199582 163464 199588
rect 163228 199504 163280 199510
rect 163228 199446 163280 199452
rect 163240 198966 163268 199446
rect 163320 199436 163372 199442
rect 163320 199378 163372 199384
rect 163228 198960 163280 198966
rect 163228 198902 163280 198908
rect 163332 196840 163360 199378
rect 163424 198150 163452 199582
rect 163688 199572 163740 199578
rect 163688 199514 163740 199520
rect 163700 199481 163728 199514
rect 163686 199472 163742 199481
rect 163596 199436 163648 199442
rect 163686 199407 163742 199416
rect 163596 199378 163648 199384
rect 163608 199073 163636 199378
rect 163686 199336 163742 199345
rect 163686 199271 163688 199280
rect 163740 199271 163742 199280
rect 163688 199242 163740 199248
rect 163594 199064 163650 199073
rect 163594 198999 163650 199008
rect 163412 198144 163464 198150
rect 163412 198086 163464 198092
rect 163594 196888 163650 196897
rect 163332 196812 163544 196840
rect 163594 196823 163650 196832
rect 163318 196480 163374 196489
rect 163228 196444 163280 196450
rect 163318 196415 163374 196424
rect 163228 196386 163280 196392
rect 162964 195486 163176 195514
rect 162768 151428 162820 151434
rect 162768 151370 162820 151376
rect 162308 145716 162360 145722
rect 162308 145658 162360 145664
rect 162490 144392 162546 144401
rect 159548 144356 159600 144362
rect 162490 144327 162546 144336
rect 159548 144298 159600 144304
rect 159180 142180 159232 142186
rect 159180 142122 159232 142128
rect 158076 141500 158128 141506
rect 158076 141442 158128 141448
rect 159192 139890 159220 142122
rect 159560 139890 159588 144298
rect 160834 144120 160890 144129
rect 160834 144055 160890 144064
rect 159638 142896 159694 142905
rect 159638 142831 159694 142840
rect 157904 139862 158332 139890
rect 158884 139862 159220 139890
rect 159436 139862 159588 139890
rect 159652 139890 159680 142831
rect 160848 139890 160876 144055
rect 161938 142760 161994 142769
rect 161938 142695 161994 142704
rect 161952 139890 161980 142695
rect 162504 139890 162532 144327
rect 162964 140214 162992 195486
rect 163136 195220 163188 195226
rect 163136 195162 163188 195168
rect 163044 195152 163096 195158
rect 163044 195094 163096 195100
rect 163056 145625 163084 195094
rect 163148 148714 163176 195162
rect 163240 148782 163268 196386
rect 163332 151366 163360 196415
rect 163410 196344 163466 196353
rect 163410 196279 163466 196288
rect 163320 151360 163372 151366
rect 163320 151302 163372 151308
rect 163424 151298 163452 196279
rect 163516 189990 163544 196812
rect 163608 191418 163636 196823
rect 163792 195158 163820 199668
rect 164022 199702 164096 199730
rect 163872 199650 163924 199656
rect 163780 195152 163832 195158
rect 163780 195094 163832 195100
rect 163884 193214 163912 199650
rect 163962 199608 164018 199617
rect 163962 199543 163964 199552
rect 164016 199543 164018 199552
rect 163964 199514 164016 199520
rect 163964 199436 164016 199442
rect 163964 199378 164016 199384
rect 163976 199345 164004 199378
rect 163962 199336 164018 199345
rect 163962 199271 164018 199280
rect 163964 199164 164016 199170
rect 163964 199106 164016 199112
rect 163976 198830 164004 199106
rect 163964 198824 164016 198830
rect 163964 198766 164016 198772
rect 164068 195226 164096 199702
rect 164160 196897 164188 199736
rect 164482 199764 164510 200124
rect 164574 199918 164602 200124
rect 164562 199912 164614 199918
rect 164562 199854 164614 199860
rect 164666 199764 164694 200124
rect 164482 199736 164556 199764
rect 164620 199753 164694 199764
rect 164332 199718 164384 199724
rect 164240 199640 164292 199646
rect 164240 199582 164292 199588
rect 164252 197169 164280 199582
rect 164344 199209 164372 199718
rect 164424 199640 164476 199646
rect 164528 199617 164556 199736
rect 164606 199744 164694 199753
rect 164662 199736 164694 199744
rect 164606 199679 164662 199688
rect 164424 199582 164476 199588
rect 164514 199608 164570 199617
rect 164330 199200 164386 199209
rect 164330 199135 164386 199144
rect 164330 197568 164386 197577
rect 164330 197503 164386 197512
rect 164238 197160 164294 197169
rect 164238 197095 164294 197104
rect 164146 196888 164202 196897
rect 164344 196874 164372 197503
rect 164436 196994 164464 199582
rect 164758 199594 164786 200124
rect 164850 199850 164878 200124
rect 164942 199850 164970 200124
rect 165034 199850 165062 200124
rect 164838 199844 164890 199850
rect 164838 199786 164890 199792
rect 164930 199844 164982 199850
rect 164930 199786 164982 199792
rect 165022 199844 165074 199850
rect 165022 199786 165074 199792
rect 165126 199764 165154 200124
rect 165218 199923 165246 200124
rect 165204 199914 165260 199923
rect 165204 199849 165260 199858
rect 165310 199850 165338 200124
rect 165298 199844 165350 199850
rect 165298 199786 165350 199792
rect 165126 199753 165200 199764
rect 164882 199744 164938 199753
rect 165126 199744 165214 199753
rect 165126 199736 165158 199744
rect 164882 199679 164938 199688
rect 165158 199679 165214 199688
rect 164514 199543 164570 199552
rect 164608 199572 164660 199578
rect 164608 199514 164660 199520
rect 164712 199566 164786 199594
rect 164516 199504 164568 199510
rect 164516 199446 164568 199452
rect 164528 198694 164556 199446
rect 164620 199073 164648 199514
rect 164606 199064 164662 199073
rect 164606 198999 164662 199008
rect 164516 198688 164568 198694
rect 164516 198630 164568 198636
rect 164712 197130 164740 199566
rect 164792 199504 164844 199510
rect 164792 199446 164844 199452
rect 164700 197124 164752 197130
rect 164700 197066 164752 197072
rect 164424 196988 164476 196994
rect 164424 196930 164476 196936
rect 164804 196874 164832 199446
rect 164146 196823 164202 196832
rect 164252 196846 164372 196874
rect 164436 196846 164832 196874
rect 164056 195220 164108 195226
rect 164056 195162 164108 195168
rect 163884 193186 164096 193214
rect 164068 191834 164096 193186
rect 164068 191806 164188 191834
rect 164160 191554 164188 191806
rect 164148 191548 164200 191554
rect 164148 191490 164200 191496
rect 163596 191412 163648 191418
rect 163596 191354 163648 191360
rect 164148 191412 164200 191418
rect 164148 191354 164200 191360
rect 163504 189984 163556 189990
rect 163504 189926 163556 189932
rect 163412 151292 163464 151298
rect 163412 151234 163464 151240
rect 163228 148776 163280 148782
rect 163228 148718 163280 148724
rect 163136 148708 163188 148714
rect 163136 148650 163188 148656
rect 163042 145616 163098 145625
rect 163042 145551 163098 145560
rect 163964 144560 164016 144566
rect 163964 144502 164016 144508
rect 163594 142896 163650 142905
rect 163594 142831 163650 142840
rect 162952 140208 163004 140214
rect 162952 140150 163004 140156
rect 159652 139862 159988 139890
rect 160540 139862 160876 139890
rect 161644 139862 161980 139890
rect 162196 139862 162532 139890
rect 162582 139904 162638 139913
rect 163608 139890 163636 142831
rect 163976 139890 164004 144502
rect 164160 140282 164188 191354
rect 164252 141642 164280 196846
rect 164332 196784 164384 196790
rect 164332 196726 164384 196732
rect 164344 144673 164372 196726
rect 164436 148510 164464 196846
rect 164516 196716 164568 196722
rect 164896 196704 164924 199679
rect 165160 199640 165212 199646
rect 165402 199628 165430 200124
rect 165494 199730 165522 200124
rect 165586 199923 165614 200124
rect 165572 199914 165628 199923
rect 165572 199849 165628 199858
rect 165678 199782 165706 200124
rect 165666 199776 165718 199782
rect 165494 199702 165568 199730
rect 165770 199753 165798 200124
rect 165666 199718 165718 199724
rect 165756 199744 165812 199753
rect 165402 199600 165476 199628
rect 165160 199582 165212 199588
rect 164976 199504 165028 199510
rect 164976 199446 165028 199452
rect 164516 196658 164568 196664
rect 164620 196676 164924 196704
rect 164424 148504 164476 148510
rect 164424 148446 164476 148452
rect 164528 148306 164556 196658
rect 164620 148646 164648 196676
rect 164884 196512 164936 196518
rect 164988 196489 165016 199446
rect 165172 197305 165200 199582
rect 165344 199504 165396 199510
rect 165250 199472 165306 199481
rect 165344 199446 165396 199452
rect 165250 199407 165306 199416
rect 165158 197296 165214 197305
rect 165158 197231 165214 197240
rect 164884 196454 164936 196460
rect 164974 196480 165030 196489
rect 164896 191834 164924 196454
rect 164974 196415 165030 196424
rect 165264 194954 165292 199407
rect 165356 199034 165384 199446
rect 165344 199028 165396 199034
rect 165344 198970 165396 198976
rect 165448 198734 165476 199600
rect 165356 198706 165476 198734
rect 165356 196790 165384 198706
rect 165540 198642 165568 199702
rect 165756 199679 165812 199688
rect 165620 199640 165672 199646
rect 165620 199582 165672 199588
rect 165448 198614 165568 198642
rect 165344 196784 165396 196790
rect 165344 196726 165396 196732
rect 165448 196518 165476 198614
rect 165528 198552 165580 198558
rect 165528 198494 165580 198500
rect 165436 196512 165488 196518
rect 165436 196454 165488 196460
rect 165252 194948 165304 194954
rect 165252 194890 165304 194896
rect 164712 191806 164924 191834
rect 164712 190058 164740 191806
rect 164700 190052 164752 190058
rect 164700 189994 164752 190000
rect 165540 180794 165568 198494
rect 165632 196722 165660 199582
rect 165712 199572 165764 199578
rect 165712 199514 165764 199520
rect 165724 198354 165752 199514
rect 165862 199492 165890 200124
rect 165954 199628 165982 200124
rect 166046 199923 166074 200124
rect 166032 199914 166088 199923
rect 166032 199849 166088 199858
rect 166138 199730 166166 200124
rect 166092 199702 166166 199730
rect 165954 199600 166028 199628
rect 165862 199481 165936 199492
rect 165862 199472 165950 199481
rect 165862 199464 165894 199472
rect 165894 199407 165950 199416
rect 165712 198348 165764 198354
rect 165712 198290 165764 198296
rect 165620 196716 165672 196722
rect 165620 196658 165672 196664
rect 165712 196716 165764 196722
rect 165712 196658 165764 196664
rect 165264 180766 165568 180794
rect 165264 152386 165292 180766
rect 165724 152454 165752 196658
rect 166000 196654 166028 199600
rect 166092 199345 166120 199702
rect 166230 199628 166258 200124
rect 166322 199923 166350 200124
rect 166308 199914 166364 199923
rect 166414 199918 166442 200124
rect 166506 199918 166534 200124
rect 166598 199918 166626 200124
rect 166690 199918 166718 200124
rect 166782 199918 166810 200124
rect 166308 199849 166364 199858
rect 166402 199912 166454 199918
rect 166402 199854 166454 199860
rect 166494 199912 166546 199918
rect 166494 199854 166546 199860
rect 166586 199912 166638 199918
rect 166586 199854 166638 199860
rect 166678 199912 166730 199918
rect 166678 199854 166730 199860
rect 166770 199912 166822 199918
rect 166770 199854 166822 199860
rect 166356 199776 166408 199782
rect 166356 199718 166408 199724
rect 166540 199776 166592 199782
rect 166874 199730 166902 200124
rect 166966 199753 166994 200124
rect 167058 199918 167086 200124
rect 167150 199923 167178 200124
rect 167046 199912 167098 199918
rect 167046 199854 167098 199860
rect 167136 199914 167192 199923
rect 167136 199849 167192 199858
rect 166540 199718 166592 199724
rect 166184 199600 166258 199628
rect 166078 199336 166134 199345
rect 166078 199271 166134 199280
rect 165988 196648 166040 196654
rect 165988 196590 166040 196596
rect 166184 196500 166212 199600
rect 166264 199504 166316 199510
rect 166264 199446 166316 199452
rect 166276 198937 166304 199446
rect 166262 198928 166318 198937
rect 166262 198863 166318 198872
rect 166264 198484 166316 198490
rect 166264 198426 166316 198432
rect 165908 196472 166212 196500
rect 165908 155582 165936 196472
rect 166078 196344 166134 196353
rect 166078 196279 166134 196288
rect 165988 195152 166040 195158
rect 165988 195094 166040 195100
rect 166000 155650 166028 195094
rect 166092 187610 166120 196279
rect 166276 195974 166304 198426
rect 166368 197334 166396 199718
rect 166448 199708 166500 199714
rect 166448 199650 166500 199656
rect 166356 197328 166408 197334
rect 166356 197270 166408 197276
rect 166276 195946 166396 195974
rect 166262 195800 166318 195809
rect 166262 195735 166318 195744
rect 166276 191622 166304 195735
rect 166264 191616 166316 191622
rect 166264 191558 166316 191564
rect 166368 190454 166396 195946
rect 166460 195158 166488 199650
rect 166448 195152 166500 195158
rect 166448 195094 166500 195100
rect 166552 193214 166580 199718
rect 166632 199708 166684 199714
rect 166632 199650 166684 199656
rect 166828 199702 166902 199730
rect 166952 199744 167008 199753
rect 166644 197033 166672 199650
rect 166724 199572 166776 199578
rect 166724 199514 166776 199520
rect 166630 197024 166686 197033
rect 166630 196959 166686 196968
rect 166736 196722 166764 199514
rect 166724 196716 166776 196722
rect 166724 196658 166776 196664
rect 166828 193866 166856 199702
rect 167242 199730 167270 200124
rect 167334 199850 167362 200124
rect 167322 199844 167374 199850
rect 167322 199786 167374 199792
rect 166952 199679 167008 199688
rect 167196 199702 167270 199730
rect 166908 199640 166960 199646
rect 166908 199582 166960 199588
rect 166920 198801 166948 199582
rect 167090 199472 167146 199481
rect 167090 199407 167146 199416
rect 166906 198792 166962 198801
rect 166906 198727 166962 198736
rect 167104 198626 167132 199407
rect 167092 198620 167144 198626
rect 167092 198562 167144 198568
rect 167092 198348 167144 198354
rect 167092 198290 167144 198296
rect 167000 196716 167052 196722
rect 167000 196658 167052 196664
rect 166908 196648 166960 196654
rect 166908 196590 166960 196596
rect 166816 193860 166868 193866
rect 166816 193802 166868 193808
rect 166552 193186 166672 193214
rect 166644 190454 166672 193186
rect 166368 190426 166488 190454
rect 166644 190426 166764 190454
rect 166080 187604 166132 187610
rect 166080 187546 166132 187552
rect 166080 158228 166132 158234
rect 166080 158170 166132 158176
rect 165988 155644 166040 155650
rect 165988 155586 166040 155592
rect 165896 155576 165948 155582
rect 165896 155518 165948 155524
rect 165712 152448 165764 152454
rect 165712 152390 165764 152396
rect 165252 152380 165304 152386
rect 165252 152322 165304 152328
rect 164608 148640 164660 148646
rect 164608 148582 164660 148588
rect 164516 148300 164568 148306
rect 164516 148242 164568 148248
rect 164330 144664 164386 144673
rect 164330 144599 164386 144608
rect 165528 144628 165580 144634
rect 165528 144570 165580 144576
rect 165250 143032 165306 143041
rect 165250 142967 165306 142976
rect 164240 141636 164292 141642
rect 164240 141578 164292 141584
rect 164148 140276 164200 140282
rect 164148 140218 164200 140224
rect 165264 139890 165292 142967
rect 165540 140162 165568 144570
rect 166092 140162 166120 158170
rect 166460 141506 166488 190426
rect 166632 143064 166684 143070
rect 166632 143006 166684 143012
rect 166448 141500 166500 141506
rect 166448 141442 166500 141448
rect 166644 140162 166672 143006
rect 162638 139862 162748 139890
rect 163300 139862 163636 139890
rect 163852 139862 164004 139890
rect 164956 139862 165292 139890
rect 165494 140134 165568 140162
rect 166046 140134 166120 140162
rect 166598 140134 166672 140162
rect 165494 139876 165522 140134
rect 166046 139876 166074 140134
rect 166598 139876 166626 140134
rect 162582 139839 162638 139848
rect 164606 139768 164662 139777
rect 157168 139726 157228 139754
rect 164404 139726 164606 139754
rect 164606 139703 164662 139712
rect 161296 139664 161348 139670
rect 161092 139612 161296 139618
rect 161092 139606 161348 139612
rect 161092 139590 161336 139606
rect 166736 139369 166764 190426
rect 166920 152590 166948 196590
rect 166908 152584 166960 152590
rect 166908 152526 166960 152532
rect 167012 148481 167040 196658
rect 167104 149569 167132 198290
rect 167196 197606 167224 199702
rect 167426 199696 167454 200124
rect 167518 199918 167546 200124
rect 167610 199918 167638 200124
rect 167506 199912 167558 199918
rect 167506 199854 167558 199860
rect 167598 199912 167650 199918
rect 167598 199854 167650 199860
rect 167552 199708 167604 199714
rect 167426 199668 167500 199696
rect 167276 199640 167328 199646
rect 167276 199582 167328 199588
rect 167184 197600 167236 197606
rect 167184 197542 167236 197548
rect 167184 194880 167236 194886
rect 167184 194822 167236 194828
rect 167196 151473 167224 194822
rect 167288 155786 167316 199582
rect 167368 199572 167420 199578
rect 167368 199514 167420 199520
rect 167276 155780 167328 155786
rect 167276 155722 167328 155728
rect 167380 155514 167408 199514
rect 167472 191350 167500 199668
rect 167702 199696 167730 200124
rect 167794 199714 167822 200124
rect 167886 199923 167914 200124
rect 167872 199914 167928 199923
rect 167872 199849 167928 199858
rect 167978 199764 168006 200124
rect 168070 199923 168098 200124
rect 168056 199914 168112 199923
rect 168162 199918 168190 200124
rect 168254 199918 168282 200124
rect 168346 199923 168374 200124
rect 168056 199849 168112 199858
rect 168150 199912 168202 199918
rect 168150 199854 168202 199860
rect 168242 199912 168294 199918
rect 168242 199854 168294 199860
rect 168332 199914 168388 199923
rect 168332 199849 168388 199858
rect 167932 199736 168006 199764
rect 167552 199650 167604 199656
rect 167656 199668 167730 199696
rect 167782 199708 167834 199714
rect 167460 191344 167512 191350
rect 167460 191286 167512 191292
rect 167564 155718 167592 199650
rect 167656 196654 167684 199668
rect 167782 199650 167834 199656
rect 167826 199608 167882 199617
rect 167736 199572 167788 199578
rect 167826 199543 167882 199552
rect 167736 199514 167788 199520
rect 167644 196648 167696 196654
rect 167644 196590 167696 196596
rect 167642 196208 167698 196217
rect 167642 196143 167698 196152
rect 167656 191418 167684 196143
rect 167748 194585 167776 199514
rect 167840 197470 167868 199543
rect 167828 197464 167880 197470
rect 167828 197406 167880 197412
rect 167932 197282 167960 199736
rect 168438 199714 168466 200124
rect 168530 199782 168558 200124
rect 168518 199776 168570 199782
rect 168622 199753 168650 200124
rect 168714 199764 168742 200124
rect 168806 199918 168834 200124
rect 168898 199918 168926 200124
rect 168990 199923 169018 200124
rect 168794 199912 168846 199918
rect 168794 199854 168846 199860
rect 168886 199912 168938 199918
rect 168886 199854 168938 199860
rect 168976 199914 169032 199923
rect 168976 199849 169032 199858
rect 169082 199850 169110 200124
rect 169174 199923 169202 200124
rect 169160 199914 169216 199923
rect 169070 199844 169122 199850
rect 169160 199849 169216 199858
rect 169266 199850 169294 200124
rect 169070 199786 169122 199792
rect 169254 199844 169306 199850
rect 169254 199786 169306 199792
rect 168932 199776 168984 199782
rect 168714 199753 168788 199764
rect 168518 199718 168570 199724
rect 168608 199744 168664 199753
rect 168196 199708 168248 199714
rect 168196 199650 168248 199656
rect 168426 199708 168478 199714
rect 168714 199744 168802 199753
rect 168714 199736 168746 199744
rect 168608 199679 168664 199688
rect 169358 199730 169386 200124
rect 169450 199850 169478 200124
rect 169542 199850 169570 200124
rect 169438 199844 169490 199850
rect 169438 199786 169490 199792
rect 169530 199844 169582 199850
rect 169530 199786 169582 199792
rect 169634 199764 169662 200124
rect 169726 199923 169754 200124
rect 169712 199914 169768 199923
rect 169712 199849 169768 199858
rect 169634 199753 169754 199764
rect 169634 199744 169768 199753
rect 169634 199736 169712 199744
rect 168932 199718 168984 199724
rect 168746 199679 168802 199688
rect 168840 199708 168892 199714
rect 168426 199650 168478 199656
rect 168840 199650 168892 199656
rect 168104 199640 168156 199646
rect 168010 199608 168066 199617
rect 168104 199582 168156 199588
rect 168010 199543 168066 199552
rect 167840 197254 167960 197282
rect 167840 194886 167868 197254
rect 167920 197192 167972 197198
rect 167920 197134 167972 197140
rect 167932 195809 167960 197134
rect 167918 195800 167974 195809
rect 167918 195735 167974 195744
rect 167828 194880 167880 194886
rect 167828 194822 167880 194828
rect 167734 194576 167790 194585
rect 167734 194511 167790 194520
rect 168024 193225 168052 199543
rect 168116 198354 168144 199582
rect 168104 198348 168156 198354
rect 168104 198290 168156 198296
rect 168104 198144 168156 198150
rect 168104 198086 168156 198092
rect 168116 197198 168144 198086
rect 168104 197192 168156 197198
rect 168104 197134 168156 197140
rect 168208 196722 168236 199650
rect 168564 199640 168616 199646
rect 168470 199608 168526 199617
rect 168288 199572 168340 199578
rect 168288 199514 168340 199520
rect 168380 199572 168432 199578
rect 168564 199582 168616 199588
rect 168656 199640 168708 199646
rect 168656 199582 168708 199588
rect 168746 199608 168802 199617
rect 168470 199543 168526 199552
rect 168380 199514 168432 199520
rect 168300 198966 168328 199514
rect 168288 198960 168340 198966
rect 168288 198902 168340 198908
rect 168392 198393 168420 199514
rect 168484 199510 168512 199543
rect 168472 199504 168524 199510
rect 168472 199446 168524 199452
rect 168472 199028 168524 199034
rect 168472 198970 168524 198976
rect 168484 198830 168512 198970
rect 168472 198824 168524 198830
rect 168472 198766 168524 198772
rect 168378 198384 168434 198393
rect 168378 198319 168434 198328
rect 168380 197464 168432 197470
rect 168380 197406 168432 197412
rect 168196 196716 168248 196722
rect 168196 196658 168248 196664
rect 168286 196480 168342 196489
rect 168286 196415 168342 196424
rect 168010 193216 168066 193225
rect 168010 193151 168066 193160
rect 167644 191412 167696 191418
rect 167644 191354 167696 191360
rect 167552 155712 167604 155718
rect 167552 155654 167604 155660
rect 167368 155508 167420 155514
rect 167368 155450 167420 155456
rect 168300 155242 168328 196415
rect 168392 192273 168420 197406
rect 168472 196716 168524 196722
rect 168576 196704 168604 199582
rect 168668 199481 168696 199582
rect 168746 199543 168802 199552
rect 168654 199472 168710 199481
rect 168654 199407 168710 199416
rect 168654 199336 168710 199345
rect 168654 199271 168710 199280
rect 168668 199034 168696 199271
rect 168656 199028 168708 199034
rect 168656 198970 168708 198976
rect 168576 196676 168696 196704
rect 168472 196658 168524 196664
rect 168378 192264 168434 192273
rect 168378 192199 168434 192208
rect 168380 192160 168432 192166
rect 168380 192102 168432 192108
rect 168288 155236 168340 155242
rect 168288 155178 168340 155184
rect 167182 151464 167238 151473
rect 167182 151399 167238 151408
rect 167090 149560 167146 149569
rect 167090 149495 167146 149504
rect 166998 148472 167054 148481
rect 166998 148407 167054 148416
rect 168010 144528 168066 144537
rect 168010 144463 168066 144472
rect 167460 141568 167512 141574
rect 167460 141510 167512 141516
rect 167472 139890 167500 141510
rect 168024 139890 168052 144463
rect 168196 143132 168248 143138
rect 168196 143074 168248 143080
rect 167164 139862 167500 139890
rect 167716 139862 168052 139890
rect 168208 139890 168236 143074
rect 168392 142934 168420 192102
rect 168484 151638 168512 196658
rect 168564 196172 168616 196178
rect 168564 196114 168616 196120
rect 168576 191185 168604 196114
rect 168668 191282 168696 196676
rect 168760 193361 168788 199543
rect 168852 198490 168880 199650
rect 168840 198484 168892 198490
rect 168840 198426 168892 198432
rect 168840 198280 168892 198286
rect 168840 198222 168892 198228
rect 168852 195265 168880 198222
rect 168838 195256 168894 195265
rect 168944 195226 168972 199718
rect 169024 199708 169076 199714
rect 169024 199650 169076 199656
rect 169312 199702 169386 199730
rect 169036 196450 169064 199650
rect 169116 199640 169168 199646
rect 169114 199608 169116 199617
rect 169168 199608 169170 199617
rect 169114 199543 169170 199552
rect 169116 199504 169168 199510
rect 169116 199446 169168 199452
rect 169128 196489 169156 199446
rect 169208 199436 169260 199442
rect 169208 199378 169260 199384
rect 169220 199345 169248 199378
rect 169206 199336 169262 199345
rect 169206 199271 169262 199280
rect 169312 196722 169340 199702
rect 169712 199679 169768 199688
rect 169392 199640 169444 199646
rect 169392 199582 169444 199588
rect 169484 199640 169536 199646
rect 169484 199582 169536 199588
rect 169666 199608 169722 199617
rect 169300 196716 169352 196722
rect 169300 196658 169352 196664
rect 169114 196480 169170 196489
rect 169024 196444 169076 196450
rect 169114 196415 169170 196424
rect 169024 196386 169076 196392
rect 169404 196382 169432 199582
rect 169392 196376 169444 196382
rect 169022 196344 169078 196353
rect 169392 196318 169444 196324
rect 169022 196279 169078 196288
rect 168838 195191 168894 195200
rect 168932 195220 168984 195226
rect 168932 195162 168984 195168
rect 168746 193352 168802 193361
rect 168746 193287 168802 193296
rect 169036 191834 169064 196279
rect 169390 196072 169446 196081
rect 169390 196007 169446 196016
rect 169404 195974 169432 196007
rect 169392 195968 169444 195974
rect 169392 195910 169444 195916
rect 168944 191806 169064 191834
rect 168656 191276 168708 191282
rect 168656 191218 168708 191224
rect 168562 191176 168618 191185
rect 168562 191111 168618 191120
rect 168944 191026 168972 191806
rect 168576 190998 168972 191026
rect 168576 155378 168604 190998
rect 169496 180794 169524 199582
rect 169576 199572 169628 199578
rect 169818 199594 169846 200124
rect 169910 199923 169938 200124
rect 169896 199914 169952 199923
rect 169896 199849 169952 199858
rect 170002 199628 170030 200124
rect 170094 199923 170122 200124
rect 170080 199914 170136 199923
rect 170080 199849 170136 199858
rect 170186 199850 170214 200124
rect 170278 199923 170306 200124
rect 170264 199914 170320 199923
rect 170174 199844 170226 199850
rect 170264 199849 170320 199858
rect 170174 199786 170226 199792
rect 170370 199764 170398 200124
rect 170462 199850 170490 200124
rect 170450 199844 170502 199850
rect 170450 199786 170502 199792
rect 170324 199736 170398 199764
rect 170220 199708 170272 199714
rect 170220 199650 170272 199656
rect 170002 199600 170076 199628
rect 169818 199566 169892 199594
rect 169666 199543 169722 199552
rect 169576 199514 169628 199520
rect 169588 196722 169616 199514
rect 169576 196716 169628 196722
rect 169576 196658 169628 196664
rect 169574 196480 169630 196489
rect 169574 196415 169630 196424
rect 169588 191834 169616 196415
rect 169680 192166 169708 199543
rect 169760 199436 169812 199442
rect 169760 199378 169812 199384
rect 169772 199073 169800 199378
rect 169758 199064 169814 199073
rect 169758 198999 169814 199008
rect 169864 199016 169892 199566
rect 169944 199504 169996 199510
rect 169942 199472 169944 199481
rect 169996 199472 169998 199481
rect 169942 199407 169998 199416
rect 169864 198988 169984 199016
rect 169760 197804 169812 197810
rect 169760 197746 169812 197752
rect 169772 197538 169800 197746
rect 169760 197532 169812 197538
rect 169760 197474 169812 197480
rect 169852 196716 169904 196722
rect 169852 196658 169904 196664
rect 169864 196518 169892 196658
rect 169852 196512 169904 196518
rect 169852 196454 169904 196460
rect 169850 196344 169906 196353
rect 169850 196279 169906 196288
rect 169758 196208 169814 196217
rect 169758 196143 169814 196152
rect 169772 193089 169800 196143
rect 169758 193080 169814 193089
rect 169758 193015 169814 193024
rect 169668 192160 169720 192166
rect 169668 192102 169720 192108
rect 169588 191806 169800 191834
rect 168668 180766 169524 180794
rect 168564 155372 168616 155378
rect 168564 155314 168616 155320
rect 168668 155310 168696 180766
rect 168748 158432 168800 158438
rect 168748 158374 168800 158380
rect 168656 155304 168708 155310
rect 168656 155246 168708 155252
rect 168472 151632 168524 151638
rect 168472 151574 168524 151580
rect 168380 142928 168432 142934
rect 168380 142870 168432 142876
rect 168760 139890 168788 158374
rect 169668 143268 169720 143274
rect 169668 143210 169720 143216
rect 169680 139890 169708 143210
rect 169772 140049 169800 191806
rect 169864 147626 169892 196279
rect 169852 147620 169904 147626
rect 169852 147562 169904 147568
rect 169956 147393 169984 198988
rect 170048 198150 170076 199600
rect 170126 199608 170182 199617
rect 170126 199543 170182 199552
rect 170036 198144 170088 198150
rect 170036 198086 170088 198092
rect 170140 196654 170168 199543
rect 170232 198626 170260 199650
rect 170220 198620 170272 198626
rect 170220 198562 170272 198568
rect 170036 196648 170088 196654
rect 170036 196590 170088 196596
rect 170128 196648 170180 196654
rect 170128 196590 170180 196596
rect 170048 192137 170076 196590
rect 170220 196512 170272 196518
rect 170220 196454 170272 196460
rect 170126 196208 170182 196217
rect 170126 196143 170182 196152
rect 170034 192128 170090 192137
rect 170034 192063 170090 192072
rect 170036 158296 170088 158302
rect 170036 158238 170088 158244
rect 169942 147384 169998 147393
rect 169942 147319 169998 147328
rect 170048 143546 170076 158238
rect 170140 147257 170168 196143
rect 170232 192710 170260 196454
rect 170220 192704 170272 192710
rect 170220 192646 170272 192652
rect 170220 155848 170272 155854
rect 170220 155790 170272 155796
rect 170126 147248 170182 147257
rect 170126 147183 170182 147192
rect 170036 143540 170088 143546
rect 170036 143482 170088 143488
rect 169758 140040 169814 140049
rect 169758 139975 169814 139984
rect 170232 139890 170260 155790
rect 170324 147665 170352 199736
rect 170554 199628 170582 200124
rect 170646 199923 170674 200124
rect 170632 199914 170688 199923
rect 170632 199849 170688 199858
rect 170738 199782 170766 200124
rect 170830 199850 170858 200124
rect 170922 199855 170950 200124
rect 171014 199918 171042 200124
rect 171106 199918 171134 200124
rect 171002 199912 171054 199918
rect 170818 199844 170870 199850
rect 170818 199786 170870 199792
rect 170908 199846 170964 199855
rect 171002 199854 171054 199860
rect 171094 199912 171146 199918
rect 171094 199854 171146 199860
rect 170726 199776 170778 199782
rect 170908 199781 170964 199790
rect 171198 199764 171226 200124
rect 171290 199923 171318 200124
rect 171276 199914 171332 199923
rect 171276 199849 171332 199858
rect 171198 199753 171272 199764
rect 171198 199744 171286 199753
rect 171198 199736 171230 199744
rect 170726 199718 170778 199724
rect 171048 199708 171100 199714
rect 171382 199696 171410 200124
rect 171474 199918 171502 200124
rect 171566 199918 171594 200124
rect 171462 199912 171514 199918
rect 171462 199854 171514 199860
rect 171554 199912 171606 199918
rect 171554 199854 171606 199860
rect 171658 199764 171686 200124
rect 171750 199850 171778 200124
rect 171738 199844 171790 199850
rect 171738 199786 171790 199792
rect 171230 199679 171286 199688
rect 171048 199650 171100 199656
rect 171336 199668 171410 199696
rect 171566 199736 171686 199764
rect 171566 199696 171594 199736
rect 171842 199730 171870 200124
rect 171934 199923 171962 200124
rect 171920 199914 171976 199923
rect 172026 199918 172054 200124
rect 171920 199849 171976 199858
rect 172014 199912 172066 199918
rect 172014 199854 172066 199860
rect 172118 199764 172146 200124
rect 172072 199753 172146 199764
rect 172210 199753 172238 200124
rect 172302 199764 172330 200124
rect 172394 199918 172422 200124
rect 172382 199912 172434 199918
rect 172382 199854 172434 199860
rect 172382 199776 172434 199782
rect 171796 199702 171870 199730
rect 172058 199744 172146 199753
rect 171566 199668 171640 199696
rect 170554 199600 170628 199628
rect 170404 199572 170456 199578
rect 170404 199514 170456 199520
rect 170416 198098 170444 199514
rect 170496 199504 170548 199510
rect 170496 199446 170548 199452
rect 170508 198286 170536 199446
rect 170496 198280 170548 198286
rect 170600 198257 170628 199600
rect 170678 199608 170734 199617
rect 170678 199543 170734 199552
rect 170772 199572 170824 199578
rect 170692 198694 170720 199543
rect 170772 199514 170824 199520
rect 170680 198688 170732 198694
rect 170680 198630 170732 198636
rect 170496 198222 170548 198228
rect 170586 198248 170642 198257
rect 170586 198183 170642 198192
rect 170416 198070 170720 198098
rect 170496 198008 170548 198014
rect 170496 197950 170548 197956
rect 170310 147656 170366 147665
rect 170310 147591 170366 147600
rect 170312 143540 170364 143546
rect 170312 143482 170364 143488
rect 168208 139862 168268 139890
rect 168760 139862 168820 139890
rect 169372 139862 169708 139890
rect 169924 139862 170260 139890
rect 170324 139890 170352 143482
rect 170508 141778 170536 197950
rect 170692 192030 170720 198070
rect 170784 192914 170812 199514
rect 170954 199472 171010 199481
rect 170954 199407 171010 199416
rect 170864 198688 170916 198694
rect 170862 198656 170864 198665
rect 170916 198656 170918 198665
rect 170862 198591 170918 198600
rect 170968 198490 170996 199407
rect 170864 198484 170916 198490
rect 170864 198426 170916 198432
rect 170956 198484 171008 198490
rect 170956 198426 171008 198432
rect 170876 194138 170904 198426
rect 170956 198280 171008 198286
rect 170956 198222 171008 198228
rect 170864 194132 170916 194138
rect 170864 194074 170916 194080
rect 170772 192908 170824 192914
rect 170772 192850 170824 192856
rect 170680 192024 170732 192030
rect 170680 191966 170732 191972
rect 170968 191894 170996 198222
rect 171060 198121 171088 199650
rect 171140 199640 171192 199646
rect 171140 199582 171192 199588
rect 171232 199640 171284 199646
rect 171232 199582 171284 199588
rect 171152 198354 171180 199582
rect 171244 198966 171272 199582
rect 171232 198960 171284 198966
rect 171232 198902 171284 198908
rect 171230 198384 171286 198393
rect 171140 198348 171192 198354
rect 171230 198319 171286 198328
rect 171140 198290 171192 198296
rect 171140 198212 171192 198218
rect 171140 198154 171192 198160
rect 171046 198112 171102 198121
rect 171046 198047 171102 198056
rect 171048 197872 171100 197878
rect 171048 197814 171100 197820
rect 171060 196246 171088 197814
rect 171152 197810 171180 198154
rect 171140 197804 171192 197810
rect 171140 197746 171192 197752
rect 171244 197062 171272 198319
rect 171336 197577 171364 199668
rect 171508 199504 171560 199510
rect 171508 199446 171560 199452
rect 171520 198200 171548 199446
rect 171428 198172 171548 198200
rect 171322 197568 171378 197577
rect 171322 197503 171378 197512
rect 171232 197056 171284 197062
rect 171232 196998 171284 197004
rect 171428 196704 171456 198172
rect 171508 198076 171560 198082
rect 171508 198018 171560 198024
rect 171152 196676 171456 196704
rect 171048 196240 171100 196246
rect 171048 196182 171100 196188
rect 170956 191888 171008 191894
rect 170956 191830 171008 191836
rect 171152 147529 171180 196676
rect 171322 196480 171378 196489
rect 171322 196415 171378 196424
rect 171336 192098 171364 196415
rect 171324 192092 171376 192098
rect 171324 192034 171376 192040
rect 171520 191978 171548 198018
rect 171612 197849 171640 199668
rect 171692 199640 171744 199646
rect 171692 199582 171744 199588
rect 171598 197840 171654 197849
rect 171598 197775 171654 197784
rect 171598 196072 171654 196081
rect 171598 196007 171654 196016
rect 171612 193050 171640 196007
rect 171600 193044 171652 193050
rect 171600 192986 171652 192992
rect 171244 191950 171548 191978
rect 171138 147520 171194 147529
rect 171244 147490 171272 191950
rect 171324 191820 171376 191826
rect 171324 191762 171376 191768
rect 171138 147455 171194 147464
rect 171232 147484 171284 147490
rect 171232 147426 171284 147432
rect 171336 147121 171364 191762
rect 171704 180794 171732 199582
rect 171796 197792 171824 199702
rect 172114 199736 172146 199744
rect 172196 199744 172252 199753
rect 172058 199679 172114 199688
rect 172302 199736 172382 199764
rect 172382 199718 172434 199724
rect 172196 199679 172252 199688
rect 171876 199640 171928 199646
rect 171876 199582 171928 199588
rect 172152 199640 172204 199646
rect 172152 199582 172204 199588
rect 172244 199640 172296 199646
rect 172486 199628 172514 200124
rect 172578 199764 172606 200124
rect 172670 199923 172698 200124
rect 172656 199914 172712 199923
rect 172656 199849 172712 199858
rect 172762 199764 172790 200124
rect 172854 199918 172882 200124
rect 172842 199912 172894 199918
rect 172946 199889 172974 200124
rect 172842 199854 172894 199860
rect 172932 199880 172988 199889
rect 173038 199850 173066 200124
rect 172932 199815 172988 199824
rect 173026 199844 173078 199850
rect 173026 199786 173078 199792
rect 172578 199753 172652 199764
rect 172578 199744 172666 199753
rect 172578 199736 172610 199744
rect 172610 199679 172666 199688
rect 172716 199736 172790 199764
rect 172486 199600 172560 199628
rect 172244 199582 172296 199588
rect 171888 198082 171916 199582
rect 172060 199572 172112 199578
rect 172060 199514 172112 199520
rect 172072 198966 172100 199514
rect 172060 198960 172112 198966
rect 172060 198902 172112 198908
rect 172060 198416 172112 198422
rect 172060 198358 172112 198364
rect 171876 198076 171928 198082
rect 171876 198018 171928 198024
rect 171796 197764 172008 197792
rect 171876 197668 171928 197674
rect 171876 197610 171928 197616
rect 171782 197432 171838 197441
rect 171782 197367 171838 197376
rect 171428 180766 171732 180794
rect 171322 147112 171378 147121
rect 171428 147082 171456 180766
rect 171508 155916 171560 155922
rect 171508 155858 171560 155864
rect 171322 147047 171378 147056
rect 171416 147076 171468 147082
rect 171416 147018 171468 147024
rect 170956 143336 171008 143342
rect 170956 143278 171008 143284
rect 170496 141772 170548 141778
rect 170496 141714 170548 141720
rect 170968 139890 170996 143278
rect 171520 139890 171548 155858
rect 171796 145761 171824 197367
rect 171888 190454 171916 197610
rect 171980 191962 172008 197764
rect 172072 196489 172100 198358
rect 172164 197985 172192 199582
rect 172256 198801 172284 199582
rect 172336 199572 172388 199578
rect 172336 199514 172388 199520
rect 172242 198792 172298 198801
rect 172242 198727 172298 198736
rect 172150 197976 172206 197985
rect 172150 197911 172206 197920
rect 172152 197804 172204 197810
rect 172152 197746 172204 197752
rect 172058 196480 172114 196489
rect 172058 196415 172114 196424
rect 172164 195974 172192 197746
rect 172072 195946 172192 195974
rect 172072 195702 172100 195946
rect 172060 195696 172112 195702
rect 172060 195638 172112 195644
rect 172348 193214 172376 199514
rect 172428 199504 172480 199510
rect 172428 199446 172480 199452
rect 172440 196704 172468 199446
rect 172532 198286 172560 199600
rect 172716 199594 172744 199736
rect 173130 199730 173158 200124
rect 173222 199889 173250 200124
rect 173208 199880 173264 199889
rect 173208 199815 173264 199824
rect 172946 199702 173158 199730
rect 173210 199776 173262 199782
rect 173210 199718 173262 199724
rect 172946 199628 172974 199702
rect 172624 199566 172744 199594
rect 172808 199600 172974 199628
rect 172624 198626 172652 199566
rect 172704 199504 172756 199510
rect 172704 199446 172756 199452
rect 172716 198966 172744 199446
rect 172704 198960 172756 198966
rect 172704 198902 172756 198908
rect 172612 198620 172664 198626
rect 172612 198562 172664 198568
rect 172612 198348 172664 198354
rect 172612 198290 172664 198296
rect 172520 198280 172572 198286
rect 172520 198222 172572 198228
rect 172624 197985 172652 198290
rect 172610 197976 172666 197985
rect 172610 197911 172666 197920
rect 172808 197441 172836 199600
rect 173222 199560 173250 199718
rect 173084 199532 173250 199560
rect 172980 199504 173032 199510
rect 172980 199446 173032 199452
rect 172992 198558 173020 199446
rect 173084 198937 173112 199532
rect 173314 199322 173342 200124
rect 173406 199560 173434 200124
rect 173498 199628 173526 200124
rect 173590 199730 173618 200124
rect 173682 199889 173710 200124
rect 173774 199918 173802 200124
rect 173866 199918 173894 200124
rect 173958 199918 173986 200124
rect 173762 199912 173814 199918
rect 173668 199880 173724 199889
rect 173762 199854 173814 199860
rect 173854 199912 173906 199918
rect 173854 199854 173906 199860
rect 173946 199912 173998 199918
rect 173946 199854 173998 199860
rect 173668 199815 173724 199824
rect 173808 199776 173860 199782
rect 173728 199736 173808 199764
rect 173590 199702 173664 199730
rect 173498 199600 173572 199628
rect 173406 199532 173480 199560
rect 173452 199322 173480 199532
rect 173268 199294 173342 199322
rect 173406 199294 173480 199322
rect 173070 198928 173126 198937
rect 173070 198863 173126 198872
rect 172980 198552 173032 198558
rect 172980 198494 173032 198500
rect 173268 198393 173296 199294
rect 173406 199152 173434 199294
rect 173360 199124 173434 199152
rect 173254 198384 173310 198393
rect 173254 198319 173310 198328
rect 172794 197432 172850 197441
rect 172794 197367 172850 197376
rect 173360 196790 173388 199124
rect 172796 196784 172848 196790
rect 172796 196726 172848 196732
rect 173348 196784 173400 196790
rect 173348 196726 173400 196732
rect 172440 196676 172652 196704
rect 172518 196344 172574 196353
rect 172518 196279 172574 196288
rect 172256 193186 172376 193214
rect 171968 191956 172020 191962
rect 171968 191898 172020 191904
rect 172256 191826 172284 193186
rect 172244 191820 172296 191826
rect 172244 191762 172296 191768
rect 171888 190426 172376 190454
rect 171782 145752 171838 145761
rect 171782 145687 171838 145696
rect 172348 144770 172376 190426
rect 172532 146033 172560 196279
rect 172624 147558 172652 196676
rect 172702 196344 172758 196353
rect 172702 196279 172758 196288
rect 172716 149734 172744 196279
rect 172808 150006 172836 196726
rect 173544 196722 173572 199600
rect 173636 198354 173664 199702
rect 173624 198348 173676 198354
rect 173624 198290 173676 198296
rect 172888 196716 172940 196722
rect 172888 196658 172940 196664
rect 173532 196716 173584 196722
rect 173532 196658 173584 196664
rect 172900 190262 172928 196658
rect 173162 196208 173218 196217
rect 173162 196143 173218 196152
rect 173176 192846 173204 196143
rect 173728 195650 173756 199736
rect 173808 199718 173860 199724
rect 173900 199776 173952 199782
rect 174050 199764 174078 200124
rect 174142 199918 174170 200124
rect 174130 199912 174182 199918
rect 174130 199854 174182 199860
rect 174234 199764 174262 200124
rect 173900 199718 173952 199724
rect 174004 199736 174078 199764
rect 174188 199736 174262 199764
rect 174326 199764 174354 200124
rect 174418 199923 174446 200124
rect 174404 199914 174460 199923
rect 174510 199918 174538 200124
rect 174602 199923 174630 200124
rect 174404 199849 174460 199858
rect 174498 199912 174550 199918
rect 174498 199854 174550 199860
rect 174588 199914 174644 199923
rect 174588 199849 174644 199858
rect 174694 199850 174722 200124
rect 174786 199918 174814 200124
rect 174878 199918 174906 200124
rect 174970 199918 174998 200124
rect 174774 199912 174826 199918
rect 174774 199854 174826 199860
rect 174866 199912 174918 199918
rect 174866 199854 174918 199860
rect 174958 199912 175010 199918
rect 174958 199854 175010 199860
rect 174682 199844 174734 199850
rect 174682 199786 174734 199792
rect 174452 199776 174504 199782
rect 174326 199736 174400 199764
rect 173808 199572 173860 199578
rect 173808 199514 173860 199520
rect 173820 198422 173848 199514
rect 173808 198416 173860 198422
rect 173808 198358 173860 198364
rect 173808 197736 173860 197742
rect 173808 197678 173860 197684
rect 173820 195770 173848 197678
rect 173912 197554 173940 199718
rect 174004 199578 174032 199736
rect 174188 199594 174216 199736
rect 173992 199572 174044 199578
rect 173992 199514 174044 199520
rect 174096 199566 174216 199594
rect 174268 199640 174320 199646
rect 174268 199582 174320 199588
rect 173912 197526 174032 197554
rect 173900 197464 173952 197470
rect 173900 197406 173952 197412
rect 173808 195764 173860 195770
rect 173808 195706 173860 195712
rect 173532 195628 173584 195634
rect 173728 195622 173848 195650
rect 173532 195570 173584 195576
rect 173438 194440 173494 194449
rect 173438 194375 173494 194384
rect 173452 194002 173480 194375
rect 173440 193996 173492 194002
rect 173440 193938 173492 193944
rect 173164 192840 173216 192846
rect 173164 192782 173216 192788
rect 172888 190256 172940 190262
rect 172888 190198 172940 190204
rect 173544 180794 173572 195570
rect 173716 195560 173768 195566
rect 173716 195502 173768 195508
rect 173728 194886 173756 195502
rect 173716 194880 173768 194886
rect 173716 194822 173768 194828
rect 173820 194206 173848 195622
rect 173808 194200 173860 194206
rect 173808 194142 173860 194148
rect 173622 194032 173678 194041
rect 173622 193967 173678 193976
rect 173636 193934 173664 193967
rect 173624 193928 173676 193934
rect 173624 193870 173676 193876
rect 173360 180766 173572 180794
rect 172888 158364 172940 158370
rect 172888 158306 172940 158312
rect 172796 150000 172848 150006
rect 172796 149942 172848 149948
rect 172704 149728 172756 149734
rect 172704 149670 172756 149676
rect 172612 147552 172664 147558
rect 172612 147494 172664 147500
rect 172518 146024 172574 146033
rect 172518 145959 172574 145968
rect 172336 144764 172388 144770
rect 172336 144706 172388 144712
rect 172428 144696 172480 144702
rect 172428 144638 172480 144644
rect 172440 139890 172468 144638
rect 172900 143546 172928 158306
rect 173360 151814 173388 180766
rect 173360 151786 173480 151814
rect 172888 143540 172940 143546
rect 172888 143482 172940 143488
rect 173164 143200 173216 143206
rect 173164 143142 173216 143148
rect 170324 139862 170476 139890
rect 170968 139862 171028 139890
rect 171520 139862 171580 139890
rect 172132 139862 172468 139890
rect 173176 139890 173204 143142
rect 173176 139862 173236 139890
rect 172684 139738 173020 139754
rect 172684 139732 173032 139738
rect 172684 139726 172980 139732
rect 172980 139674 173032 139680
rect 173452 139369 173480 151786
rect 173912 145897 173940 197406
rect 174004 196704 174032 197526
rect 174096 197470 174124 199566
rect 174280 199510 174308 199582
rect 174176 199504 174228 199510
rect 174176 199446 174228 199452
rect 174268 199504 174320 199510
rect 174268 199446 174320 199452
rect 174188 199073 174216 199446
rect 174266 199336 174322 199345
rect 174266 199271 174322 199280
rect 174174 199064 174230 199073
rect 174174 198999 174230 199008
rect 174280 198966 174308 199271
rect 174268 198960 174320 198966
rect 174174 198928 174230 198937
rect 174268 198902 174320 198908
rect 174174 198863 174230 198872
rect 174188 197946 174216 198863
rect 174176 197940 174228 197946
rect 174176 197882 174228 197888
rect 174084 197464 174136 197470
rect 174084 197406 174136 197412
rect 174004 196676 174216 196704
rect 173992 195152 174044 195158
rect 173992 195094 174044 195100
rect 174004 149802 174032 195094
rect 174084 194608 174136 194614
rect 174084 194550 174136 194556
rect 174096 149870 174124 194550
rect 174188 150385 174216 196676
rect 174372 194070 174400 199736
rect 175062 199764 175090 200124
rect 174452 199718 174504 199724
rect 174542 199744 174598 199753
rect 174360 194064 174412 194070
rect 174360 194006 174412 194012
rect 174268 193724 174320 193730
rect 174268 193666 174320 193672
rect 174280 190126 174308 193666
rect 174464 193214 174492 199718
rect 175016 199736 175090 199764
rect 174542 199679 174544 199688
rect 174596 199679 174598 199688
rect 174912 199708 174964 199714
rect 174544 199650 174596 199656
rect 174912 199650 174964 199656
rect 174544 199572 174596 199578
rect 174544 199514 174596 199520
rect 174556 194313 174584 199514
rect 174728 199504 174780 199510
rect 174728 199446 174780 199452
rect 174820 199504 174872 199510
rect 174820 199446 174872 199452
rect 174634 199336 174690 199345
rect 174634 199271 174690 199280
rect 174648 194449 174676 199271
rect 174740 195158 174768 199446
rect 174728 195152 174780 195158
rect 174728 195094 174780 195100
rect 174634 194440 174690 194449
rect 174634 194375 174690 194384
rect 174542 194304 174598 194313
rect 174542 194239 174598 194248
rect 174832 193730 174860 199446
rect 174924 198218 174952 199650
rect 174912 198212 174964 198218
rect 174912 198154 174964 198160
rect 175016 194614 175044 199736
rect 175154 199594 175182 200124
rect 175246 199923 175274 200124
rect 175232 199914 175288 199923
rect 175338 199918 175366 200124
rect 175232 199849 175288 199858
rect 175326 199912 175378 199918
rect 175326 199854 175378 199860
rect 175430 199850 175458 200124
rect 175522 199918 175550 200124
rect 175510 199912 175562 199918
rect 175510 199854 175562 199860
rect 175418 199844 175470 199850
rect 175418 199786 175470 199792
rect 175614 199764 175642 200124
rect 175568 199736 175642 199764
rect 175568 199730 175596 199736
rect 175522 199702 175596 199730
rect 175108 199566 175182 199594
rect 175372 199640 175424 199646
rect 175522 199628 175550 199702
rect 175706 199628 175734 200124
rect 175798 199730 175826 200124
rect 175890 199923 175918 200124
rect 175876 199914 175932 199923
rect 175982 199918 176010 200124
rect 176074 199918 176102 200124
rect 175876 199849 175932 199858
rect 175970 199912 176022 199918
rect 175970 199854 176022 199860
rect 176062 199912 176114 199918
rect 176062 199854 176114 199860
rect 176016 199776 176068 199782
rect 175798 199702 175964 199730
rect 176016 199718 176068 199724
rect 175936 199646 175964 199702
rect 175924 199640 175976 199646
rect 175522 199600 175596 199628
rect 175706 199600 175872 199628
rect 175372 199582 175424 199588
rect 175004 194608 175056 194614
rect 175004 194550 175056 194556
rect 174820 193724 174872 193730
rect 174820 193666 174872 193672
rect 174372 193186 174492 193214
rect 174268 190120 174320 190126
rect 174268 190062 174320 190068
rect 174268 155168 174320 155174
rect 174268 155110 174320 155116
rect 174174 150376 174230 150385
rect 174174 150311 174230 150320
rect 174084 149864 174136 149870
rect 174084 149806 174136 149812
rect 173992 149796 174044 149802
rect 173992 149738 174044 149744
rect 174280 147674 174308 155110
rect 174372 150113 174400 193186
rect 175108 193118 175136 199566
rect 175188 199504 175240 199510
rect 175188 199446 175240 199452
rect 175200 197713 175228 199446
rect 175384 198529 175412 199582
rect 175370 198520 175426 198529
rect 175370 198455 175426 198464
rect 175186 197704 175242 197713
rect 175186 197639 175242 197648
rect 175188 197532 175240 197538
rect 175188 197474 175240 197480
rect 175200 195838 175228 197474
rect 175372 197464 175424 197470
rect 175372 197406 175424 197412
rect 175462 197432 175518 197441
rect 175188 195832 175240 195838
rect 175188 195774 175240 195780
rect 174452 193112 174504 193118
rect 174452 193054 174504 193060
rect 175096 193112 175148 193118
rect 175096 193054 175148 193060
rect 174464 189718 174492 193054
rect 174542 192128 174598 192137
rect 174542 192063 174598 192072
rect 174452 189712 174504 189718
rect 174452 189654 174504 189660
rect 174358 150104 174414 150113
rect 174358 150039 174414 150048
rect 174280 147646 174492 147674
rect 173898 145888 173954 145897
rect 173898 145823 173954 145832
rect 173532 143540 173584 143546
rect 173532 143482 173584 143488
rect 174268 143540 174320 143546
rect 174268 143482 174320 143488
rect 173544 139890 173572 143482
rect 174280 139890 174308 143482
rect 174464 139890 174492 147646
rect 174556 141545 174584 192063
rect 175384 149938 175412 197406
rect 175462 197367 175518 197376
rect 175372 149932 175424 149938
rect 175372 149874 175424 149880
rect 175476 149705 175504 197367
rect 175568 196790 175596 199600
rect 175648 199504 175700 199510
rect 175648 199446 175700 199452
rect 175556 196784 175608 196790
rect 175556 196726 175608 196732
rect 175660 196602 175688 199446
rect 175568 196574 175688 196602
rect 175568 190330 175596 196574
rect 175844 196518 175872 199600
rect 175924 199582 175976 199588
rect 175924 199504 175976 199510
rect 175924 199446 175976 199452
rect 175936 199209 175964 199446
rect 175922 199200 175978 199209
rect 175922 199135 175978 199144
rect 176028 198801 176056 199718
rect 176166 199696 176194 200124
rect 176120 199668 176194 199696
rect 176014 198792 176070 198801
rect 176014 198727 176070 198736
rect 176120 197470 176148 199668
rect 176258 199628 176286 200124
rect 176350 199764 176378 200124
rect 176442 199923 176470 200124
rect 176428 199914 176484 199923
rect 176428 199849 176484 199858
rect 176350 199736 176424 199764
rect 176212 199600 176286 199628
rect 176108 197464 176160 197470
rect 176108 197406 176160 197412
rect 176212 197384 176240 199600
rect 176396 197742 176424 199736
rect 176534 199628 176562 200124
rect 176626 199696 176654 200124
rect 176718 199764 176746 200124
rect 176810 199918 176838 200124
rect 176902 199918 176930 200124
rect 176798 199912 176850 199918
rect 176798 199854 176850 199860
rect 176890 199912 176942 199918
rect 176890 199854 176942 199860
rect 176844 199776 176896 199782
rect 176718 199736 176792 199764
rect 176626 199668 176700 199696
rect 176534 199600 176608 199628
rect 176384 197736 176436 197742
rect 176384 197678 176436 197684
rect 176212 197356 176332 197384
rect 175832 196512 175884 196518
rect 175832 196454 175884 196460
rect 176200 195900 176252 195906
rect 176200 195842 176252 195848
rect 175648 195084 175700 195090
rect 175648 195026 175700 195032
rect 175556 190324 175608 190330
rect 175556 190266 175608 190272
rect 175660 189825 175688 195026
rect 176108 194880 176160 194886
rect 176108 194822 176160 194828
rect 175922 193080 175978 193089
rect 175922 193015 175978 193024
rect 175936 192273 175964 193015
rect 175922 192264 175978 192273
rect 175922 192199 175978 192208
rect 175646 189816 175702 189825
rect 175646 189751 175702 189760
rect 175462 149696 175518 149705
rect 175462 149631 175518 149640
rect 176120 146266 176148 194822
rect 176212 194818 176240 195842
rect 176200 194812 176252 194818
rect 176200 194754 176252 194760
rect 176304 194274 176332 197356
rect 176580 196874 176608 199600
rect 176672 198082 176700 199668
rect 176764 199646 176792 199736
rect 176994 199764 177022 200124
rect 177086 199889 177114 200124
rect 177072 199880 177128 199889
rect 177072 199815 177128 199824
rect 177178 199764 177206 200124
rect 176844 199718 176896 199724
rect 176948 199736 177022 199764
rect 177132 199736 177206 199764
rect 176752 199640 176804 199646
rect 176752 199582 176804 199588
rect 176660 198076 176712 198082
rect 176660 198018 176712 198024
rect 176396 196846 176608 196874
rect 176396 195090 176424 196846
rect 176476 196784 176528 196790
rect 176856 196772 176884 199718
rect 176476 196726 176528 196732
rect 176580 196744 176884 196772
rect 176384 195084 176436 195090
rect 176384 195026 176436 195032
rect 176292 194268 176344 194274
rect 176292 194210 176344 194216
rect 176108 146260 176160 146266
rect 176108 146202 176160 146208
rect 176488 146169 176516 196726
rect 176580 195158 176608 196744
rect 176948 196704 176976 199736
rect 177132 197402 177160 199736
rect 177270 199696 177298 200124
rect 177362 199832 177390 200124
rect 177454 199900 177482 200124
rect 177546 199968 177574 200124
rect 177546 199940 177620 199968
rect 177454 199872 177528 199900
rect 177362 199804 177436 199832
rect 177224 199668 177298 199696
rect 177120 197396 177172 197402
rect 177120 197338 177172 197344
rect 177120 196784 177172 196790
rect 177120 196726 177172 196732
rect 176764 196676 176976 196704
rect 177028 196716 177080 196722
rect 176660 196580 176712 196586
rect 176660 196522 176712 196528
rect 176568 195152 176620 195158
rect 176568 195094 176620 195100
rect 176672 149841 176700 196522
rect 176764 150414 176792 196676
rect 177028 196658 177080 196664
rect 176936 196308 176988 196314
rect 176936 196250 176988 196256
rect 176844 196172 176896 196178
rect 176844 196114 176896 196120
rect 176856 152658 176884 196114
rect 176844 152652 176896 152658
rect 176844 152594 176896 152600
rect 176948 152522 176976 196250
rect 177040 155446 177068 196658
rect 177132 189961 177160 196726
rect 177224 196586 177252 199668
rect 177408 196790 177436 199804
rect 177396 196784 177448 196790
rect 177396 196726 177448 196732
rect 177212 196580 177264 196586
rect 177212 196522 177264 196528
rect 177304 196580 177356 196586
rect 177304 196522 177356 196528
rect 177212 195152 177264 195158
rect 177212 195094 177264 195100
rect 177224 190466 177252 195094
rect 177212 190460 177264 190466
rect 177212 190402 177264 190408
rect 177316 190398 177344 196522
rect 177500 196314 177528 199872
rect 177592 196722 177620 199940
rect 177672 199844 177724 199850
rect 177672 199786 177724 199792
rect 177684 199646 177712 199786
rect 177672 199640 177724 199646
rect 177672 199582 177724 199588
rect 177672 197736 177724 197742
rect 177672 197678 177724 197684
rect 177580 196716 177632 196722
rect 177580 196658 177632 196664
rect 177488 196308 177540 196314
rect 177488 196250 177540 196256
rect 177684 195129 177712 197678
rect 177776 196178 177804 200246
rect 177868 198694 177896 200534
rect 178040 200048 178092 200054
rect 178040 199990 178092 199996
rect 177948 199640 178000 199646
rect 177946 199608 177948 199617
rect 178000 199608 178002 199617
rect 177946 199543 178002 199552
rect 177856 198688 177908 198694
rect 177856 198630 177908 198636
rect 177764 196172 177816 196178
rect 177764 196114 177816 196120
rect 177670 195120 177726 195129
rect 177670 195055 177726 195064
rect 177580 194880 177632 194886
rect 177580 194822 177632 194828
rect 177304 190392 177356 190398
rect 177304 190334 177356 190340
rect 177118 189952 177174 189961
rect 177118 189887 177174 189896
rect 177028 155440 177080 155446
rect 177028 155382 177080 155388
rect 176936 152516 176988 152522
rect 176936 152458 176988 152464
rect 176752 150408 176804 150414
rect 176752 150350 176804 150356
rect 176658 149832 176714 149841
rect 176658 149767 176714 149776
rect 177592 148238 177620 194822
rect 178052 192982 178080 199990
rect 178222 199880 178278 199889
rect 178222 199815 178278 199824
rect 178236 196586 178264 199815
rect 178224 196580 178276 196586
rect 178224 196522 178276 196528
rect 178040 192976 178092 192982
rect 178040 192918 178092 192924
rect 177580 148232 177632 148238
rect 177580 148174 177632 148180
rect 178408 146192 178460 146198
rect 176474 146160 176530 146169
rect 178408 146134 178460 146140
rect 176474 146095 176530 146104
rect 177212 146124 177264 146130
rect 177212 146066 177264 146072
rect 177120 144832 177172 144838
rect 177120 144774 177172 144780
rect 176292 143472 176344 143478
rect 176292 143414 176344 143420
rect 175740 143404 175792 143410
rect 175740 143346 175792 143352
rect 174542 141536 174598 141545
rect 174542 141471 174598 141480
rect 175752 139890 175780 143346
rect 176304 139890 176332 143414
rect 176476 141840 176528 141846
rect 176476 141782 176528 141788
rect 173544 139862 173788 139890
rect 174280 139862 174340 139890
rect 174464 139862 174892 139890
rect 175444 139862 175780 139890
rect 175996 139862 176332 139890
rect 176488 139890 176516 141782
rect 177132 140162 177160 144774
rect 177086 140134 177160 140162
rect 176488 139862 176548 139890
rect 177086 139876 177114 140134
rect 177224 139890 177252 146066
rect 178316 145512 178368 145518
rect 178316 145454 178368 145460
rect 178224 145444 178276 145450
rect 178224 145386 178276 145392
rect 178236 140162 178264 145386
rect 178328 143410 178356 145454
rect 178316 143404 178368 143410
rect 178316 143346 178368 143352
rect 178420 142154 178448 146134
rect 178190 140134 178264 140162
rect 178328 142126 178448 142154
rect 177224 139862 177652 139890
rect 178190 139876 178218 140134
rect 178328 139890 178356 142126
rect 178696 140350 178724 200602
rect 178776 200592 178828 200598
rect 178776 200534 178828 200540
rect 178788 140418 178816 200534
rect 178880 199918 178908 200670
rect 178868 199912 178920 199918
rect 178868 199854 178920 199860
rect 179050 199744 179106 199753
rect 179050 199679 179106 199688
rect 179064 199073 179092 199679
rect 179050 199064 179106 199073
rect 179050 198999 179106 199008
rect 178868 198960 178920 198966
rect 178868 198902 178920 198908
rect 178880 143410 178908 198902
rect 179420 197328 179472 197334
rect 179420 197270 179472 197276
rect 178960 196240 179012 196246
rect 178960 196182 179012 196188
rect 178972 152726 179000 196182
rect 179432 193118 179460 197270
rect 179984 195566 180012 200670
rect 180154 200560 180210 200569
rect 180154 200495 180210 200504
rect 180168 199850 180196 200495
rect 180156 199844 180208 199850
rect 180156 199786 180208 199792
rect 180156 199504 180208 199510
rect 180156 199446 180208 199452
rect 180064 198756 180116 198762
rect 180064 198698 180116 198704
rect 179972 195560 180024 195566
rect 179972 195502 180024 195508
rect 179420 193112 179472 193118
rect 179420 193054 179472 193060
rect 178960 152720 179012 152726
rect 178960 152662 179012 152668
rect 179604 147416 179656 147422
rect 179604 147358 179656 147364
rect 178960 147280 179012 147286
rect 178960 147222 179012 147228
rect 178868 143404 178920 143410
rect 178868 143346 178920 143352
rect 178776 140412 178828 140418
rect 178776 140354 178828 140360
rect 178684 140344 178736 140350
rect 178684 140286 178736 140292
rect 178972 139890 179000 147222
rect 179512 147212 179564 147218
rect 179512 147154 179564 147160
rect 179418 146840 179474 146849
rect 179418 146775 179474 146784
rect 179432 143274 179460 146775
rect 179524 143342 179552 147154
rect 179616 143478 179644 147358
rect 179696 147348 179748 147354
rect 179696 147290 179748 147296
rect 179708 143546 179736 147290
rect 179788 145376 179840 145382
rect 179788 145318 179840 145324
rect 179696 143540 179748 143546
rect 179696 143482 179748 143488
rect 179604 143472 179656 143478
rect 179604 143414 179656 143420
rect 179512 143336 179564 143342
rect 179512 143278 179564 143284
rect 179420 143268 179472 143274
rect 179420 143210 179472 143216
rect 179800 142154 179828 145318
rect 179432 142126 179828 142154
rect 179432 139890 179460 142126
rect 180076 140486 180104 198698
rect 180168 141710 180196 199446
rect 180260 147150 180288 200670
rect 180338 200424 180394 200433
rect 180338 200359 180394 200368
rect 180352 199782 180380 200359
rect 187700 200320 187752 200326
rect 187700 200262 187752 200268
rect 186688 200252 186740 200258
rect 186688 200194 186740 200200
rect 181996 199980 182048 199986
rect 181996 199922 182048 199928
rect 180340 199776 180392 199782
rect 180340 199718 180392 199724
rect 181076 199436 181128 199442
rect 181076 199378 181128 199384
rect 180432 197260 180484 197266
rect 180432 197202 180484 197208
rect 180340 194812 180392 194818
rect 180340 194754 180392 194760
rect 180248 147144 180300 147150
rect 180248 147086 180300 147092
rect 180352 144809 180380 194754
rect 180444 148170 180472 197202
rect 180892 149184 180944 149190
rect 180892 149126 180944 149132
rect 180432 148164 180484 148170
rect 180432 148106 180484 148112
rect 180432 147484 180484 147490
rect 180432 147426 180484 147432
rect 180444 147082 180472 147426
rect 180432 147076 180484 147082
rect 180432 147018 180484 147024
rect 180338 144800 180394 144809
rect 180338 144735 180394 144744
rect 180340 141908 180392 141914
rect 180340 141850 180392 141856
rect 180156 141704 180208 141710
rect 180156 141646 180208 141652
rect 180064 140480 180116 140486
rect 180064 140422 180116 140428
rect 178328 139862 178756 139890
rect 178972 139862 179308 139890
rect 179432 139862 179860 139890
rect 180064 139528 180116 139534
rect 180352 139482 180380 141850
rect 180904 139890 180932 149126
rect 181088 139890 181116 199378
rect 181168 198076 181220 198082
rect 181168 198018 181220 198024
rect 181444 198076 181496 198082
rect 181444 198018 181496 198024
rect 181180 196790 181208 198018
rect 181456 197878 181484 198018
rect 181444 197872 181496 197878
rect 181444 197814 181496 197820
rect 181168 196784 181220 196790
rect 181168 196726 181220 196732
rect 182008 196722 182036 199922
rect 182916 199504 182968 199510
rect 182916 199446 182968 199452
rect 182824 198824 182876 198830
rect 182824 198766 182876 198772
rect 182456 197396 182508 197402
rect 182456 197338 182508 197344
rect 181996 196716 182048 196722
rect 181996 196658 182048 196664
rect 182272 196512 182324 196518
rect 182272 196454 182324 196460
rect 181444 194404 181496 194410
rect 181444 194346 181496 194352
rect 181456 143138 181484 194346
rect 181536 194336 181588 194342
rect 181536 194278 181588 194284
rect 181548 143478 181576 194278
rect 182284 193905 182312 196454
rect 182468 195634 182496 197338
rect 182456 195628 182508 195634
rect 182456 195570 182508 195576
rect 182270 193896 182326 193905
rect 182270 193831 182326 193840
rect 182088 150068 182140 150074
rect 182088 150010 182140 150016
rect 182100 149190 182128 150010
rect 182088 149184 182140 149190
rect 182088 149126 182140 149132
rect 182272 144968 182324 144974
rect 182272 144910 182324 144916
rect 181536 143472 181588 143478
rect 181536 143414 181588 143420
rect 181720 143336 181772 143342
rect 181720 143278 181772 143284
rect 181352 143132 181404 143138
rect 181352 143074 181404 143080
rect 181444 143132 181496 143138
rect 181444 143074 181496 143080
rect 181364 142730 181392 143074
rect 181352 142724 181404 142730
rect 181352 142666 181404 142672
rect 181732 140894 181760 143278
rect 181720 140888 181772 140894
rect 181720 140830 181772 140836
rect 181732 139890 181760 140830
rect 182284 139890 182312 144910
rect 182836 140593 182864 198766
rect 182928 140826 182956 199446
rect 186596 198960 186648 198966
rect 186596 198902 186648 198908
rect 184296 198756 184348 198762
rect 184296 198698 184348 198704
rect 183008 196376 183060 196382
rect 183008 196318 183060 196324
rect 182916 140820 182968 140826
rect 182916 140762 182968 140768
rect 182822 140584 182878 140593
rect 182822 140519 182878 140528
rect 182928 139890 182956 140762
rect 183020 140321 183048 196318
rect 183100 195968 183152 195974
rect 183100 195910 183152 195916
rect 183006 140312 183062 140321
rect 183006 140247 183062 140256
rect 183112 140162 183140 195910
rect 183192 195220 183244 195226
rect 183192 195162 183244 195168
rect 183204 140457 183232 195162
rect 183834 194848 183890 194857
rect 183834 194783 183890 194792
rect 183848 194750 183876 194783
rect 183836 194744 183888 194750
rect 183836 194686 183888 194692
rect 184204 191548 184256 191554
rect 184204 191490 184256 191496
rect 183560 154556 183612 154562
rect 183560 154498 183612 154504
rect 183572 153270 183600 154498
rect 183560 153264 183612 153270
rect 183560 153206 183612 153212
rect 183468 145580 183520 145586
rect 183468 145522 183520 145528
rect 183480 144974 183508 145522
rect 183468 144968 183520 144974
rect 183468 144910 183520 144916
rect 183572 140758 183600 153206
rect 184216 151814 184244 191490
rect 184308 154562 184336 198698
rect 186504 194744 186556 194750
rect 186504 194686 186556 194692
rect 185676 192772 185728 192778
rect 185676 192714 185728 192720
rect 185584 189576 185636 189582
rect 185584 189518 185636 189524
rect 184296 154556 184348 154562
rect 184296 154498 184348 154504
rect 184664 153196 184716 153202
rect 184664 153138 184716 153144
rect 184572 152992 184624 152998
rect 184572 152934 184624 152940
rect 184388 152856 184440 152862
rect 184388 152798 184440 152804
rect 184296 152380 184348 152386
rect 184296 152322 184348 152328
rect 184124 151786 184244 151814
rect 184124 144906 184152 151786
rect 184308 146962 184336 152322
rect 184216 146934 184336 146962
rect 184112 144900 184164 144906
rect 184112 144842 184164 144848
rect 184020 142248 184072 142254
rect 184020 142190 184072 142196
rect 183560 140752 183612 140758
rect 183560 140694 183612 140700
rect 183190 140448 183246 140457
rect 183190 140383 183246 140392
rect 183112 140134 183324 140162
rect 180904 139862 180964 139890
rect 181088 139862 181516 139890
rect 181732 139862 182068 139890
rect 182284 139862 182620 139890
rect 182928 139862 183172 139890
rect 181272 139505 181300 139862
rect 183296 139534 183324 140134
rect 184032 139890 184060 142190
rect 184112 142044 184164 142050
rect 184112 141986 184164 141992
rect 183572 139862 184060 139890
rect 183572 139602 183600 139862
rect 183560 139596 183612 139602
rect 183560 139538 183612 139544
rect 183284 139528 183336 139534
rect 181258 139496 181314 139505
rect 180116 139476 180412 139482
rect 180064 139470 180412 139476
rect 180076 139454 180412 139470
rect 183284 139470 183336 139476
rect 181258 139431 181314 139440
rect 184124 139369 184152 141986
rect 184216 140690 184244 146934
rect 184296 143268 184348 143274
rect 184296 143210 184348 143216
rect 184308 142322 184336 143210
rect 184296 142316 184348 142322
rect 184296 142258 184348 142264
rect 184204 140684 184256 140690
rect 184204 140626 184256 140632
rect 184308 140162 184336 142258
rect 184400 142050 184428 152798
rect 184480 152788 184532 152794
rect 184480 152730 184532 152736
rect 184492 142050 184520 152730
rect 184388 142044 184440 142050
rect 184388 141986 184440 141992
rect 184480 142044 184532 142050
rect 184480 141986 184532 141992
rect 184584 140842 184612 152934
rect 184676 141302 184704 153138
rect 185492 152924 185544 152930
rect 185492 152866 185544 152872
rect 184756 146940 184808 146946
rect 184756 146882 184808 146888
rect 184768 141370 184796 146882
rect 185398 143168 185454 143177
rect 185398 143103 185454 143112
rect 185412 142497 185440 143103
rect 185398 142488 185454 142497
rect 185398 142423 185454 142432
rect 184848 142044 184900 142050
rect 184848 141986 184900 141992
rect 184756 141364 184808 141370
rect 184756 141306 184808 141312
rect 184664 141296 184716 141302
rect 184664 141238 184716 141244
rect 184262 140134 184336 140162
rect 184400 140814 184612 140842
rect 184262 139876 184290 140134
rect 184400 139369 184428 140814
rect 184480 140752 184532 140758
rect 184480 140694 184532 140700
rect 184492 139890 184520 140694
rect 184860 140622 184888 141986
rect 185308 141772 185360 141778
rect 185308 141714 185360 141720
rect 185320 141234 185348 141714
rect 185308 141228 185360 141234
rect 185308 141170 185360 141176
rect 184848 140616 184900 140622
rect 184848 140558 184900 140564
rect 185412 140162 185440 142423
rect 185366 140134 185440 140162
rect 184492 139862 184828 139890
rect 185366 139876 185394 140134
rect 185504 139369 185532 152866
rect 185596 140554 185624 189518
rect 185688 146810 185716 192714
rect 185860 191616 185912 191622
rect 185860 191558 185912 191564
rect 185768 191480 185820 191486
rect 185768 191422 185820 191428
rect 185676 146804 185728 146810
rect 185676 146746 185728 146752
rect 185676 144764 185728 144770
rect 185676 144706 185728 144712
rect 185688 144158 185716 144706
rect 185676 144152 185728 144158
rect 185676 144094 185728 144100
rect 185780 143546 185808 191422
rect 185872 150521 185900 191558
rect 185952 153128 186004 153134
rect 185952 153070 186004 153076
rect 185858 150512 185914 150521
rect 185858 150447 185914 150456
rect 185860 146940 185912 146946
rect 185860 146882 185912 146888
rect 185768 143540 185820 143546
rect 185768 143482 185820 143488
rect 185674 143440 185730 143449
rect 185674 143375 185730 143384
rect 185688 142633 185716 143375
rect 185674 142624 185730 142633
rect 185674 142559 185730 142568
rect 185584 140548 185636 140554
rect 185584 140490 185636 140496
rect 185688 139890 185716 142559
rect 185872 140706 185900 146882
rect 185964 141778 185992 153070
rect 186136 153060 186188 153066
rect 186136 153002 186188 153008
rect 186042 152416 186098 152425
rect 186042 152351 186098 152360
rect 186056 146946 186084 152351
rect 186044 146940 186096 146946
rect 186044 146882 186096 146888
rect 186044 146804 186096 146810
rect 186044 146746 186096 146752
rect 186056 142798 186084 146746
rect 186044 142792 186096 142798
rect 186044 142734 186096 142740
rect 186148 142050 186176 153002
rect 186228 152448 186280 152454
rect 186228 152390 186280 152396
rect 186136 142044 186188 142050
rect 186136 141986 186188 141992
rect 186240 141982 186268 152390
rect 186228 141976 186280 141982
rect 186228 141918 186280 141924
rect 185952 141772 186004 141778
rect 185952 141714 186004 141720
rect 185872 140678 186084 140706
rect 185688 139862 185932 139890
rect 123114 139360 123170 139369
rect 123114 139295 123170 139304
rect 123850 139360 123906 139369
rect 123850 139295 123906 139304
rect 129186 139360 129242 139369
rect 129186 139295 129242 139304
rect 131946 139360 132002 139369
rect 131946 139295 132002 139304
rect 166722 139360 166778 139369
rect 166722 139295 166778 139304
rect 173438 139360 173494 139369
rect 173438 139295 173494 139304
rect 184110 139360 184166 139369
rect 184110 139295 184166 139304
rect 184386 139360 184442 139369
rect 184386 139295 184442 139304
rect 185490 139360 185546 139369
rect 186056 139346 186084 140678
rect 186516 140185 186544 194686
rect 186502 140176 186558 140185
rect 186502 140111 186558 140120
rect 186226 139360 186282 139369
rect 186056 139318 186226 139346
rect 185490 139295 185546 139304
rect 186226 139295 186282 139304
rect 125600 80640 125652 80646
rect 130476 80640 130528 80646
rect 125600 80582 125652 80588
rect 130014 80608 130070 80617
rect 124126 78296 124182 78305
rect 124126 78231 124182 78240
rect 122472 67108 122524 67114
rect 122472 67050 122524 67056
rect 124140 65754 124168 78231
rect 125612 77178 125640 80582
rect 130476 80582 130528 80588
rect 131120 80640 131172 80646
rect 131304 80640 131356 80646
rect 131172 80588 131304 80594
rect 182134 80640 182186 80646
rect 131120 80582 131356 80588
rect 178038 80608 178094 80617
rect 130014 80543 130070 80552
rect 129738 80200 129794 80209
rect 129738 80135 129794 80144
rect 129004 80096 129056 80102
rect 129004 80038 129056 80044
rect 128542 79928 128598 79937
rect 128542 79863 128598 79872
rect 128556 78441 128584 79863
rect 129016 78577 129044 80038
rect 129002 78568 129058 78577
rect 129002 78503 129058 78512
rect 128542 78432 128598 78441
rect 128542 78367 128598 78376
rect 129752 77926 129780 80135
rect 129924 79416 129976 79422
rect 129924 79358 129976 79364
rect 129832 78056 129884 78062
rect 129832 77998 129884 78004
rect 129740 77920 129792 77926
rect 126978 77888 127034 77897
rect 129646 77888 129702 77897
rect 126978 77823 127034 77832
rect 128544 77852 128596 77858
rect 124864 77172 124916 77178
rect 124864 77114 124916 77120
rect 125600 77172 125652 77178
rect 125600 77114 125652 77120
rect 124128 65748 124180 65754
rect 124128 65690 124180 65696
rect 122288 3732 122340 3738
rect 122288 3674 122340 3680
rect 121460 3052 121512 3058
rect 121460 2994 121512 3000
rect 122300 480 122328 3674
rect 124876 3534 124904 77114
rect 126992 76430 127020 77823
rect 129740 77862 129792 77868
rect 129646 77823 129702 77832
rect 128544 77794 128596 77800
rect 126980 76424 127032 76430
rect 126980 76366 127032 76372
rect 126992 16574 127020 76366
rect 128556 74526 128584 77794
rect 129554 77616 129610 77625
rect 129554 77551 129610 77560
rect 129002 75168 129058 75177
rect 129002 75103 129058 75112
rect 128544 74520 128596 74526
rect 128544 74462 128596 74468
rect 128452 73636 128504 73642
rect 128452 73578 128504 73584
rect 128360 71052 128412 71058
rect 128360 70994 128412 71000
rect 126992 16546 127112 16574
rect 127084 3942 127112 16546
rect 127072 3936 127124 3942
rect 127072 3878 127124 3884
rect 125876 3596 125928 3602
rect 125876 3538 125928 3544
rect 123484 3528 123536 3534
rect 123484 3470 123536 3476
rect 124864 3528 124916 3534
rect 124864 3470 124916 3476
rect 123496 480 123524 3470
rect 124680 3120 124732 3126
rect 124680 3062 124732 3068
rect 124692 480 124720 3062
rect 125888 480 125916 3538
rect 128176 3528 128228 3534
rect 128176 3470 128228 3476
rect 126980 3324 127032 3330
rect 126980 3266 127032 3272
rect 126992 480 127020 3266
rect 128188 480 128216 3470
rect 128372 490 128400 70994
rect 128464 3330 128492 73578
rect 129016 3534 129044 75103
rect 129568 71058 129596 77551
rect 129660 73642 129688 77823
rect 129648 73636 129700 73642
rect 129648 73578 129700 73584
rect 129556 71052 129608 71058
rect 129556 70994 129608 71000
rect 129844 3806 129872 77998
rect 129936 77858 129964 79358
rect 129924 77852 129976 77858
rect 129924 77794 129976 77800
rect 129936 75177 129964 77794
rect 130028 77353 130056 80543
rect 130488 80442 130516 80582
rect 131132 80566 131344 80582
rect 182186 80588 182220 80594
rect 182134 80582 182220 80588
rect 178038 80543 178094 80552
rect 178132 80572 178184 80578
rect 130476 80436 130528 80442
rect 130476 80378 130528 80384
rect 130384 80368 130436 80374
rect 130384 80310 130436 80316
rect 130396 79694 130424 80310
rect 177764 80300 177816 80306
rect 177764 80242 177816 80248
rect 132052 80158 132388 80186
rect 177776 80170 177804 80242
rect 177764 80164 177816 80170
rect 130384 79688 130436 79694
rect 130384 79630 130436 79636
rect 130292 79620 130344 79626
rect 130292 79562 130344 79568
rect 130304 78810 130332 79562
rect 130568 79552 130620 79558
rect 130568 79494 130620 79500
rect 130292 78804 130344 78810
rect 130292 78746 130344 78752
rect 130014 77344 130070 77353
rect 130014 77279 130070 77288
rect 130474 75304 130530 75313
rect 130474 75239 130530 75248
rect 129922 75168 129978 75177
rect 129922 75103 129978 75112
rect 129924 73092 129976 73098
rect 129924 73034 129976 73040
rect 129832 3800 129884 3806
rect 129832 3742 129884 3748
rect 129936 3602 129964 73034
rect 130488 64874 130516 75239
rect 130580 75070 130608 79494
rect 131028 79484 131080 79490
rect 131028 79426 131080 79432
rect 130660 78056 130712 78062
rect 130660 77998 130712 78004
rect 130752 78056 130804 78062
rect 130752 77998 130804 78004
rect 130842 78024 130898 78033
rect 130672 77926 130700 77998
rect 130660 77920 130712 77926
rect 130660 77862 130712 77868
rect 130660 77716 130712 77722
rect 130660 77658 130712 77664
rect 130568 75064 130620 75070
rect 130568 75006 130620 75012
rect 130672 74730 130700 77658
rect 130660 74724 130712 74730
rect 130660 74666 130712 74672
rect 130764 73098 130792 77998
rect 130842 77959 130898 77968
rect 130856 77353 130884 77959
rect 130936 77784 130988 77790
rect 130936 77726 130988 77732
rect 130842 77344 130898 77353
rect 130842 77279 130898 77288
rect 130752 73092 130804 73098
rect 130752 73034 130804 73040
rect 130028 64846 130516 64874
rect 130028 16574 130056 64846
rect 130028 16546 130608 16574
rect 129924 3596 129976 3602
rect 129924 3538 129976 3544
rect 129004 3528 129056 3534
rect 129004 3470 129056 3476
rect 128452 3324 128504 3330
rect 128452 3266 128504 3272
rect 121062 354 121174 480
rect 120736 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 128372 462 128952 490
rect 130580 480 130608 16546
rect 130856 3738 130884 77279
rect 130948 75313 130976 77726
rect 131040 77722 131068 79426
rect 131212 77988 131264 77994
rect 131212 77930 131264 77936
rect 131028 77716 131080 77722
rect 131028 77658 131080 77664
rect 131028 75472 131080 75478
rect 131028 75414 131080 75420
rect 131120 75472 131172 75478
rect 131120 75414 131172 75420
rect 130934 75304 130990 75313
rect 130934 75239 130990 75248
rect 130936 75064 130988 75070
rect 130936 75006 130988 75012
rect 130844 3732 130896 3738
rect 130844 3674 130896 3680
rect 130948 3602 130976 75006
rect 131040 74866 131068 75414
rect 131132 75342 131160 75414
rect 131120 75336 131172 75342
rect 131120 75278 131172 75284
rect 131028 74860 131080 74866
rect 131028 74802 131080 74808
rect 131028 74724 131080 74730
rect 131028 74666 131080 74672
rect 131040 3806 131068 74666
rect 131028 3800 131080 3806
rect 131028 3742 131080 3748
rect 130936 3596 130988 3602
rect 130936 3538 130988 3544
rect 131132 3398 131160 75278
rect 131120 3392 131172 3398
rect 131120 3334 131172 3340
rect 131224 490 131252 77930
rect 132052 75857 132080 80158
rect 177764 80106 177816 80112
rect 178052 80102 178080 80543
rect 182146 80566 182220 80582
rect 178132 80514 178184 80520
rect 178040 80096 178092 80102
rect 132466 79914 132494 80036
rect 132558 79966 132586 80036
rect 132420 79886 132494 79914
rect 132546 79960 132598 79966
rect 132650 79937 132678 80036
rect 132742 79966 132770 80036
rect 132834 79966 132862 80036
rect 132926 79966 132954 80036
rect 133018 79966 133046 80036
rect 132730 79960 132782 79966
rect 132546 79902 132598 79908
rect 132636 79928 132692 79937
rect 132038 75848 132094 75857
rect 132038 75783 132094 75792
rect 131304 74996 131356 75002
rect 131304 74938 131356 74944
rect 131316 3874 131344 74938
rect 132420 73710 132448 79886
rect 132730 79902 132782 79908
rect 132822 79960 132874 79966
rect 132822 79902 132874 79908
rect 132914 79960 132966 79966
rect 132914 79902 132966 79908
rect 133006 79960 133058 79966
rect 133006 79902 133058 79908
rect 133110 79898 133138 80036
rect 133202 79971 133230 80036
rect 133188 79962 133244 79971
rect 132636 79863 132692 79872
rect 133098 79892 133150 79898
rect 133188 79897 133244 79906
rect 133098 79834 133150 79840
rect 132500 79824 132552 79830
rect 133294 79812 133322 80036
rect 133386 79966 133414 80036
rect 133478 79966 133506 80036
rect 133570 79971 133598 80036
rect 133374 79960 133426 79966
rect 133374 79902 133426 79908
rect 133466 79960 133518 79966
rect 133466 79902 133518 79908
rect 133556 79962 133612 79971
rect 133556 79897 133612 79906
rect 133662 79812 133690 80036
rect 133754 79898 133782 80036
rect 133846 79898 133874 80036
rect 133938 79898 133966 80036
rect 134030 79898 134058 80036
rect 133742 79892 133794 79898
rect 133742 79834 133794 79840
rect 133834 79892 133886 79898
rect 133834 79834 133886 79840
rect 133926 79892 133978 79898
rect 133926 79834 133978 79840
rect 134018 79892 134070 79898
rect 134018 79834 134070 79840
rect 133248 79801 133322 79812
rect 132500 79766 132552 79772
rect 132866 79792 132922 79801
rect 132512 78305 132540 79766
rect 132776 79756 132828 79762
rect 133234 79792 133322 79801
rect 132866 79727 132868 79736
rect 132776 79698 132828 79704
rect 132920 79727 132922 79736
rect 132960 79756 133012 79762
rect 132868 79698 132920 79704
rect 132960 79698 133012 79704
rect 133144 79756 133196 79762
rect 133290 79784 133322 79792
rect 133418 79792 133474 79801
rect 133234 79727 133290 79736
rect 133616 79784 133690 79812
rect 133616 79778 133644 79784
rect 133418 79727 133474 79736
rect 133570 79750 133644 79778
rect 134122 79778 134150 80036
rect 134214 79971 134242 80036
rect 134200 79962 134256 79971
rect 134200 79897 134256 79906
rect 134306 79812 134334 80036
rect 134398 79966 134426 80036
rect 134386 79960 134438 79966
rect 134386 79902 134438 79908
rect 134490 79898 134518 80036
rect 134582 79966 134610 80036
rect 134570 79960 134622 79966
rect 134570 79902 134622 79908
rect 134478 79892 134530 79898
rect 134478 79834 134530 79840
rect 134306 79784 134380 79812
rect 134352 79778 134380 79784
rect 134674 79778 134702 80036
rect 134766 79903 134794 80036
rect 134752 79894 134808 79903
rect 134752 79829 134808 79838
rect 133880 79756 133932 79762
rect 133144 79698 133196 79704
rect 132684 79620 132736 79626
rect 132684 79562 132736 79568
rect 132498 78296 132554 78305
rect 132498 78231 132554 78240
rect 132592 77376 132644 77382
rect 132592 77318 132644 77324
rect 132500 77308 132552 77314
rect 132500 77250 132552 77256
rect 132408 73704 132460 73710
rect 132408 73646 132460 73652
rect 132512 73098 132540 77250
rect 132604 75478 132632 77318
rect 132592 75472 132644 75478
rect 132592 75414 132644 75420
rect 132696 74534 132724 79562
rect 132788 77382 132816 79698
rect 132868 79484 132920 79490
rect 132868 79426 132920 79432
rect 132880 77654 132908 79426
rect 132868 77648 132920 77654
rect 132868 77590 132920 77596
rect 132776 77376 132828 77382
rect 132776 77318 132828 77324
rect 132776 76560 132828 76566
rect 132776 76502 132828 76508
rect 132788 76226 132816 76502
rect 132776 76220 132828 76226
rect 132776 76162 132828 76168
rect 132776 76084 132828 76090
rect 132776 76026 132828 76032
rect 132604 74506 132724 74534
rect 131396 73092 131448 73098
rect 131396 73034 131448 73040
rect 132500 73092 132552 73098
rect 132500 73034 132552 73040
rect 131408 72554 131436 73034
rect 131396 72548 131448 72554
rect 131396 72490 131448 72496
rect 131304 3868 131356 3874
rect 131304 3810 131356 3816
rect 131408 3670 131436 72490
rect 132604 72282 132632 74506
rect 132592 72276 132644 72282
rect 132592 72218 132644 72224
rect 132788 68474 132816 76026
rect 132776 68468 132828 68474
rect 132776 68410 132828 68416
rect 132684 67584 132736 67590
rect 132684 67526 132736 67532
rect 131488 65544 131540 65550
rect 131488 65486 131540 65492
rect 131396 3664 131448 3670
rect 131396 3606 131448 3612
rect 131500 3126 131528 65486
rect 132696 4826 132724 67526
rect 132880 37942 132908 77590
rect 132972 77294 133000 79698
rect 133050 79656 133106 79665
rect 133050 79591 133106 79600
rect 133064 77450 133092 79591
rect 133052 77444 133104 77450
rect 133052 77386 133104 77392
rect 132972 77266 133092 77294
rect 132960 76560 133012 76566
rect 132960 76502 133012 76508
rect 132972 60722 133000 76502
rect 133064 65958 133092 77266
rect 133156 72350 133184 79698
rect 133328 79688 133380 79694
rect 133234 79656 133290 79665
rect 133328 79630 133380 79636
rect 133234 79591 133290 79600
rect 133248 77466 133276 79591
rect 133340 77761 133368 79630
rect 133326 77752 133382 77761
rect 133326 77687 133382 77696
rect 133248 77438 133368 77466
rect 133236 77376 133288 77382
rect 133236 77318 133288 77324
rect 133144 72344 133196 72350
rect 133144 72286 133196 72292
rect 133248 67590 133276 77318
rect 133340 74534 133368 77438
rect 133432 77314 133460 79727
rect 133570 79676 133598 79750
rect 134122 79750 134196 79778
rect 134352 79750 134472 79778
rect 133880 79698 133932 79704
rect 133570 79648 133644 79676
rect 133420 77308 133472 77314
rect 133420 77250 133472 77256
rect 133616 76090 133644 79648
rect 133892 79608 133920 79698
rect 134064 79688 134116 79694
rect 134064 79630 134116 79636
rect 133800 79580 133920 79608
rect 133800 76566 133828 79580
rect 133972 79552 134024 79558
rect 133972 79494 134024 79500
rect 133880 79484 133932 79490
rect 133880 79426 133932 79432
rect 133892 77858 133920 79426
rect 133880 77852 133932 77858
rect 133880 77794 133932 77800
rect 133880 77648 133932 77654
rect 133880 77590 133932 77596
rect 133788 76560 133840 76566
rect 133788 76502 133840 76508
rect 133604 76084 133656 76090
rect 133604 76026 133656 76032
rect 133340 74506 133460 74534
rect 133432 71126 133460 74506
rect 133420 71120 133472 71126
rect 133420 71062 133472 71068
rect 133236 67584 133288 67590
rect 133236 67526 133288 67532
rect 133052 65952 133104 65958
rect 133052 65894 133104 65900
rect 132960 60716 133012 60722
rect 132960 60658 133012 60664
rect 132868 37936 132920 37942
rect 132868 37878 132920 37884
rect 133892 7614 133920 77590
rect 133984 76673 134012 79494
rect 134076 77353 134104 79630
rect 134168 78577 134196 79750
rect 134248 79688 134300 79694
rect 134248 79630 134300 79636
rect 134340 79688 134392 79694
rect 134340 79630 134392 79636
rect 134154 78568 134210 78577
rect 134154 78503 134210 78512
rect 134154 78432 134210 78441
rect 134154 78367 134210 78376
rect 134062 77344 134118 77353
rect 134062 77279 134118 77288
rect 133970 76664 134026 76673
rect 133970 76599 134026 76608
rect 134168 66162 134196 78367
rect 134260 68610 134288 79630
rect 134352 78305 134380 79630
rect 134444 78985 134472 79750
rect 134524 79756 134576 79762
rect 134524 79698 134576 79704
rect 134628 79750 134702 79778
rect 134430 78976 134486 78985
rect 134430 78911 134486 78920
rect 134338 78296 134394 78305
rect 134338 78231 134394 78240
rect 134444 78180 134472 78911
rect 134352 78152 134472 78180
rect 134352 77654 134380 78152
rect 134536 77976 134564 79698
rect 134444 77948 134564 77976
rect 134340 77648 134392 77654
rect 134340 77590 134392 77596
rect 134340 76424 134392 76430
rect 134340 76366 134392 76372
rect 134248 68604 134300 68610
rect 134248 68546 134300 68552
rect 134352 66230 134380 76366
rect 134444 70990 134472 77948
rect 134522 77888 134578 77897
rect 134522 77823 134524 77832
rect 134576 77823 134578 77832
rect 134524 77794 134576 77800
rect 134432 70984 134484 70990
rect 134432 70926 134484 70932
rect 134628 70394 134656 79750
rect 134858 79744 134886 80036
rect 134950 79971 134978 80036
rect 134936 79962 134992 79971
rect 135042 79966 135070 80036
rect 135134 79966 135162 80036
rect 134936 79897 134992 79906
rect 135030 79960 135082 79966
rect 135030 79902 135082 79908
rect 135122 79960 135174 79966
rect 135122 79902 135174 79908
rect 134812 79716 134886 79744
rect 135076 79756 135128 79762
rect 134708 79552 134760 79558
rect 134708 79494 134760 79500
rect 134720 77081 134748 79494
rect 134706 77072 134762 77081
rect 134706 77007 134762 77016
rect 134444 70366 134656 70394
rect 134340 66224 134392 66230
rect 134340 66166 134392 66172
rect 134156 66156 134208 66162
rect 134156 66098 134208 66104
rect 134064 66088 134116 66094
rect 134064 66030 134116 66036
rect 133972 49020 134024 49026
rect 133972 48962 134024 48968
rect 133880 7608 133932 7614
rect 133880 7550 133932 7556
rect 132684 4820 132736 4826
rect 132684 4762 132736 4768
rect 132960 3868 133012 3874
rect 132960 3810 133012 3816
rect 131488 3120 131540 3126
rect 131488 3062 131540 3068
rect 128924 354 128952 462
rect 129342 354 129454 480
rect 128924 326 129454 354
rect 129342 -960 129454 326
rect 130538 -960 130650 480
rect 131224 462 131344 490
rect 132972 480 133000 3810
rect 131316 354 131344 462
rect 131734 354 131846 480
rect 131316 326 131846 354
rect 131734 -960 131846 326
rect 132930 -960 133042 480
rect 133984 354 134012 48962
rect 134076 33794 134104 66030
rect 134168 35222 134196 66098
rect 134444 62014 134472 70366
rect 134812 66094 134840 79716
rect 135226 79744 135254 80036
rect 135318 79937 135346 80036
rect 135410 79966 135438 80036
rect 135398 79960 135450 79966
rect 135304 79928 135360 79937
rect 135398 79902 135450 79908
rect 135304 79863 135360 79872
rect 135502 79778 135530 80036
rect 135594 79966 135622 80036
rect 135686 79971 135714 80036
rect 135582 79960 135634 79966
rect 135582 79902 135634 79908
rect 135672 79962 135728 79971
rect 135778 79966 135806 80036
rect 135870 79966 135898 80036
rect 135962 79971 135990 80036
rect 135672 79897 135728 79906
rect 135766 79960 135818 79966
rect 135766 79902 135818 79908
rect 135858 79960 135910 79966
rect 135858 79902 135910 79908
rect 135948 79962 136004 79971
rect 136054 79966 136082 80036
rect 135948 79897 136004 79906
rect 136042 79960 136094 79966
rect 136042 79902 136094 79908
rect 135076 79698 135128 79704
rect 135180 79716 135254 79744
rect 135410 79750 135530 79778
rect 135720 79824 135772 79830
rect 136146 79812 136174 80036
rect 135720 79766 135772 79772
rect 135994 79792 136050 79801
rect 134982 79656 135038 79665
rect 134982 79591 135038 79600
rect 134996 71398 135024 79591
rect 135088 75682 135116 79698
rect 135180 76430 135208 79716
rect 135410 79676 135438 79750
rect 135410 79648 135484 79676
rect 135260 79620 135312 79626
rect 135260 79562 135312 79568
rect 135272 78198 135300 79562
rect 135352 79552 135404 79558
rect 135352 79494 135404 79500
rect 135260 78192 135312 78198
rect 135260 78134 135312 78140
rect 135364 77353 135392 79494
rect 135350 77344 135406 77353
rect 135350 77279 135406 77288
rect 135456 76430 135484 79648
rect 135628 79552 135680 79558
rect 135534 79520 135590 79529
rect 135628 79494 135680 79500
rect 135534 79455 135590 79464
rect 135168 76424 135220 76430
rect 135168 76366 135220 76372
rect 135444 76424 135496 76430
rect 135444 76366 135496 76372
rect 135076 75676 135128 75682
rect 135076 75618 135128 75624
rect 135352 75676 135404 75682
rect 135352 75618 135404 75624
rect 135364 74866 135392 75618
rect 135352 74860 135404 74866
rect 135352 74802 135404 74808
rect 134984 71392 135036 71398
rect 134984 71334 135036 71340
rect 135260 67516 135312 67522
rect 135260 67458 135312 67464
rect 134800 66088 134852 66094
rect 134800 66030 134852 66036
rect 134432 62008 134484 62014
rect 134432 61950 134484 61956
rect 134156 35216 134208 35222
rect 134156 35158 134208 35164
rect 134064 33788 134116 33794
rect 134064 33730 134116 33736
rect 135272 480 135300 67458
rect 135364 8974 135392 74802
rect 135548 66026 135576 79455
rect 135640 77382 135668 79494
rect 135628 77376 135680 77382
rect 135628 77318 135680 77324
rect 135628 76560 135680 76566
rect 135628 76502 135680 76508
rect 135640 68950 135668 76502
rect 135628 68944 135680 68950
rect 135628 68886 135680 68892
rect 135536 66020 135588 66026
rect 135536 65962 135588 65968
rect 135548 31074 135576 65962
rect 135732 60654 135760 79766
rect 135812 79756 135864 79762
rect 135994 79727 136050 79736
rect 136100 79784 136174 79812
rect 135812 79698 135864 79704
rect 135824 77625 135852 79698
rect 135904 79620 135956 79626
rect 135904 79562 135956 79568
rect 135810 77616 135866 77625
rect 135810 77551 135866 77560
rect 135812 77308 135864 77314
rect 135812 77250 135864 77256
rect 135720 60648 135772 60654
rect 135720 60590 135772 60596
rect 135824 59362 135852 77250
rect 135916 75682 135944 79562
rect 135904 75676 135956 75682
rect 135904 75618 135956 75624
rect 136008 70378 136036 79727
rect 136100 76566 136128 79784
rect 136238 79744 136266 80036
rect 136330 79830 136358 80036
rect 136422 79966 136450 80036
rect 136514 79971 136542 80036
rect 136410 79960 136462 79966
rect 136410 79902 136462 79908
rect 136500 79962 136556 79971
rect 136606 79966 136634 80036
rect 136500 79897 136556 79906
rect 136594 79960 136646 79966
rect 136594 79902 136646 79908
rect 136318 79824 136370 79830
rect 136698 79812 136726 80036
rect 136790 79966 136818 80036
rect 136778 79960 136830 79966
rect 136778 79902 136830 79908
rect 136318 79766 136370 79772
rect 136652 79784 136726 79812
rect 136192 79716 136266 79744
rect 136192 77314 136220 79716
rect 136548 79688 136600 79694
rect 136454 79656 136510 79665
rect 136548 79630 136600 79636
rect 136454 79591 136510 79600
rect 136364 79552 136416 79558
rect 136270 79520 136326 79529
rect 136364 79494 136416 79500
rect 136270 79455 136326 79464
rect 136284 78334 136312 79455
rect 136272 78328 136324 78334
rect 136272 78270 136324 78276
rect 136272 77376 136324 77382
rect 136272 77318 136324 77324
rect 136180 77308 136232 77314
rect 136180 77250 136232 77256
rect 136088 76560 136140 76566
rect 136088 76502 136140 76508
rect 136088 76424 136140 76430
rect 136088 76366 136140 76372
rect 135996 70372 136048 70378
rect 135996 70314 136048 70320
rect 136100 67318 136128 76366
rect 136284 70394 136312 77318
rect 136376 73846 136404 79494
rect 136364 73840 136416 73846
rect 136364 73782 136416 73788
rect 136468 72962 136496 79591
rect 136560 78266 136588 79630
rect 136548 78260 136600 78266
rect 136548 78202 136600 78208
rect 136652 76566 136680 79784
rect 136882 79744 136910 80036
rect 136974 79898 137002 80036
rect 137066 79937 137094 80036
rect 137158 79966 137186 80036
rect 137250 79966 137278 80036
rect 137342 79971 137370 80036
rect 137146 79960 137198 79966
rect 137052 79928 137108 79937
rect 136962 79892 137014 79898
rect 137146 79902 137198 79908
rect 137238 79960 137290 79966
rect 137238 79902 137290 79908
rect 137328 79962 137384 79971
rect 137434 79966 137462 80036
rect 137526 79966 137554 80036
rect 137328 79897 137384 79906
rect 137422 79960 137474 79966
rect 137422 79902 137474 79908
rect 137514 79960 137566 79966
rect 137514 79902 137566 79908
rect 137618 79898 137646 80036
rect 137052 79863 137108 79872
rect 137606 79892 137658 79898
rect 136962 79834 137014 79840
rect 137606 79834 137658 79840
rect 137376 79824 137428 79830
rect 137006 79792 137062 79801
rect 136882 79716 136956 79744
rect 137710 79801 137738 80036
rect 137376 79766 137428 79772
rect 137696 79792 137752 79801
rect 137006 79727 137062 79736
rect 137100 79756 137152 79762
rect 136732 79688 136784 79694
rect 136928 79665 136956 79716
rect 136732 79630 136784 79636
rect 136914 79656 136970 79665
rect 136744 78305 136772 79630
rect 136824 79620 136876 79626
rect 136914 79591 136970 79600
rect 136824 79562 136876 79568
rect 136730 78296 136786 78305
rect 136730 78231 136786 78240
rect 136732 78192 136784 78198
rect 136732 78134 136784 78140
rect 136640 76560 136692 76566
rect 136640 76502 136692 76508
rect 136456 72956 136508 72962
rect 136456 72898 136508 72904
rect 136192 70366 136312 70394
rect 136744 70394 136772 78134
rect 136836 76362 136864 79562
rect 136916 79552 136968 79558
rect 136916 79494 136968 79500
rect 136928 78470 136956 79494
rect 136916 78464 136968 78470
rect 136916 78406 136968 78412
rect 136824 76356 136876 76362
rect 136824 76298 136876 76304
rect 137020 75342 137048 79727
rect 137100 79698 137152 79704
rect 137008 75336 137060 75342
rect 137008 75278 137060 75284
rect 137008 74996 137060 75002
rect 137008 74938 137060 74944
rect 136744 70366 136956 70394
rect 136088 67312 136140 67318
rect 136088 67254 136140 67260
rect 136192 62082 136220 70366
rect 136928 65793 136956 70366
rect 136914 65784 136970 65793
rect 136914 65719 136970 65728
rect 136180 62076 136232 62082
rect 136180 62018 136232 62024
rect 135812 59356 135864 59362
rect 135812 59298 135864 59304
rect 136928 42090 136956 65719
rect 137020 59294 137048 74938
rect 137112 64802 137140 79698
rect 137192 79688 137244 79694
rect 137192 79630 137244 79636
rect 137282 79656 137338 79665
rect 137204 78402 137232 79630
rect 137282 79591 137338 79600
rect 137192 78396 137244 78402
rect 137192 78338 137244 78344
rect 137296 78198 137324 79591
rect 137284 78192 137336 78198
rect 137284 78134 137336 78140
rect 137388 77926 137416 79766
rect 137468 79756 137520 79762
rect 137696 79727 137752 79736
rect 137468 79698 137520 79704
rect 137376 77920 137428 77926
rect 137376 77862 137428 77868
rect 137480 77110 137508 79698
rect 137802 79676 137830 80036
rect 137894 79903 137922 80036
rect 137880 79894 137936 79903
rect 137986 79898 138014 80036
rect 138078 79966 138106 80036
rect 138170 79966 138198 80036
rect 138066 79960 138118 79966
rect 138066 79902 138118 79908
rect 138158 79960 138210 79966
rect 138158 79902 138210 79908
rect 137880 79829 137936 79838
rect 137974 79892 138026 79898
rect 137974 79834 138026 79840
rect 138262 79812 138290 80036
rect 138124 79784 138290 79812
rect 138354 79801 138382 80036
rect 138340 79792 138396 79801
rect 137928 79756 137980 79762
rect 137928 79698 137980 79704
rect 137756 79648 137830 79676
rect 137652 79620 137704 79626
rect 137652 79562 137704 79568
rect 137558 79520 137614 79529
rect 137558 79455 137614 79464
rect 137468 77104 137520 77110
rect 137468 77046 137520 77052
rect 137468 76560 137520 76566
rect 137468 76502 137520 76508
rect 137192 75336 137244 75342
rect 137192 75278 137244 75284
rect 137204 70242 137232 75278
rect 137192 70236 137244 70242
rect 137192 70178 137244 70184
rect 137480 64870 137508 76502
rect 137572 75614 137600 79455
rect 137664 76498 137692 79562
rect 137652 76492 137704 76498
rect 137652 76434 137704 76440
rect 137560 75608 137612 75614
rect 137560 75550 137612 75556
rect 137756 75002 137784 79648
rect 137940 78577 137968 79698
rect 138020 79688 138072 79694
rect 138020 79630 138072 79636
rect 137926 78568 137982 78577
rect 137926 78503 137982 78512
rect 138032 75914 138060 79630
rect 138124 79558 138152 79784
rect 138340 79727 138396 79736
rect 138446 79744 138474 80036
rect 138538 79937 138566 80036
rect 138630 79966 138658 80036
rect 138722 79966 138750 80036
rect 138814 79966 138842 80036
rect 138618 79960 138670 79966
rect 138524 79928 138580 79937
rect 138618 79902 138670 79908
rect 138710 79960 138762 79966
rect 138710 79902 138762 79908
rect 138802 79960 138854 79966
rect 138802 79902 138854 79908
rect 138524 79863 138580 79872
rect 138572 79824 138624 79830
rect 138570 79792 138572 79801
rect 138756 79824 138808 79830
rect 138624 79792 138626 79801
rect 138446 79716 138520 79744
rect 138756 79766 138808 79772
rect 138570 79727 138626 79736
rect 138296 79688 138348 79694
rect 138296 79630 138348 79636
rect 138204 79620 138256 79626
rect 138204 79562 138256 79568
rect 138112 79552 138164 79558
rect 138112 79494 138164 79500
rect 138216 78826 138244 79562
rect 137940 75886 138060 75914
rect 138124 78798 138244 78826
rect 137744 74996 137796 75002
rect 137744 74938 137796 74944
rect 137940 71602 137968 75886
rect 138124 75274 138152 78798
rect 138204 78736 138256 78742
rect 138204 78678 138256 78684
rect 138216 75914 138244 78678
rect 138308 77314 138336 79630
rect 138492 77704 138520 79716
rect 138572 79688 138624 79694
rect 138572 79630 138624 79636
rect 138664 79688 138716 79694
rect 138664 79630 138716 79636
rect 138584 78742 138612 79630
rect 138572 78736 138624 78742
rect 138572 78678 138624 78684
rect 138676 78674 138704 79630
rect 138664 78668 138716 78674
rect 138664 78610 138716 78616
rect 138768 77926 138796 79766
rect 138906 79676 138934 80036
rect 138998 79971 139026 80036
rect 138984 79962 139040 79971
rect 138984 79897 139040 79906
rect 139090 79898 139118 80036
rect 139182 79903 139210 80036
rect 139274 79966 139302 80036
rect 139366 79966 139394 80036
rect 139262 79960 139314 79966
rect 139078 79892 139130 79898
rect 139078 79834 139130 79840
rect 139168 79894 139224 79903
rect 139262 79902 139314 79908
rect 139354 79960 139406 79966
rect 139458 79937 139486 80036
rect 139550 79966 139578 80036
rect 139642 79966 139670 80036
rect 139734 79971 139762 80036
rect 139538 79960 139590 79966
rect 139354 79902 139406 79908
rect 139444 79928 139500 79937
rect 139538 79902 139590 79908
rect 139630 79960 139682 79966
rect 139630 79902 139682 79908
rect 139720 79962 139776 79971
rect 139826 79966 139854 80036
rect 139918 79966 139946 80036
rect 139720 79897 139776 79906
rect 139814 79960 139866 79966
rect 139814 79902 139866 79908
rect 139906 79960 139958 79966
rect 139906 79902 139958 79908
rect 139444 79863 139500 79872
rect 139168 79829 139224 79838
rect 140010 79812 140038 80036
rect 140102 79966 140130 80036
rect 140194 79966 140222 80036
rect 140286 79971 140314 80036
rect 140090 79960 140142 79966
rect 140090 79902 140142 79908
rect 140182 79960 140234 79966
rect 140182 79902 140234 79908
rect 140272 79962 140328 79971
rect 140378 79966 140406 80036
rect 140272 79897 140328 79906
rect 140366 79960 140418 79966
rect 140366 79902 140418 79908
rect 139964 79784 140038 79812
rect 139032 79756 139084 79762
rect 139032 79698 139084 79704
rect 139124 79756 139176 79762
rect 139124 79698 139176 79704
rect 139584 79756 139636 79762
rect 139584 79698 139636 79704
rect 139768 79756 139820 79762
rect 139768 79698 139820 79704
rect 138860 79648 138934 79676
rect 138756 77920 138808 77926
rect 138756 77862 138808 77868
rect 138492 77676 138612 77704
rect 138296 77308 138348 77314
rect 138296 77250 138348 77256
rect 138480 77308 138532 77314
rect 138480 77250 138532 77256
rect 138216 75886 138336 75914
rect 138204 75744 138256 75750
rect 138204 75686 138256 75692
rect 138020 75268 138072 75274
rect 138020 75210 138072 75216
rect 138112 75268 138164 75274
rect 138112 75210 138164 75216
rect 138032 75002 138060 75210
rect 138020 74996 138072 75002
rect 138020 74938 138072 74944
rect 138216 72486 138244 75686
rect 138204 72480 138256 72486
rect 138204 72422 138256 72428
rect 137928 71596 137980 71602
rect 137928 71538 137980 71544
rect 138020 68672 138072 68678
rect 138020 68614 138072 68620
rect 137468 64864 137520 64870
rect 137468 64806 137520 64812
rect 137100 64796 137152 64802
rect 137100 64738 137152 64744
rect 137008 59288 137060 59294
rect 137008 59230 137060 59236
rect 136916 42084 136968 42090
rect 136916 42026 136968 42032
rect 138032 39370 138060 68614
rect 138110 66056 138166 66065
rect 138110 65991 138166 66000
rect 138124 40730 138152 65991
rect 138112 40724 138164 40730
rect 138112 40666 138164 40672
rect 138112 40044 138164 40050
rect 138112 39986 138164 39992
rect 138020 39364 138072 39370
rect 138020 39306 138072 39312
rect 135536 31068 135588 31074
rect 135536 31010 135588 31016
rect 135352 8968 135404 8974
rect 135352 8910 135404 8916
rect 138124 6914 138152 39986
rect 138216 15910 138244 72422
rect 138308 67250 138336 75886
rect 138492 75698 138520 77250
rect 138400 75670 138520 75698
rect 138296 67244 138348 67250
rect 138296 67186 138348 67192
rect 138400 56574 138428 75670
rect 138480 75268 138532 75274
rect 138480 75210 138532 75216
rect 138492 66065 138520 75210
rect 138584 68678 138612 77676
rect 138572 68672 138624 68678
rect 138572 68614 138624 68620
rect 138860 67182 138888 79648
rect 138938 78024 138994 78033
rect 138938 77959 138994 77968
rect 138952 75818 138980 77959
rect 138940 75812 138992 75818
rect 138940 75754 138992 75760
rect 139044 70174 139072 79698
rect 139136 73778 139164 79698
rect 139214 79656 139270 79665
rect 139214 79591 139270 79600
rect 139228 75750 139256 79591
rect 139490 79384 139546 79393
rect 139490 79319 139546 79328
rect 139308 77920 139360 77926
rect 139308 77862 139360 77868
rect 139216 75744 139268 75750
rect 139216 75686 139268 75692
rect 139320 74934 139348 77862
rect 139504 77790 139532 79319
rect 139596 78577 139624 79698
rect 139674 79656 139730 79665
rect 139674 79591 139730 79600
rect 139688 79422 139716 79591
rect 139676 79416 139728 79422
rect 139676 79358 139728 79364
rect 139582 78568 139638 78577
rect 139582 78503 139638 78512
rect 139584 78396 139636 78402
rect 139584 78338 139636 78344
rect 139492 77784 139544 77790
rect 139492 77726 139544 77732
rect 139308 74928 139360 74934
rect 139308 74870 139360 74876
rect 139596 74526 139624 78338
rect 139780 75750 139808 79698
rect 139964 79608 139992 79784
rect 140470 79778 140498 80036
rect 140562 79966 140590 80036
rect 140550 79960 140602 79966
rect 140550 79902 140602 79908
rect 140654 79812 140682 80036
rect 140608 79784 140682 79812
rect 140136 79756 140188 79762
rect 140470 79750 140544 79778
rect 140136 79698 140188 79704
rect 140044 79688 140096 79694
rect 140044 79630 140096 79636
rect 139872 79580 139992 79608
rect 139768 75744 139820 75750
rect 139768 75686 139820 75692
rect 139584 74520 139636 74526
rect 139584 74462 139636 74468
rect 139124 73772 139176 73778
rect 139124 73714 139176 73720
rect 139596 70394 139624 74462
rect 139596 70366 139808 70394
rect 139032 70168 139084 70174
rect 139032 70110 139084 70116
rect 138848 67176 138900 67182
rect 138848 67118 138900 67124
rect 138478 66056 138534 66065
rect 138478 65991 138534 66000
rect 139582 65648 139638 65657
rect 139582 65583 139638 65592
rect 138388 56568 138440 56574
rect 138388 56510 138440 56516
rect 138664 55276 138716 55282
rect 138664 55218 138716 55224
rect 138204 15904 138256 15910
rect 138204 15846 138256 15852
rect 138124 6886 138612 6914
rect 137652 3664 137704 3670
rect 137652 3606 137704 3612
rect 136456 3188 136508 3194
rect 136456 3130 136508 3136
rect 136468 480 136496 3130
rect 137664 480 137692 3606
rect 138584 3482 138612 6886
rect 138676 3670 138704 55218
rect 139596 36582 139624 65583
rect 139584 36576 139636 36582
rect 139584 36518 139636 36524
rect 139780 6186 139808 70366
rect 139872 60586 139900 79580
rect 139952 78668 140004 78674
rect 139952 78610 140004 78616
rect 139964 70106 139992 78610
rect 140056 76702 140084 79630
rect 140148 78674 140176 79698
rect 140412 79688 140464 79694
rect 140226 79656 140282 79665
rect 140412 79630 140464 79636
rect 140226 79591 140282 79600
rect 140320 79620 140372 79626
rect 140240 79558 140268 79591
rect 140320 79562 140372 79568
rect 140228 79552 140280 79558
rect 140228 79494 140280 79500
rect 140228 79416 140280 79422
rect 140228 79358 140280 79364
rect 140136 78668 140188 78674
rect 140136 78610 140188 78616
rect 140136 78192 140188 78198
rect 140136 78134 140188 78140
rect 140044 76696 140096 76702
rect 140044 76638 140096 76644
rect 140044 75880 140096 75886
rect 140044 75822 140096 75828
rect 140056 71670 140084 75822
rect 140044 71664 140096 71670
rect 140044 71606 140096 71612
rect 139952 70100 140004 70106
rect 139952 70042 140004 70048
rect 140044 69080 140096 69086
rect 140044 69022 140096 69028
rect 139860 60580 139912 60586
rect 139860 60522 139912 60528
rect 139768 6180 139820 6186
rect 139768 6122 139820 6128
rect 140056 3874 140084 69022
rect 140148 65822 140176 78134
rect 140240 75886 140268 79358
rect 140228 75880 140280 75886
rect 140228 75822 140280 75828
rect 140228 75744 140280 75750
rect 140228 75686 140280 75692
rect 140136 65816 140188 65822
rect 140136 65758 140188 65764
rect 140240 65657 140268 75686
rect 140332 72894 140360 79562
rect 140424 78402 140452 79630
rect 140516 79422 140544 79750
rect 140504 79416 140556 79422
rect 140504 79358 140556 79364
rect 140504 78668 140556 78674
rect 140504 78610 140556 78616
rect 140412 78396 140464 78402
rect 140412 78338 140464 78344
rect 140516 77897 140544 78610
rect 140502 77888 140558 77897
rect 140502 77823 140558 77832
rect 140412 77648 140464 77654
rect 140412 77590 140464 77596
rect 140424 74186 140452 77590
rect 140608 74390 140636 79784
rect 140746 79744 140774 80036
rect 140838 79971 140866 80036
rect 140824 79962 140880 79971
rect 140824 79897 140880 79906
rect 140700 79716 140774 79744
rect 140930 79744 140958 80036
rect 141022 79898 141050 80036
rect 141010 79892 141062 79898
rect 141010 79834 141062 79840
rect 140930 79716 141004 79744
rect 140700 77654 140728 79716
rect 140780 79620 140832 79626
rect 140780 79562 140832 79568
rect 140872 79620 140924 79626
rect 140872 79562 140924 79568
rect 140792 78198 140820 79562
rect 140780 78192 140832 78198
rect 140780 78134 140832 78140
rect 140688 77648 140740 77654
rect 140688 77590 140740 77596
rect 140884 76226 140912 79562
rect 140976 76945 141004 79716
rect 141114 79676 141142 80036
rect 141206 79744 141234 80036
rect 141298 79898 141326 80036
rect 141390 79937 141418 80036
rect 141376 79928 141432 79937
rect 141286 79892 141338 79898
rect 141482 79898 141510 80036
rect 141376 79863 141432 79872
rect 141470 79892 141522 79898
rect 141286 79834 141338 79840
rect 141470 79834 141522 79840
rect 141574 79744 141602 80036
rect 141206 79716 141280 79744
rect 141114 79648 141188 79676
rect 141056 79552 141108 79558
rect 141056 79494 141108 79500
rect 140962 76936 141018 76945
rect 140962 76871 141018 76880
rect 140964 76696 141016 76702
rect 140964 76638 141016 76644
rect 140872 76220 140924 76226
rect 140872 76162 140924 76168
rect 140976 75138 141004 76638
rect 140964 75132 141016 75138
rect 140964 75074 141016 75080
rect 140596 74384 140648 74390
rect 140596 74326 140648 74332
rect 140412 74180 140464 74186
rect 140412 74122 140464 74128
rect 140320 72888 140372 72894
rect 140320 72830 140372 72836
rect 141068 69766 141096 79494
rect 141160 76634 141188 79648
rect 141252 79608 141280 79716
rect 141528 79716 141602 79744
rect 141332 79620 141384 79626
rect 141252 79580 141332 79608
rect 141332 79562 141384 79568
rect 141424 79620 141476 79626
rect 141424 79562 141476 79568
rect 141240 79484 141292 79490
rect 141240 79426 141292 79432
rect 141332 79484 141384 79490
rect 141332 79426 141384 79432
rect 141252 76702 141280 79426
rect 141240 76696 141292 76702
rect 141240 76638 141292 76644
rect 141148 76628 141200 76634
rect 141148 76570 141200 76576
rect 141240 75268 141292 75274
rect 141240 75210 141292 75216
rect 141148 75200 141200 75206
rect 141148 75142 141200 75148
rect 141056 69760 141108 69766
rect 141056 69702 141108 69708
rect 140226 65648 140282 65657
rect 140226 65583 140282 65592
rect 141160 65550 141188 75142
rect 141252 68338 141280 75210
rect 141344 69834 141372 79426
rect 141436 78305 141464 79562
rect 141422 78296 141478 78305
rect 141422 78231 141478 78240
rect 141422 77888 141478 77897
rect 141422 77823 141478 77832
rect 141332 69828 141384 69834
rect 141332 69770 141384 69776
rect 141436 68406 141464 77823
rect 141528 72418 141556 79716
rect 141666 79608 141694 80036
rect 141758 79898 141786 80036
rect 141746 79892 141798 79898
rect 141746 79834 141798 79840
rect 141850 79744 141878 80036
rect 141942 79812 141970 80036
rect 142034 79966 142062 80036
rect 142022 79960 142074 79966
rect 142022 79902 142074 79908
rect 142126 79812 142154 80036
rect 142218 79898 142246 80036
rect 142310 79903 142338 80036
rect 142206 79892 142258 79898
rect 142206 79834 142258 79840
rect 142296 79894 142352 79903
rect 142402 79898 142430 80036
rect 142494 79966 142522 80036
rect 142482 79960 142534 79966
rect 142482 79902 142534 79908
rect 142296 79829 142352 79838
rect 142390 79892 142442 79898
rect 142390 79834 142442 79840
rect 142586 79812 142614 80036
rect 142678 79937 142706 80036
rect 142664 79928 142720 79937
rect 142664 79863 142720 79872
rect 142770 79812 142798 80036
rect 142862 79966 142890 80036
rect 142850 79960 142902 79966
rect 142850 79902 142902 79908
rect 142954 79812 142982 80036
rect 141942 79784 142016 79812
rect 141620 79580 141694 79608
rect 141804 79716 141878 79744
rect 141620 75274 141648 79580
rect 141804 79472 141832 79716
rect 141988 79608 142016 79784
rect 141712 79444 141832 79472
rect 141896 79580 142016 79608
rect 142080 79784 142154 79812
rect 142540 79784 142614 79812
rect 142724 79784 142798 79812
rect 142908 79784 142982 79812
rect 141712 78169 141740 79444
rect 141698 78160 141754 78169
rect 141698 78095 141754 78104
rect 141896 77178 141924 79580
rect 141976 79484 142028 79490
rect 141976 79426 142028 79432
rect 141884 77172 141936 77178
rect 141884 77114 141936 77120
rect 141608 75268 141660 75274
rect 141608 75210 141660 75216
rect 141988 75206 142016 79426
rect 142080 78062 142108 79784
rect 142344 79756 142396 79762
rect 142344 79698 142396 79704
rect 142160 79688 142212 79694
rect 142160 79630 142212 79636
rect 142068 78056 142120 78062
rect 142068 77998 142120 78004
rect 142172 77976 142200 79630
rect 142252 79620 142304 79626
rect 142252 79562 142304 79568
rect 142264 79393 142292 79562
rect 142250 79384 142306 79393
rect 142250 79319 142306 79328
rect 142252 79144 142304 79150
rect 142252 79086 142304 79092
rect 142264 78198 142292 79086
rect 142252 78192 142304 78198
rect 142252 78134 142304 78140
rect 142172 77948 142292 77976
rect 142158 77888 142214 77897
rect 142264 77858 142292 77948
rect 142158 77823 142214 77832
rect 142252 77852 142304 77858
rect 141976 75200 142028 75206
rect 141976 75142 142028 75148
rect 142172 72826 142200 77823
rect 142252 77794 142304 77800
rect 142356 77489 142384 79698
rect 142540 77994 142568 79784
rect 142620 79620 142672 79626
rect 142620 79562 142672 79568
rect 142528 77988 142580 77994
rect 142528 77930 142580 77936
rect 142342 77480 142398 77489
rect 142342 77415 142398 77424
rect 142528 75676 142580 75682
rect 142528 75618 142580 75624
rect 142436 75132 142488 75138
rect 142436 75074 142488 75080
rect 142252 74520 142304 74526
rect 142252 74462 142304 74468
rect 142264 73982 142292 74462
rect 142252 73976 142304 73982
rect 142252 73918 142304 73924
rect 142160 72820 142212 72826
rect 142160 72762 142212 72768
rect 141516 72412 141568 72418
rect 141516 72354 141568 72360
rect 142172 69086 142200 72762
rect 142160 69080 142212 69086
rect 142160 69022 142212 69028
rect 142160 68876 142212 68882
rect 142160 68818 142212 68824
rect 141424 68400 141476 68406
rect 141424 68342 141476 68348
rect 141240 68332 141292 68338
rect 141240 68274 141292 68280
rect 141424 67652 141476 67658
rect 141424 67594 141476 67600
rect 141148 65544 141200 65550
rect 141148 65486 141200 65492
rect 141240 4140 141292 4146
rect 141240 4082 141292 4088
rect 140044 3868 140096 3874
rect 140044 3810 140096 3816
rect 138664 3664 138716 3670
rect 138664 3606 138716 3612
rect 140044 3528 140096 3534
rect 138584 3454 138888 3482
rect 140044 3470 140096 3476
rect 138860 480 138888 3454
rect 140056 480 140084 3470
rect 141252 480 141280 4082
rect 141436 3194 141464 67594
rect 141516 66292 141568 66298
rect 141516 66234 141568 66240
rect 141528 3534 141556 66234
rect 142172 60734 142200 68818
rect 142264 67658 142292 73918
rect 142344 73092 142396 73098
rect 142344 73034 142396 73040
rect 142356 72690 142384 73034
rect 142344 72684 142396 72690
rect 142344 72626 142396 72632
rect 142252 67652 142304 67658
rect 142252 67594 142304 67600
rect 142356 66298 142384 72626
rect 142448 69970 142476 75074
rect 142540 74254 142568 75618
rect 142528 74248 142580 74254
rect 142528 74190 142580 74196
rect 142436 69964 142488 69970
rect 142436 69906 142488 69912
rect 142344 66292 142396 66298
rect 142344 66234 142396 66240
rect 142344 66156 142396 66162
rect 142344 66098 142396 66104
rect 142172 60706 142292 60734
rect 142264 40050 142292 60706
rect 142356 55282 142384 66098
rect 142344 55276 142396 55282
rect 142344 55218 142396 55224
rect 142252 40044 142304 40050
rect 142252 39986 142304 39992
rect 142448 6914 142476 69906
rect 142540 65498 142568 74190
rect 142632 67522 142660 79562
rect 142724 79234 142752 79784
rect 142908 79744 142936 79784
rect 143046 79744 143074 80036
rect 142816 79716 142936 79744
rect 143000 79716 143074 79744
rect 143138 79744 143166 80036
rect 143230 79903 143258 80036
rect 143322 79966 143350 80036
rect 143310 79960 143362 79966
rect 143216 79894 143272 79903
rect 143310 79902 143362 79908
rect 143216 79829 143272 79838
rect 143414 79778 143442 80036
rect 143368 79750 143442 79778
rect 143506 79778 143534 80036
rect 143598 79937 143626 80036
rect 143584 79928 143640 79937
rect 143584 79863 143640 79872
rect 143690 79778 143718 80036
rect 143782 79835 143810 80036
rect 143874 79966 143902 80036
rect 143862 79960 143914 79966
rect 143862 79902 143914 79908
rect 143506 79750 143580 79778
rect 143138 79716 143212 79744
rect 142816 79558 142844 79716
rect 142804 79552 142856 79558
rect 142804 79494 142856 79500
rect 142724 79206 142936 79234
rect 142804 79144 142856 79150
rect 142804 79086 142856 79092
rect 142816 75682 142844 79086
rect 142804 75676 142856 75682
rect 142804 75618 142856 75624
rect 142908 75426 142936 79206
rect 142816 75398 142936 75426
rect 142712 75200 142764 75206
rect 142712 75142 142764 75148
rect 142724 68882 142752 75142
rect 142816 71262 142844 75398
rect 142896 75268 142948 75274
rect 142896 75210 142948 75216
rect 142804 71256 142856 71262
rect 142804 71198 142856 71204
rect 142712 68876 142764 68882
rect 142712 68818 142764 68824
rect 142710 68776 142766 68785
rect 142710 68711 142766 68720
rect 142724 68105 142752 68711
rect 142710 68096 142766 68105
rect 142710 68031 142766 68040
rect 142620 67516 142672 67522
rect 142620 67458 142672 67464
rect 142540 65470 142752 65498
rect 142528 65408 142580 65414
rect 142528 65350 142580 65356
rect 142540 49026 142568 65350
rect 142724 60734 142752 65470
rect 142816 65414 142844 71198
rect 142908 68814 142936 75210
rect 143000 69902 143028 79716
rect 143080 79552 143132 79558
rect 143080 79494 143132 79500
rect 143092 74526 143120 79494
rect 143184 75206 143212 79716
rect 143264 79620 143316 79626
rect 143264 79562 143316 79568
rect 143172 75200 143224 75206
rect 143172 75142 143224 75148
rect 143276 75138 143304 79562
rect 143368 75274 143396 79750
rect 143446 79656 143502 79665
rect 143446 79591 143502 79600
rect 143356 75268 143408 75274
rect 143356 75210 143408 75216
rect 143264 75132 143316 75138
rect 143264 75074 143316 75080
rect 143080 74520 143132 74526
rect 143080 74462 143132 74468
rect 143460 73098 143488 79591
rect 143552 79150 143580 79750
rect 143644 79750 143718 79778
rect 143768 79826 143824 79835
rect 143966 79801 143994 80036
rect 144058 79966 144086 80036
rect 144046 79960 144098 79966
rect 144046 79902 144098 79908
rect 144150 79898 144178 80036
rect 144138 79892 144190 79898
rect 144138 79834 144190 79840
rect 144046 79824 144098 79830
rect 143768 79761 143824 79770
rect 143952 79792 144008 79801
rect 143644 79608 143672 79750
rect 144098 79772 144178 79778
rect 144046 79766 144178 79772
rect 144058 79750 144178 79766
rect 143952 79727 144008 79736
rect 143908 79688 143960 79694
rect 144150 79642 144178 79750
rect 144242 79744 144270 80036
rect 144334 79966 144362 80036
rect 144426 79966 144454 80036
rect 144518 79966 144546 80036
rect 144610 79966 144638 80036
rect 144702 79966 144730 80036
rect 144322 79960 144374 79966
rect 144322 79902 144374 79908
rect 144414 79960 144466 79966
rect 144414 79902 144466 79908
rect 144506 79960 144558 79966
rect 144506 79902 144558 79908
rect 144598 79960 144650 79966
rect 144598 79902 144650 79908
rect 144690 79960 144742 79966
rect 144690 79902 144742 79908
rect 144368 79824 144420 79830
rect 144368 79766 144420 79772
rect 144460 79824 144512 79830
rect 144794 79812 144822 80036
rect 144886 79966 144914 80036
rect 144874 79960 144926 79966
rect 144874 79902 144926 79908
rect 144794 79801 144868 79812
rect 144794 79792 144882 79801
rect 144794 79784 144826 79792
rect 144460 79766 144512 79772
rect 144242 79716 144316 79744
rect 144288 79665 144316 79716
rect 143908 79630 143960 79636
rect 143816 79620 143868 79626
rect 143644 79580 143764 79608
rect 143540 79144 143592 79150
rect 143540 79086 143592 79092
rect 143538 78976 143594 78985
rect 143538 78911 143594 78920
rect 143552 78334 143580 78911
rect 143632 78736 143684 78742
rect 143632 78678 143684 78684
rect 143540 78328 143592 78334
rect 143540 78270 143592 78276
rect 143448 73092 143500 73098
rect 143448 73034 143500 73040
rect 142988 69896 143040 69902
rect 142988 69838 143040 69844
rect 142896 68808 142948 68814
rect 142896 68750 142948 68756
rect 142804 65408 142856 65414
rect 142804 65350 142856 65356
rect 142724 60706 142844 60734
rect 142528 49020 142580 49026
rect 142528 48962 142580 48968
rect 142816 8294 142844 60706
rect 142804 8288 142856 8294
rect 142804 8230 142856 8236
rect 142356 6886 142476 6914
rect 142356 4146 142384 6886
rect 142344 4140 142396 4146
rect 142344 4082 142396 4088
rect 141516 3528 141568 3534
rect 142908 3482 142936 68750
rect 143000 66162 143028 69838
rect 142988 66156 143040 66162
rect 142988 66098 143040 66104
rect 143552 11762 143580 78270
rect 143644 75018 143672 78678
rect 143736 75154 143764 79580
rect 143816 79562 143868 79568
rect 143828 77926 143856 79562
rect 143816 77920 143868 77926
rect 143816 77862 143868 77868
rect 143920 75274 143948 79630
rect 144000 79620 144052 79626
rect 144000 79562 144052 79568
rect 144104 79614 144178 79642
rect 144274 79656 144330 79665
rect 143908 75268 143960 75274
rect 143908 75210 143960 75216
rect 143736 75126 143948 75154
rect 143644 74990 143856 75018
rect 143724 74928 143776 74934
rect 143724 74870 143776 74876
rect 143736 51746 143764 74870
rect 143828 63442 143856 74990
rect 143920 69018 143948 75126
rect 143908 69012 143960 69018
rect 143908 68954 143960 68960
rect 143816 63436 143868 63442
rect 143816 63378 143868 63384
rect 143920 60734 143948 68954
rect 144012 68542 144040 79562
rect 144104 77722 144132 79614
rect 144274 79591 144330 79600
rect 144184 79552 144236 79558
rect 144184 79494 144236 79500
rect 144092 77716 144144 77722
rect 144092 77658 144144 77664
rect 144092 75268 144144 75274
rect 144092 75210 144144 75216
rect 144104 68746 144132 75210
rect 144196 75041 144224 79494
rect 144380 79472 144408 79766
rect 144288 79444 144408 79472
rect 144288 78742 144316 79444
rect 144366 79384 144422 79393
rect 144366 79319 144422 79328
rect 144276 78736 144328 78742
rect 144276 78678 144328 78684
rect 144380 76838 144408 79319
rect 144472 78033 144500 79766
rect 144826 79727 144882 79736
rect 144978 79744 145006 80036
rect 145070 79971 145098 80036
rect 145056 79962 145112 79971
rect 145056 79897 145112 79906
rect 145162 79744 145190 80036
rect 145254 79971 145282 80036
rect 145240 79962 145296 79971
rect 145240 79897 145296 79906
rect 145346 79898 145374 80036
rect 145334 79892 145386 79898
rect 145334 79834 145386 79840
rect 145438 79744 145466 80036
rect 145530 79898 145558 80036
rect 145622 79898 145650 80036
rect 145518 79892 145570 79898
rect 145518 79834 145570 79840
rect 145610 79892 145662 79898
rect 145610 79834 145662 79840
rect 145564 79756 145616 79762
rect 144978 79716 145052 79744
rect 145162 79716 145328 79744
rect 145438 79716 145512 79744
rect 144552 79688 144604 79694
rect 144550 79656 144552 79665
rect 144604 79656 144606 79665
rect 144550 79591 144606 79600
rect 144644 79620 144696 79626
rect 144644 79562 144696 79568
rect 144920 79620 144972 79626
rect 144920 79562 144972 79568
rect 144550 79520 144606 79529
rect 144550 79455 144606 79464
rect 144564 78742 144592 79455
rect 144552 78736 144604 78742
rect 144552 78678 144604 78684
rect 144458 78024 144514 78033
rect 144458 77959 144514 77968
rect 144460 77920 144512 77926
rect 144656 77897 144684 79562
rect 144734 79520 144790 79529
rect 144734 79455 144790 79464
rect 144748 79014 144776 79455
rect 144932 79150 144960 79562
rect 144920 79144 144972 79150
rect 144920 79086 144972 79092
rect 144736 79008 144788 79014
rect 144736 78950 144788 78956
rect 144460 77862 144512 77868
rect 144642 77888 144698 77897
rect 144368 76832 144420 76838
rect 144368 76774 144420 76780
rect 144380 76022 144408 76774
rect 144368 76016 144420 76022
rect 144368 75958 144420 75964
rect 144182 75032 144238 75041
rect 144182 74967 144238 74976
rect 144196 70394 144224 74967
rect 144472 70394 144500 77862
rect 144642 77823 144698 77832
rect 144748 74934 144776 78950
rect 144920 78736 144972 78742
rect 144920 78678 144972 78684
rect 144932 77602 144960 78678
rect 145024 78674 145052 79716
rect 145102 79520 145158 79529
rect 145102 79455 145158 79464
rect 145012 78668 145064 78674
rect 145012 78610 145064 78616
rect 144840 77574 144960 77602
rect 145012 77580 145064 77586
rect 144840 75818 144868 77574
rect 145012 77522 145064 77528
rect 144828 75812 144880 75818
rect 144828 75754 144880 75760
rect 144840 75546 144868 75754
rect 144828 75540 144880 75546
rect 144828 75482 144880 75488
rect 144736 74928 144788 74934
rect 144736 74870 144788 74876
rect 144196 70366 144316 70394
rect 144472 70366 144868 70394
rect 144092 68740 144144 68746
rect 144092 68682 144144 68688
rect 144000 68536 144052 68542
rect 144000 68478 144052 68484
rect 144012 66570 144040 68478
rect 144104 67658 144132 68682
rect 144092 67652 144144 67658
rect 144092 67594 144144 67600
rect 144000 66564 144052 66570
rect 144000 66506 144052 66512
rect 143920 60706 144224 60734
rect 143724 51740 143776 51746
rect 143724 51682 143776 51688
rect 144196 25702 144224 60706
rect 144288 33794 144316 70366
rect 144368 67652 144420 67658
rect 144368 67594 144420 67600
rect 144380 48278 144408 67594
rect 144368 48272 144420 48278
rect 144368 48214 144420 48220
rect 144276 33788 144328 33794
rect 144276 33730 144328 33736
rect 144184 25696 144236 25702
rect 144184 25638 144236 25644
rect 144840 19990 144868 70366
rect 145024 49026 145052 77522
rect 145116 77246 145144 79455
rect 145300 78962 145328 79716
rect 145208 78934 145328 78962
rect 145104 77240 145156 77246
rect 145104 77182 145156 77188
rect 145208 75274 145236 78934
rect 145288 78192 145340 78198
rect 145288 78134 145340 78140
rect 145196 75268 145248 75274
rect 145196 75210 145248 75216
rect 145208 75002 145236 75210
rect 145196 74996 145248 75002
rect 145196 74938 145248 74944
rect 145300 60734 145328 78134
rect 145484 75342 145512 79716
rect 145714 79744 145742 80036
rect 145564 79698 145616 79704
rect 145668 79716 145742 79744
rect 145806 79744 145834 80036
rect 145898 79812 145926 80036
rect 145990 79971 146018 80036
rect 145976 79962 146032 79971
rect 146082 79966 146110 80036
rect 146174 79971 146202 80036
rect 145976 79897 146032 79906
rect 146070 79960 146122 79966
rect 146070 79902 146122 79908
rect 146160 79962 146216 79971
rect 146266 79966 146294 80036
rect 146358 79966 146386 80036
rect 146082 79830 146110 79902
rect 146160 79897 146216 79906
rect 146254 79960 146306 79966
rect 146254 79902 146306 79908
rect 146346 79960 146398 79966
rect 146346 79902 146398 79908
rect 146450 79898 146478 80036
rect 146542 79966 146570 80036
rect 146634 79966 146662 80036
rect 146726 79971 146754 80036
rect 146530 79960 146582 79966
rect 146530 79902 146582 79908
rect 146622 79960 146674 79966
rect 146622 79902 146674 79908
rect 146712 79962 146768 79971
rect 146438 79892 146490 79898
rect 146712 79897 146768 79906
rect 146438 79834 146490 79840
rect 146070 79824 146122 79830
rect 145898 79801 145972 79812
rect 145898 79792 145986 79801
rect 145898 79784 145930 79792
rect 145806 79716 145880 79744
rect 146070 79766 146122 79772
rect 146818 79778 146846 80036
rect 146910 79898 146938 80036
rect 147002 79966 147030 80036
rect 146990 79960 147042 79966
rect 146990 79902 147042 79908
rect 146898 79892 146950 79898
rect 146898 79834 146950 79840
rect 145930 79727 145986 79736
rect 146208 79756 146260 79762
rect 145576 77586 145604 79698
rect 145668 79676 145696 79716
rect 145668 79648 145788 79676
rect 145656 79552 145708 79558
rect 145656 79494 145708 79500
rect 145668 78130 145696 79494
rect 145656 78124 145708 78130
rect 145656 78066 145708 78072
rect 145564 77580 145616 77586
rect 145564 77522 145616 77528
rect 145472 75336 145524 75342
rect 145472 75278 145524 75284
rect 145484 70394 145512 75278
rect 145484 70366 145604 70394
rect 145116 60706 145328 60734
rect 145116 55894 145144 60706
rect 145104 55888 145156 55894
rect 145104 55830 145156 55836
rect 145012 49020 145064 49026
rect 145012 48962 145064 48968
rect 145576 38214 145604 70366
rect 145668 46238 145696 78066
rect 145760 76770 145788 79648
rect 145852 78266 145880 79716
rect 146208 79698 146260 79704
rect 146576 79756 146628 79762
rect 146818 79750 146892 79778
rect 146576 79698 146628 79704
rect 145932 79688 145984 79694
rect 145932 79630 145984 79636
rect 145840 78260 145892 78266
rect 145840 78202 145892 78208
rect 145944 77178 145972 79630
rect 146024 79620 146076 79626
rect 146024 79562 146076 79568
rect 146036 79150 146064 79562
rect 146114 79520 146170 79529
rect 146114 79455 146170 79464
rect 146024 79144 146076 79150
rect 146024 79086 146076 79092
rect 146036 77450 146064 79086
rect 146128 78878 146156 79455
rect 146116 78872 146168 78878
rect 146116 78814 146168 78820
rect 146024 77444 146076 77450
rect 146024 77386 146076 77392
rect 146024 77240 146076 77246
rect 146024 77182 146076 77188
rect 145932 77172 145984 77178
rect 145932 77114 145984 77120
rect 145748 76764 145800 76770
rect 145748 76706 145800 76712
rect 145748 75268 145800 75274
rect 145748 75210 145800 75216
rect 145760 53106 145788 75210
rect 146036 63646 146064 77182
rect 146024 63640 146076 63646
rect 146024 63582 146076 63588
rect 146128 60734 146156 78814
rect 146220 76673 146248 79698
rect 146300 79620 146352 79626
rect 146352 79580 146432 79608
rect 146300 79562 146352 79568
rect 146300 79484 146352 79490
rect 146300 79426 146352 79432
rect 146312 79286 146340 79426
rect 146404 79286 146432 79580
rect 146484 79552 146536 79558
rect 146484 79494 146536 79500
rect 146300 79280 146352 79286
rect 146300 79222 146352 79228
rect 146392 79280 146444 79286
rect 146392 79222 146444 79228
rect 146312 77518 146340 79222
rect 146300 77512 146352 77518
rect 146300 77454 146352 77460
rect 146206 76664 146262 76673
rect 146206 76599 146262 76608
rect 146300 76016 146352 76022
rect 146300 75958 146352 75964
rect 146036 60706 146156 60734
rect 145748 53100 145800 53106
rect 145748 53042 145800 53048
rect 145656 46232 145708 46238
rect 145656 46174 145708 46180
rect 145564 38208 145616 38214
rect 145564 38150 145616 38156
rect 144920 25696 144972 25702
rect 144920 25638 144972 25644
rect 144828 19984 144880 19990
rect 144828 19926 144880 19932
rect 144932 16574 144960 25638
rect 146036 25566 146064 60706
rect 146024 25560 146076 25566
rect 146024 25502 146076 25508
rect 146312 16574 146340 75958
rect 146496 75614 146524 79494
rect 146484 75608 146536 75614
rect 146484 75550 146536 75556
rect 146588 75070 146616 79698
rect 146666 79656 146722 79665
rect 146666 79591 146722 79600
rect 146680 75478 146708 79591
rect 146864 79506 146892 79750
rect 147094 79608 147122 80036
rect 147186 79898 147214 80036
rect 147278 79937 147306 80036
rect 147264 79928 147320 79937
rect 147174 79892 147226 79898
rect 147370 79898 147398 80036
rect 147462 79898 147490 80036
rect 147264 79863 147320 79872
rect 147358 79892 147410 79898
rect 147174 79834 147226 79840
rect 147358 79834 147410 79840
rect 147450 79892 147502 79898
rect 147450 79834 147502 79840
rect 147554 79744 147582 80036
rect 147646 79966 147674 80036
rect 147634 79960 147686 79966
rect 147634 79902 147686 79908
rect 147634 79824 147686 79830
rect 147508 79716 147582 79744
rect 147632 79792 147634 79801
rect 147686 79792 147688 79801
rect 147632 79727 147688 79736
rect 147738 79744 147766 80036
rect 147830 79971 147858 80036
rect 147816 79962 147872 79971
rect 147816 79897 147872 79906
rect 147922 79744 147950 80036
rect 148014 79898 148042 80036
rect 148002 79892 148054 79898
rect 148002 79834 148054 79840
rect 148106 79744 148134 80036
rect 148198 79971 148226 80036
rect 148184 79962 148240 79971
rect 148290 79966 148318 80036
rect 148382 79966 148410 80036
rect 148184 79897 148240 79906
rect 148278 79960 148330 79966
rect 148278 79902 148330 79908
rect 148370 79960 148422 79966
rect 148370 79902 148422 79908
rect 148232 79824 148284 79830
rect 148232 79766 148284 79772
rect 147738 79716 147812 79744
rect 147922 79716 147996 79744
rect 147218 79656 147274 79665
rect 147094 79580 147168 79608
rect 147218 79591 147220 79600
rect 146772 79478 146892 79506
rect 147036 79484 147088 79490
rect 146772 76974 146800 79478
rect 147036 79426 147088 79432
rect 146852 77512 146904 77518
rect 147048 77489 147076 79426
rect 146852 77454 146904 77460
rect 147034 77480 147090 77489
rect 146760 76968 146812 76974
rect 146760 76910 146812 76916
rect 146772 76566 146800 76910
rect 146760 76560 146812 76566
rect 146760 76502 146812 76508
rect 146668 75472 146720 75478
rect 146668 75414 146720 75420
rect 146576 75064 146628 75070
rect 146576 75006 146628 75012
rect 146588 72486 146616 75006
rect 146576 72480 146628 72486
rect 146576 72422 146628 72428
rect 146864 64190 146892 77454
rect 146944 77444 146996 77450
rect 147034 77415 147090 77424
rect 146944 77386 146996 77392
rect 146852 64184 146904 64190
rect 146852 64126 146904 64132
rect 144932 16546 145512 16574
rect 146312 16546 146892 16574
rect 143540 11756 143592 11762
rect 143540 11698 143592 11704
rect 144736 11756 144788 11762
rect 144736 11698 144788 11704
rect 143540 8288 143592 8294
rect 143540 8230 143592 8236
rect 141516 3470 141568 3476
rect 142448 3454 142936 3482
rect 141424 3188 141476 3194
rect 141424 3130 141476 3136
rect 142448 480 142476 3454
rect 143552 480 143580 8230
rect 144748 480 144776 11698
rect 134126 354 134238 480
rect 133984 326 134238 354
rect 134126 -960 134238 326
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145484 354 145512 16546
rect 146864 3482 146892 16546
rect 146956 3874 146984 77386
rect 147140 77042 147168 79580
rect 147272 79591 147274 79600
rect 147220 79562 147272 79568
rect 147232 77294 147260 79562
rect 147404 79552 147456 79558
rect 147404 79494 147456 79500
rect 147232 77266 147352 77294
rect 147128 77036 147180 77042
rect 147128 76978 147180 76984
rect 147036 75540 147088 75546
rect 147036 75482 147088 75488
rect 146944 3868 146996 3874
rect 146944 3810 146996 3816
rect 147048 3670 147076 75482
rect 147140 71126 147168 76978
rect 147324 76634 147352 77266
rect 147312 76628 147364 76634
rect 147312 76570 147364 76576
rect 147128 71120 147180 71126
rect 147128 71062 147180 71068
rect 147126 67688 147182 67697
rect 147126 67623 147182 67632
rect 147140 5250 147168 67623
rect 147220 66564 147272 66570
rect 147220 66506 147272 66512
rect 147232 16574 147260 66506
rect 147416 49230 147444 79494
rect 147508 79422 147536 79716
rect 147784 79676 147812 79716
rect 147678 79656 147734 79665
rect 147784 79648 147904 79676
rect 147678 79591 147734 79600
rect 147588 79552 147640 79558
rect 147588 79494 147640 79500
rect 147496 79416 147548 79422
rect 147496 79358 147548 79364
rect 147508 75274 147536 79358
rect 147600 77353 147628 79494
rect 147692 78946 147720 79591
rect 147772 79552 147824 79558
rect 147876 79529 147904 79648
rect 147772 79494 147824 79500
rect 147862 79520 147918 79529
rect 147784 79354 147812 79494
rect 147862 79455 147918 79464
rect 147862 79384 147918 79393
rect 147772 79348 147824 79354
rect 147862 79319 147918 79328
rect 147772 79290 147824 79296
rect 147680 78940 147732 78946
rect 147680 78882 147732 78888
rect 147586 77344 147642 77353
rect 147586 77279 147642 77288
rect 147496 75268 147548 75274
rect 147496 75210 147548 75216
rect 147404 49224 147456 49230
rect 147404 49166 147456 49172
rect 147692 48906 147720 78882
rect 147784 49094 147812 79290
rect 147876 74322 147904 79319
rect 147968 78674 147996 79716
rect 148060 79716 148134 79744
rect 147956 78668 148008 78674
rect 147956 78610 148008 78616
rect 147956 78396 148008 78402
rect 147956 78338 148008 78344
rect 147864 74316 147916 74322
rect 147864 74258 147916 74264
rect 147864 73024 147916 73030
rect 147864 72966 147916 72972
rect 147876 66910 147904 72966
rect 147968 71534 147996 78338
rect 148060 75206 148088 79716
rect 148138 79384 148194 79393
rect 148138 79319 148194 79328
rect 148048 75200 148100 75206
rect 148048 75142 148100 75148
rect 148152 72622 148180 79319
rect 148140 72616 148192 72622
rect 148140 72558 148192 72564
rect 147956 71528 148008 71534
rect 147956 71470 148008 71476
rect 148244 71466 148272 79766
rect 148324 79756 148376 79762
rect 148474 79744 148502 80036
rect 148566 79937 148594 80036
rect 148552 79928 148608 79937
rect 148552 79863 148608 79872
rect 148658 79778 148686 80036
rect 148750 79971 148778 80036
rect 148736 79962 148792 79971
rect 148736 79897 148792 79906
rect 148842 79830 148870 80036
rect 148830 79824 148882 79830
rect 148658 79750 148732 79778
rect 148830 79766 148882 79772
rect 148474 79716 148548 79744
rect 148324 79698 148376 79704
rect 148336 79490 148364 79698
rect 148414 79656 148470 79665
rect 148414 79591 148470 79600
rect 148324 79484 148376 79490
rect 148324 79426 148376 79432
rect 148324 78668 148376 78674
rect 148324 78610 148376 78616
rect 148336 77294 148364 78610
rect 148428 77722 148456 79591
rect 148416 77716 148468 77722
rect 148416 77658 148468 77664
rect 148336 77266 148456 77294
rect 148324 77172 148376 77178
rect 148324 77114 148376 77120
rect 148232 71460 148284 71466
rect 148232 71402 148284 71408
rect 147864 66904 147916 66910
rect 147864 66846 147916 66852
rect 147772 49088 147824 49094
rect 147772 49030 147824 49036
rect 147692 48878 147812 48906
rect 147680 48272 147732 48278
rect 147680 48214 147732 48220
rect 147692 16574 147720 48214
rect 147784 47734 147812 48878
rect 147772 47728 147824 47734
rect 147772 47670 147824 47676
rect 147232 16546 147352 16574
rect 147692 16546 147904 16574
rect 147140 5222 147260 5250
rect 147036 3664 147088 3670
rect 147036 3606 147088 3612
rect 147232 3534 147260 5222
rect 147220 3528 147272 3534
rect 146864 3454 147168 3482
rect 147220 3470 147272 3476
rect 147140 480 147168 3454
rect 147324 3398 147352 16546
rect 147312 3392 147364 3398
rect 147312 3334 147364 3340
rect 145902 354 146014 480
rect 145484 326 146014 354
rect 145902 -960 146014 326
rect 147098 -960 147210 480
rect 147876 354 147904 16546
rect 148336 3466 148364 77114
rect 148428 72758 148456 77266
rect 148520 73030 148548 79716
rect 148704 79642 148732 79750
rect 148934 79744 148962 80036
rect 149026 79812 149054 80036
rect 149118 79966 149146 80036
rect 149106 79960 149158 79966
rect 149210 79937 149238 80036
rect 149302 79966 149330 80036
rect 149290 79960 149342 79966
rect 149106 79902 149158 79908
rect 149196 79928 149252 79937
rect 149290 79902 149342 79908
rect 149196 79863 149252 79872
rect 149152 79824 149204 79830
rect 149026 79784 149100 79812
rect 148934 79716 149008 79744
rect 148704 79614 148916 79642
rect 148690 79520 148746 79529
rect 148690 79455 148746 79464
rect 148784 79484 148836 79490
rect 148600 79416 148652 79422
rect 148600 79358 148652 79364
rect 148612 77489 148640 79358
rect 148704 79082 148732 79455
rect 148784 79426 148836 79432
rect 148692 79076 148744 79082
rect 148692 79018 148744 79024
rect 148704 77518 148732 79018
rect 148692 77512 148744 77518
rect 148598 77480 148654 77489
rect 148692 77454 148744 77460
rect 148598 77415 148654 77424
rect 148692 74316 148744 74322
rect 148692 74258 148744 74264
rect 148508 73024 148560 73030
rect 148508 72966 148560 72972
rect 148416 72752 148468 72758
rect 148416 72694 148468 72700
rect 148600 72616 148652 72622
rect 148600 72558 148652 72564
rect 148508 71460 148560 71466
rect 148508 71402 148560 71408
rect 148520 69578 148548 71402
rect 148612 69698 148640 72558
rect 148600 69692 148652 69698
rect 148600 69634 148652 69640
rect 148520 69550 148640 69578
rect 148506 69456 148562 69465
rect 148506 69391 148562 69400
rect 148416 63436 148468 63442
rect 148416 63378 148468 63384
rect 148324 3460 148376 3466
rect 148324 3402 148376 3408
rect 148428 3058 148456 63378
rect 148520 32706 148548 69391
rect 148612 41070 148640 69550
rect 148704 58954 148732 74258
rect 148796 70394 148824 79426
rect 148888 77353 148916 79614
rect 148980 77625 149008 79716
rect 149072 78577 149100 79784
rect 149152 79766 149204 79772
rect 149244 79824 149296 79830
rect 149244 79766 149296 79772
rect 149058 78568 149114 78577
rect 149058 78503 149114 78512
rect 149164 78402 149192 79766
rect 149256 79354 149284 79766
rect 149394 79744 149422 80036
rect 149348 79716 149422 79744
rect 149244 79348 149296 79354
rect 149244 79290 149296 79296
rect 149348 78713 149376 79716
rect 149486 79676 149514 80036
rect 149578 79744 149606 80036
rect 149670 79898 149698 80036
rect 149762 79966 149790 80036
rect 149750 79960 149802 79966
rect 149750 79902 149802 79908
rect 149854 79898 149882 80036
rect 149658 79892 149710 79898
rect 149658 79834 149710 79840
rect 149842 79892 149894 79898
rect 149842 79834 149894 79840
rect 149946 79744 149974 80036
rect 150038 79966 150066 80036
rect 150026 79960 150078 79966
rect 150026 79902 150078 79908
rect 150130 79898 150158 80036
rect 150118 79892 150170 79898
rect 150118 79834 150170 79840
rect 150222 79744 150250 80036
rect 150314 79778 150342 80036
rect 150406 79966 150434 80036
rect 150394 79960 150446 79966
rect 150394 79902 150446 79908
rect 150498 79898 150526 80036
rect 150590 79971 150618 80036
rect 150576 79962 150632 79971
rect 150682 79966 150710 80036
rect 150486 79892 150538 79898
rect 150576 79897 150632 79906
rect 150670 79960 150722 79966
rect 150670 79902 150722 79908
rect 150774 79903 150802 80036
rect 150486 79834 150538 79840
rect 150760 79894 150816 79903
rect 150624 79824 150676 79830
rect 150760 79829 150816 79838
rect 150314 79750 150480 79778
rect 150866 79778 150894 80036
rect 150624 79766 150676 79772
rect 149578 79716 149652 79744
rect 149946 79716 150112 79744
rect 149440 79648 149514 79676
rect 149334 78704 149390 78713
rect 149334 78639 149390 78648
rect 149152 78396 149204 78402
rect 149152 78338 149204 78344
rect 149348 78282 149376 78639
rect 149072 78254 149376 78282
rect 148966 77616 149022 77625
rect 148966 77551 149022 77560
rect 148968 77512 149020 77518
rect 148968 77454 149020 77460
rect 148874 77344 148930 77353
rect 148874 77279 148930 77288
rect 148796 70366 148916 70394
rect 148888 70145 148916 70366
rect 148874 70136 148930 70145
rect 148874 70071 148930 70080
rect 148888 69465 148916 70071
rect 148874 69456 148930 69465
rect 148874 69391 148930 69400
rect 148980 61674 149008 77454
rect 148968 61668 149020 61674
rect 148968 61610 149020 61616
rect 148692 58948 148744 58954
rect 148692 58890 148744 58896
rect 149072 42362 149100 78254
rect 149440 77330 149468 79648
rect 149520 79552 149572 79558
rect 149520 79494 149572 79500
rect 149256 77302 149468 77330
rect 149152 74180 149204 74186
rect 149152 74122 149204 74128
rect 149164 74089 149192 74122
rect 149150 74080 149206 74089
rect 149150 74015 149206 74024
rect 149256 73914 149284 77302
rect 149336 75132 149388 75138
rect 149336 75074 149388 75080
rect 149244 73908 149296 73914
rect 149244 73850 149296 73856
rect 149348 70394 149376 75074
rect 149532 71233 149560 79494
rect 149624 77353 149652 79716
rect 150084 79665 150112 79716
rect 150176 79716 150250 79744
rect 150070 79656 150126 79665
rect 149796 79620 149848 79626
rect 149796 79562 149848 79568
rect 149888 79620 149940 79626
rect 149888 79562 149940 79568
rect 149980 79620 150032 79626
rect 150070 79591 150126 79600
rect 149980 79562 150032 79568
rect 149704 79484 149756 79490
rect 149704 79426 149756 79432
rect 149610 77344 149666 77353
rect 149610 77279 149666 77288
rect 149716 76906 149744 79426
rect 149704 76900 149756 76906
rect 149704 76842 149756 76848
rect 149716 75342 149744 76842
rect 149704 75336 149756 75342
rect 149704 75278 149756 75284
rect 149612 73160 149664 73166
rect 149612 73102 149664 73108
rect 149518 71224 149574 71233
rect 149518 71159 149574 71168
rect 149532 70394 149560 71159
rect 149164 70366 149376 70394
rect 149440 70366 149560 70394
rect 149164 67386 149192 70366
rect 149152 67380 149204 67386
rect 149152 67322 149204 67328
rect 149164 67114 149192 67322
rect 149152 67108 149204 67114
rect 149152 67050 149204 67056
rect 149440 65686 149468 70366
rect 149428 65680 149480 65686
rect 149428 65622 149480 65628
rect 149624 64326 149652 73102
rect 149808 71738 149836 79562
rect 149900 73166 149928 79562
rect 149992 75138 150020 79562
rect 150072 79552 150124 79558
rect 150072 79494 150124 79500
rect 150084 77353 150112 79494
rect 150070 77344 150126 77353
rect 150070 77279 150126 77288
rect 149980 75132 150032 75138
rect 149980 75074 150032 75080
rect 150176 73930 150204 79716
rect 150348 79688 150400 79694
rect 150254 79656 150310 79665
rect 150348 79630 150400 79636
rect 150254 79591 150310 79600
rect 150268 74066 150296 79591
rect 150360 77489 150388 79630
rect 150452 78577 150480 79750
rect 150438 78568 150494 78577
rect 150438 78503 150494 78512
rect 150346 77480 150402 77489
rect 150346 77415 150402 77424
rect 150532 76696 150584 76702
rect 150532 76638 150584 76644
rect 150440 76424 150492 76430
rect 150440 76366 150492 76372
rect 150268 74038 150388 74066
rect 149980 73908 150032 73914
rect 149980 73850 150032 73856
rect 150084 73902 150204 73930
rect 149888 73160 149940 73166
rect 149888 73102 149940 73108
rect 149796 71732 149848 71738
rect 149796 71674 149848 71680
rect 149808 70650 149836 71674
rect 149796 70644 149848 70650
rect 149796 70586 149848 70592
rect 149702 67552 149758 67561
rect 149702 67487 149758 67496
rect 149612 64320 149664 64326
rect 149612 64262 149664 64268
rect 149060 42356 149112 42362
rect 149060 42298 149112 42304
rect 148600 41064 148652 41070
rect 148600 41006 148652 41012
rect 148508 32700 148560 32706
rect 148508 32642 148560 32648
rect 149716 4146 149744 67487
rect 149888 67108 149940 67114
rect 149888 67050 149940 67056
rect 149796 63640 149848 63646
rect 149796 63582 149848 63588
rect 149704 4140 149756 4146
rect 149704 4082 149756 4088
rect 149808 3874 149836 63582
rect 149900 7886 149928 67050
rect 149992 17474 150020 73850
rect 150084 71330 150112 73902
rect 150360 71641 150388 74038
rect 150346 71632 150402 71641
rect 150346 71567 150402 71576
rect 150164 71528 150216 71534
rect 150164 71470 150216 71476
rect 150072 71324 150124 71330
rect 150072 71266 150124 71272
rect 150084 29986 150112 71266
rect 150176 47666 150204 71470
rect 150256 70644 150308 70650
rect 150256 70586 150308 70592
rect 150268 49162 150296 70586
rect 150360 50386 150388 71567
rect 150348 50380 150400 50386
rect 150348 50322 150400 50328
rect 150256 49156 150308 49162
rect 150256 49098 150308 49104
rect 150164 47660 150216 47666
rect 150164 47602 150216 47608
rect 150452 39642 150480 76366
rect 150544 65890 150572 76638
rect 150636 67590 150664 79766
rect 150728 79750 150894 79778
rect 150728 77489 150756 79750
rect 150958 79676 150986 80036
rect 151050 79778 151078 80036
rect 151142 79898 151170 80036
rect 151130 79892 151182 79898
rect 151130 79834 151182 79840
rect 151050 79750 151124 79778
rect 150912 79648 150986 79676
rect 150806 79520 150862 79529
rect 150806 79455 150862 79464
rect 150714 77480 150770 77489
rect 150714 77415 150770 77424
rect 150820 70394 150848 79455
rect 150912 77654 150940 79648
rect 151096 79608 151124 79750
rect 151234 79744 151262 80036
rect 151004 79580 151124 79608
rect 151188 79716 151262 79744
rect 151326 79744 151354 80036
rect 151418 79812 151446 80036
rect 151510 79966 151538 80036
rect 151498 79960 151550 79966
rect 151498 79902 151550 79908
rect 151602 79812 151630 80036
rect 151694 79966 151722 80036
rect 151786 79966 151814 80036
rect 151682 79960 151734 79966
rect 151682 79902 151734 79908
rect 151774 79960 151826 79966
rect 151774 79902 151826 79908
rect 151418 79784 151492 79812
rect 151326 79716 151400 79744
rect 150900 77648 150952 77654
rect 150900 77590 150952 77596
rect 150900 72752 150952 72758
rect 150900 72694 150952 72700
rect 150912 71058 150940 72694
rect 150900 71052 150952 71058
rect 150900 70994 150952 71000
rect 150728 70366 150848 70394
rect 150728 69306 150756 70366
rect 151004 70038 151032 79580
rect 151082 78160 151138 78169
rect 151082 78095 151138 78104
rect 151096 75410 151124 78095
rect 151084 75404 151136 75410
rect 151084 75346 151136 75352
rect 151188 73953 151216 79716
rect 151266 79656 151322 79665
rect 151266 79591 151322 79600
rect 151280 78849 151308 79591
rect 151266 78840 151322 78849
rect 151266 78775 151322 78784
rect 151280 76430 151308 78775
rect 151268 76424 151320 76430
rect 151268 76366 151320 76372
rect 151174 73944 151230 73953
rect 151174 73879 151230 73888
rect 151188 71890 151216 73879
rect 151188 71862 151308 71890
rect 151174 71768 151230 71777
rect 151174 71703 151230 71712
rect 150992 70032 151044 70038
rect 150992 69974 151044 69980
rect 151004 69834 151032 69974
rect 150992 69828 151044 69834
rect 150992 69770 151044 69776
rect 151188 69714 151216 71703
rect 151280 70394 151308 71862
rect 151372 71777 151400 79716
rect 151464 79665 151492 79784
rect 151556 79784 151630 79812
rect 151878 79801 151906 80036
rect 151970 79966 151998 80036
rect 152062 79966 152090 80036
rect 151958 79960 152010 79966
rect 151958 79902 152010 79908
rect 152050 79960 152102 79966
rect 152050 79902 152102 79908
rect 152004 79824 152056 79830
rect 151864 79792 151920 79801
rect 151450 79656 151506 79665
rect 151450 79591 151506 79600
rect 151452 79484 151504 79490
rect 151452 79426 151504 79432
rect 151358 71768 151414 71777
rect 151358 71703 151414 71712
rect 151464 71194 151492 79426
rect 151556 76537 151584 79784
rect 152004 79766 152056 79772
rect 151864 79727 151920 79736
rect 151636 79688 151688 79694
rect 151636 79630 151688 79636
rect 151820 79688 151872 79694
rect 151820 79630 151872 79636
rect 151648 76702 151676 79630
rect 151728 79484 151780 79490
rect 151728 79426 151780 79432
rect 151636 76696 151688 76702
rect 151636 76638 151688 76644
rect 151542 76528 151598 76537
rect 151542 76463 151598 76472
rect 151636 75064 151688 75070
rect 151636 75006 151688 75012
rect 151648 74050 151676 75006
rect 151740 74497 151768 79426
rect 151832 75070 151860 79630
rect 152016 76809 152044 79766
rect 152154 79744 152182 80036
rect 152246 79966 152274 80036
rect 152234 79960 152286 79966
rect 152234 79902 152286 79908
rect 152338 79898 152366 80036
rect 152326 79892 152378 79898
rect 152326 79834 152378 79840
rect 152278 79792 152334 79801
rect 152154 79716 152228 79744
rect 152430 79778 152458 80036
rect 152278 79727 152334 79736
rect 152384 79750 152458 79778
rect 152096 79620 152148 79626
rect 152096 79562 152148 79568
rect 152108 79218 152136 79562
rect 152096 79212 152148 79218
rect 152096 79154 152148 79160
rect 152200 76906 152228 79716
rect 152188 76900 152240 76906
rect 152188 76842 152240 76848
rect 152002 76800 152058 76809
rect 152002 76735 152058 76744
rect 151912 76696 151964 76702
rect 151912 76638 151964 76644
rect 151820 75064 151872 75070
rect 151820 75006 151872 75012
rect 151726 74488 151782 74497
rect 151726 74423 151782 74432
rect 151636 74044 151688 74050
rect 151636 73986 151688 73992
rect 151452 71188 151504 71194
rect 151452 71130 151504 71136
rect 151280 70366 151400 70394
rect 151372 69902 151400 70366
rect 151360 69896 151412 69902
rect 151360 69838 151412 69844
rect 151188 69686 151400 69714
rect 150728 69278 151216 69306
rect 151188 68649 151216 69278
rect 151174 68640 151230 68649
rect 151174 68575 151230 68584
rect 150624 67584 150676 67590
rect 150624 67526 150676 67532
rect 151084 67584 151136 67590
rect 151084 67526 151136 67532
rect 150636 67182 150664 67526
rect 150624 67176 150676 67182
rect 150624 67118 150676 67124
rect 150532 65884 150584 65890
rect 150532 65826 150584 65832
rect 150544 65482 150572 65826
rect 150532 65476 150584 65482
rect 150532 65418 150584 65424
rect 150440 39636 150492 39642
rect 150440 39578 150492 39584
rect 150072 29980 150124 29986
rect 150072 29922 150124 29928
rect 149980 17468 150032 17474
rect 149980 17410 150032 17416
rect 151096 10606 151124 67526
rect 151188 12034 151216 68575
rect 151268 65476 151320 65482
rect 151268 65418 151320 65424
rect 151280 16114 151308 65418
rect 151372 28558 151400 69686
rect 151464 43518 151492 71130
rect 151544 69828 151596 69834
rect 151544 69770 151596 69776
rect 151556 54670 151584 69770
rect 151648 58886 151676 73986
rect 151740 62966 151768 74423
rect 151924 67454 151952 76638
rect 152004 75200 152056 75206
rect 152004 75142 152056 75148
rect 152016 68921 152044 75142
rect 152292 73642 152320 79727
rect 152280 73636 152332 73642
rect 152280 73578 152332 73584
rect 152384 70394 152412 79750
rect 152522 79676 152550 80036
rect 152614 79966 152642 80036
rect 152602 79960 152654 79966
rect 152706 79937 152734 80036
rect 152602 79902 152654 79908
rect 152692 79928 152748 79937
rect 152692 79863 152748 79872
rect 152602 79824 152654 79830
rect 152600 79792 152602 79801
rect 152654 79792 152656 79801
rect 152798 79778 152826 80036
rect 152890 79966 152918 80036
rect 152878 79960 152930 79966
rect 152878 79902 152930 79908
rect 152982 79898 153010 80036
rect 152970 79892 153022 79898
rect 152970 79834 153022 79840
rect 153074 79778 153102 80036
rect 152798 79750 152964 79778
rect 152600 79727 152656 79736
rect 152476 79648 152550 79676
rect 152648 79688 152700 79694
rect 152476 76702 152504 79648
rect 152648 79630 152700 79636
rect 152740 79688 152792 79694
rect 152740 79630 152792 79636
rect 152832 79688 152884 79694
rect 152832 79630 152884 79636
rect 152556 76764 152608 76770
rect 152556 76706 152608 76712
rect 152464 76696 152516 76702
rect 152464 76638 152516 76644
rect 152568 75914 152596 76706
rect 152108 70366 152412 70394
rect 152476 75886 152596 75914
rect 152108 70310 152136 70366
rect 152096 70304 152148 70310
rect 152096 70246 152148 70252
rect 152002 68912 152058 68921
rect 152002 68847 152058 68856
rect 151912 67448 151964 67454
rect 151912 67390 151964 67396
rect 151728 62960 151780 62966
rect 151728 62902 151780 62908
rect 151636 58880 151688 58886
rect 151636 58822 151688 58828
rect 151544 54664 151596 54670
rect 151544 54606 151596 54612
rect 151452 43512 151504 43518
rect 151452 43454 151504 43460
rect 151360 28552 151412 28558
rect 151360 28494 151412 28500
rect 151268 16108 151320 16114
rect 151268 16050 151320 16056
rect 151176 12028 151228 12034
rect 151176 11970 151228 11976
rect 151084 10600 151136 10606
rect 151084 10542 151136 10548
rect 149888 7880 149940 7886
rect 149888 7822 149940 7828
rect 152476 3942 152504 75886
rect 152660 74526 152688 79630
rect 152752 77489 152780 79630
rect 152738 77480 152794 77489
rect 152738 77415 152794 77424
rect 152648 74520 152700 74526
rect 152648 74462 152700 74468
rect 152648 70304 152700 70310
rect 152648 70246 152700 70252
rect 152556 67448 152608 67454
rect 152556 67390 152608 67396
rect 152568 6594 152596 67390
rect 152660 13394 152688 70246
rect 152844 69873 152872 79630
rect 152936 78198 152964 79750
rect 153028 79750 153102 79778
rect 152924 78192 152976 78198
rect 152924 78134 152976 78140
rect 152924 78056 152976 78062
rect 152924 77998 152976 78004
rect 152936 74118 152964 77998
rect 153028 75206 153056 79750
rect 153166 79744 153194 80036
rect 153258 79966 153286 80036
rect 153246 79960 153298 79966
rect 153246 79902 153298 79908
rect 153350 79812 153378 80036
rect 153442 79966 153470 80036
rect 153534 79966 153562 80036
rect 153430 79960 153482 79966
rect 153430 79902 153482 79908
rect 153522 79960 153574 79966
rect 153522 79902 153574 79908
rect 153626 79812 153654 80036
rect 153718 79898 153746 80036
rect 153810 79966 153838 80036
rect 153798 79960 153850 79966
rect 153798 79902 153850 79908
rect 153902 79898 153930 80036
rect 153994 79966 154022 80036
rect 154086 79971 154114 80036
rect 153982 79960 154034 79966
rect 153982 79902 154034 79908
rect 154072 79962 154128 79971
rect 153706 79892 153758 79898
rect 153706 79834 153758 79840
rect 153890 79892 153942 79898
rect 154072 79897 154128 79906
rect 153890 79834 153942 79840
rect 153304 79801 153378 79812
rect 153290 79792 153378 79801
rect 153166 79716 153240 79744
rect 153346 79784 153378 79792
rect 153580 79784 153654 79812
rect 153290 79727 153346 79736
rect 153108 79620 153160 79626
rect 153108 79562 153160 79568
rect 153016 75200 153068 75206
rect 153016 75142 153068 75148
rect 152924 74112 152976 74118
rect 152924 74054 152976 74060
rect 152830 69864 152886 69873
rect 152830 69799 152886 69808
rect 152738 68912 152794 68921
rect 152738 68847 152794 68856
rect 152752 18834 152780 68847
rect 152844 32638 152872 69799
rect 152936 44878 152964 74054
rect 153016 73636 153068 73642
rect 153016 73578 153068 73584
rect 153028 70553 153056 73578
rect 153014 70544 153070 70553
rect 153014 70479 153070 70488
rect 152924 44872 152976 44878
rect 152924 44814 152976 44820
rect 153028 38146 153056 70479
rect 153120 64802 153148 79562
rect 153212 78062 153240 79716
rect 153384 79688 153436 79694
rect 153384 79630 153436 79636
rect 153474 79656 153530 79665
rect 153292 79484 153344 79490
rect 153292 79426 153344 79432
rect 153304 79257 153332 79426
rect 153290 79248 153346 79257
rect 153290 79183 153346 79192
rect 153200 78056 153252 78062
rect 153200 77998 153252 78004
rect 153304 77874 153332 79183
rect 153212 77846 153332 77874
rect 153108 64796 153160 64802
rect 153108 64738 153160 64744
rect 153016 38140 153068 38146
rect 153016 38082 153068 38088
rect 152832 32632 152884 32638
rect 152832 32574 152884 32580
rect 153212 24410 153240 77846
rect 153292 76832 153344 76838
rect 153292 76774 153344 76780
rect 153304 25770 153332 76774
rect 153396 68105 153424 79630
rect 153474 79591 153530 79600
rect 153488 73545 153516 79591
rect 153474 73536 153530 73545
rect 153474 73471 153530 73480
rect 153580 71194 153608 79784
rect 153936 79756 153988 79762
rect 154086 79744 154114 79897
rect 153936 79698 153988 79704
rect 154040 79716 154114 79744
rect 153660 79688 153712 79694
rect 153658 79656 153660 79665
rect 153712 79656 153714 79665
rect 153842 79656 153898 79665
rect 153658 79591 153714 79600
rect 153752 79620 153804 79626
rect 153842 79591 153898 79600
rect 153752 79562 153804 79568
rect 153660 79552 153712 79558
rect 153660 79494 153712 79500
rect 153568 71188 153620 71194
rect 153568 71130 153620 71136
rect 153580 70394 153608 71130
rect 153488 70366 153608 70394
rect 153382 68096 153438 68105
rect 153382 68031 153438 68040
rect 153488 66842 153516 70366
rect 153672 70009 153700 79494
rect 153764 74390 153792 79562
rect 153856 74458 153884 79591
rect 153948 79393 153976 79698
rect 153934 79384 153990 79393
rect 153934 79319 153990 79328
rect 153936 79280 153988 79286
rect 153936 79222 153988 79228
rect 153948 78470 153976 79222
rect 153936 78464 153988 78470
rect 153936 78406 153988 78412
rect 153844 74452 153896 74458
rect 153844 74394 153896 74400
rect 153752 74384 153804 74390
rect 153752 74326 153804 74332
rect 153856 74254 153884 74394
rect 153844 74248 153896 74254
rect 153844 74190 153896 74196
rect 153948 70394 153976 78406
rect 154040 76838 154068 79716
rect 154178 79608 154206 80036
rect 154270 79812 154298 80036
rect 154362 79966 154390 80036
rect 154454 79971 154482 80036
rect 154350 79960 154402 79966
rect 154350 79902 154402 79908
rect 154440 79962 154496 79971
rect 154440 79897 154496 79906
rect 154546 79812 154574 80036
rect 154270 79801 154344 79812
rect 154270 79792 154358 79801
rect 154270 79784 154302 79792
rect 154302 79727 154358 79736
rect 154500 79784 154574 79812
rect 154132 79580 154206 79608
rect 154394 79656 154450 79665
rect 154394 79591 154450 79600
rect 154132 79286 154160 79580
rect 154304 79552 154356 79558
rect 154210 79520 154266 79529
rect 154304 79494 154356 79500
rect 154210 79455 154266 79464
rect 154120 79280 154172 79286
rect 154120 79222 154172 79228
rect 154224 77294 154252 79455
rect 154132 77266 154252 77294
rect 154028 76832 154080 76838
rect 154028 76774 154080 76780
rect 154132 75585 154160 77266
rect 154316 77217 154344 79494
rect 154302 77208 154358 77217
rect 154302 77143 154358 77152
rect 154118 75576 154174 75585
rect 154118 75511 154174 75520
rect 153856 70366 153976 70394
rect 153658 70000 153714 70009
rect 153658 69935 153714 69944
rect 153476 66836 153528 66842
rect 153476 66778 153528 66784
rect 153292 25764 153344 25770
rect 153292 25706 153344 25712
rect 153200 24404 153252 24410
rect 153200 24346 153252 24352
rect 153856 20194 153884 70366
rect 154026 70000 154082 70009
rect 154026 69935 154082 69944
rect 153934 68096 153990 68105
rect 153934 68031 153990 68040
rect 153844 20188 153896 20194
rect 153844 20130 153896 20136
rect 152740 18828 152792 18834
rect 152740 18770 152792 18776
rect 153948 14754 153976 68031
rect 154040 36718 154068 69935
rect 154132 58818 154160 75511
rect 154316 64874 154344 77143
rect 154408 74361 154436 79591
rect 154500 76401 154528 79784
rect 154638 79744 154666 80036
rect 154730 79830 154758 80036
rect 154822 79966 154850 80036
rect 154810 79960 154862 79966
rect 154810 79902 154862 79908
rect 154914 79898 154942 80036
rect 155006 79971 155034 80036
rect 154992 79962 155048 79971
rect 155098 79966 155126 80036
rect 155190 79966 155218 80036
rect 155282 79971 155310 80036
rect 154902 79892 154954 79898
rect 154992 79897 155048 79906
rect 155086 79960 155138 79966
rect 155086 79902 155138 79908
rect 155178 79960 155230 79966
rect 155178 79902 155230 79908
rect 155268 79962 155324 79971
rect 155268 79897 155324 79906
rect 154718 79824 154770 79830
rect 154718 79766 154770 79772
rect 154808 79826 154864 79835
rect 154902 79834 154954 79840
rect 154808 79761 154864 79770
rect 154592 79716 154666 79744
rect 154948 79756 155000 79762
rect 154486 76392 154542 76401
rect 154486 76327 154542 76336
rect 154592 75546 154620 79716
rect 155374 79744 155402 80036
rect 155466 79966 155494 80036
rect 155454 79960 155506 79966
rect 155558 79937 155586 80036
rect 155650 79966 155678 80036
rect 155638 79960 155690 79966
rect 155454 79902 155506 79908
rect 155544 79928 155600 79937
rect 155638 79902 155690 79908
rect 155742 79898 155770 80036
rect 155834 79898 155862 80036
rect 155926 79971 155954 80036
rect 155912 79962 155968 79971
rect 155544 79863 155600 79872
rect 155730 79892 155782 79898
rect 155730 79834 155782 79840
rect 155822 79892 155874 79898
rect 155912 79897 155968 79906
rect 155822 79834 155874 79840
rect 155500 79824 155552 79830
rect 155500 79766 155552 79772
rect 155592 79824 155644 79830
rect 155592 79766 155644 79772
rect 155374 79716 155448 79744
rect 154948 79698 155000 79704
rect 154672 79620 154724 79626
rect 154672 79562 154724 79568
rect 154764 79620 154816 79626
rect 154764 79562 154816 79568
rect 154580 75540 154632 75546
rect 154580 75482 154632 75488
rect 154684 75392 154712 79562
rect 154592 75364 154712 75392
rect 154488 74384 154540 74390
rect 154394 74352 154450 74361
rect 154488 74326 154540 74332
rect 154394 74287 154450 74296
rect 154396 74248 154448 74254
rect 154396 74190 154448 74196
rect 154408 67114 154436 74190
rect 154500 72758 154528 74326
rect 154488 72752 154540 72758
rect 154488 72694 154540 72700
rect 154396 67108 154448 67114
rect 154396 67050 154448 67056
rect 154500 66994 154528 72694
rect 154224 64846 154344 64874
rect 154408 66966 154528 66994
rect 154224 61538 154252 64846
rect 154212 61532 154264 61538
rect 154212 61474 154264 61480
rect 154120 58812 154172 58818
rect 154120 58754 154172 58760
rect 154028 36712 154080 36718
rect 154028 36654 154080 36660
rect 154408 27130 154436 66966
rect 154488 66836 154540 66842
rect 154488 66778 154540 66784
rect 154396 27124 154448 27130
rect 154396 27066 154448 27072
rect 153936 14748 153988 14754
rect 153936 14690 153988 14696
rect 152648 13388 152700 13394
rect 152648 13330 152700 13336
rect 152556 6588 152608 6594
rect 152556 6530 152608 6536
rect 154500 5030 154528 66778
rect 154592 46918 154620 75364
rect 154672 75064 154724 75070
rect 154672 75006 154724 75012
rect 154684 60722 154712 75006
rect 154776 63442 154804 79562
rect 154854 78160 154910 78169
rect 154854 78095 154910 78104
rect 154868 66201 154896 78095
rect 154960 77314 154988 79698
rect 155132 79484 155184 79490
rect 155132 79426 155184 79432
rect 154948 77308 155000 77314
rect 154948 77250 155000 77256
rect 154948 76492 155000 76498
rect 154948 76434 155000 76440
rect 154854 66192 154910 66201
rect 154854 66127 154910 66136
rect 154868 64874 154896 66127
rect 154960 65958 154988 76434
rect 155144 70394 155172 79426
rect 155420 76498 155448 79716
rect 155512 77246 155540 79766
rect 155500 77240 155552 77246
rect 155500 77182 155552 77188
rect 155408 76492 155460 76498
rect 155408 76434 155460 76440
rect 155500 75540 155552 75546
rect 155500 75482 155552 75488
rect 155512 71505 155540 75482
rect 155604 75070 155632 79766
rect 155776 79756 155828 79762
rect 156018 79744 156046 80036
rect 156110 79971 156138 80036
rect 156096 79962 156152 79971
rect 156202 79966 156230 80036
rect 156294 79971 156322 80036
rect 156096 79897 156152 79906
rect 156190 79960 156242 79966
rect 156190 79902 156242 79908
rect 156280 79962 156336 79971
rect 156386 79966 156414 80036
rect 156280 79897 156336 79906
rect 156374 79960 156426 79966
rect 156374 79902 156426 79908
rect 156478 79898 156506 80036
rect 156466 79892 156518 79898
rect 156466 79834 156518 79840
rect 156570 79744 156598 80036
rect 156662 79898 156690 80036
rect 156754 79971 156782 80036
rect 156740 79962 156796 79971
rect 156846 79966 156874 80036
rect 156650 79892 156702 79898
rect 156740 79897 156796 79906
rect 156834 79960 156886 79966
rect 156834 79902 156886 79908
rect 156938 79898 156966 80036
rect 156650 79834 156702 79840
rect 156926 79892 156978 79898
rect 156926 79834 156978 79840
rect 157030 79744 157058 80036
rect 155776 79698 155828 79704
rect 155880 79716 156046 79744
rect 156524 79716 156598 79744
rect 156984 79716 157058 79744
rect 155682 79656 155738 79665
rect 155682 79591 155738 79600
rect 155592 75064 155644 75070
rect 155592 75006 155644 75012
rect 155696 72282 155724 79591
rect 155788 73154 155816 79698
rect 155880 74254 155908 79716
rect 156236 79688 156288 79694
rect 156236 79630 156288 79636
rect 156418 79656 156474 79665
rect 156052 79552 156104 79558
rect 156052 79494 156104 79500
rect 156144 79552 156196 79558
rect 156144 79494 156196 79500
rect 155960 79484 156012 79490
rect 155960 79426 156012 79432
rect 155972 78033 156000 79426
rect 156064 79257 156092 79494
rect 156050 79248 156106 79257
rect 156050 79183 156106 79192
rect 156052 79076 156104 79082
rect 156052 79018 156104 79024
rect 155958 78024 156014 78033
rect 155958 77959 156014 77968
rect 155960 76492 156012 76498
rect 155960 76434 156012 76440
rect 155868 74248 155920 74254
rect 155868 74190 155920 74196
rect 155788 73126 155908 73154
rect 155880 72690 155908 73126
rect 155868 72684 155920 72690
rect 155868 72626 155920 72632
rect 155684 72276 155736 72282
rect 155684 72218 155736 72224
rect 155498 71496 155554 71505
rect 155498 71431 155554 71440
rect 155052 70366 155172 70394
rect 155052 69018 155080 70366
rect 155040 69012 155092 69018
rect 155040 68954 155092 68960
rect 154948 65952 155000 65958
rect 154948 65894 155000 65900
rect 155512 64874 155540 71431
rect 155880 70394 155908 72626
rect 154868 64846 155264 64874
rect 154764 63436 154816 63442
rect 154764 63378 154816 63384
rect 154672 60716 154724 60722
rect 154672 60658 154724 60664
rect 154580 46912 154632 46918
rect 154580 46854 154632 46860
rect 155236 20058 155264 64846
rect 155328 64846 155540 64874
rect 155788 70366 155908 70394
rect 155328 42294 155356 64846
rect 155316 42288 155368 42294
rect 155316 42230 155368 42236
rect 155788 31346 155816 70366
rect 155868 69012 155920 69018
rect 155868 68954 155920 68960
rect 155776 31340 155828 31346
rect 155776 31282 155828 31288
rect 155880 20126 155908 68954
rect 155868 20120 155920 20126
rect 155868 20062 155920 20068
rect 155224 20052 155276 20058
rect 155224 19994 155276 20000
rect 154580 19984 154632 19990
rect 154580 19926 154632 19932
rect 154592 16574 154620 19926
rect 154592 16546 155448 16574
rect 154488 5024 154540 5030
rect 154488 4966 154540 4972
rect 153016 4140 153068 4146
rect 153016 4082 153068 4088
rect 152464 3936 152516 3942
rect 152464 3878 152516 3884
rect 149612 3868 149664 3874
rect 149612 3810 149664 3816
rect 149796 3868 149848 3874
rect 149796 3810 149848 3816
rect 149624 3670 149652 3810
rect 150624 3800 150676 3806
rect 150624 3742 150676 3748
rect 149520 3664 149572 3670
rect 149520 3606 149572 3612
rect 149612 3664 149664 3670
rect 149612 3606 149664 3612
rect 148416 3052 148468 3058
rect 148416 2994 148468 3000
rect 149532 480 149560 3606
rect 150636 480 150664 3742
rect 151820 3392 151872 3398
rect 151820 3334 151872 3340
rect 151832 480 151860 3334
rect 153028 480 153056 4082
rect 154212 3052 154264 3058
rect 154212 2994 154264 3000
rect 154224 480 154252 2994
rect 155420 480 155448 16546
rect 155972 14686 156000 76434
rect 156064 75426 156092 79018
rect 156156 75546 156184 79494
rect 156248 78305 156276 79630
rect 156418 79591 156474 79600
rect 156326 79520 156382 79529
rect 156326 79455 156382 79464
rect 156234 78296 156290 78305
rect 156234 78231 156290 78240
rect 156236 78192 156288 78198
rect 156236 78134 156288 78140
rect 156144 75540 156196 75546
rect 156144 75482 156196 75488
rect 156064 75398 156184 75426
rect 156052 75200 156104 75206
rect 156052 75142 156104 75148
rect 156064 55214 156092 75142
rect 156156 62014 156184 75398
rect 156248 74390 156276 78134
rect 156340 74866 156368 79455
rect 156328 74860 156380 74866
rect 156328 74802 156380 74808
rect 156236 74384 156288 74390
rect 156236 74326 156288 74332
rect 156432 72554 156460 79591
rect 156524 77994 156552 79716
rect 156694 79656 156750 79665
rect 156604 79620 156656 79626
rect 156878 79656 156934 79665
rect 156694 79591 156750 79600
rect 156788 79620 156840 79626
rect 156604 79562 156656 79568
rect 156512 77988 156564 77994
rect 156512 77930 156564 77936
rect 156616 75313 156644 79562
rect 156708 79082 156736 79591
rect 156878 79591 156934 79600
rect 156788 79562 156840 79568
rect 156696 79076 156748 79082
rect 156696 79018 156748 79024
rect 156800 78928 156828 79562
rect 156708 78900 156828 78928
rect 156602 75304 156658 75313
rect 156602 75239 156658 75248
rect 156708 73030 156736 78900
rect 156892 78792 156920 79591
rect 156800 78764 156920 78792
rect 156800 75721 156828 78764
rect 156880 77988 156932 77994
rect 156880 77930 156932 77936
rect 156786 75712 156842 75721
rect 156786 75647 156842 75656
rect 156788 75540 156840 75546
rect 156788 75482 156840 75488
rect 156800 74186 156828 75482
rect 156892 74338 156920 77930
rect 156984 75206 157012 79716
rect 157122 79642 157150 80036
rect 157214 79830 157242 80036
rect 157306 79937 157334 80036
rect 157398 79966 157426 80036
rect 157490 79971 157518 80036
rect 157386 79960 157438 79966
rect 157292 79928 157348 79937
rect 157386 79902 157438 79908
rect 157476 79962 157532 79971
rect 157476 79897 157532 79906
rect 157292 79863 157348 79872
rect 157202 79824 157254 79830
rect 157582 79778 157610 80036
rect 157674 79966 157702 80036
rect 157662 79960 157714 79966
rect 157662 79902 157714 79908
rect 157766 79898 157794 80036
rect 157754 79892 157806 79898
rect 157754 79834 157806 79840
rect 157202 79766 157254 79772
rect 157536 79750 157610 79778
rect 157858 79778 157886 80036
rect 157950 79966 157978 80036
rect 158042 79966 158070 80036
rect 157938 79960 157990 79966
rect 157938 79902 157990 79908
rect 158030 79960 158082 79966
rect 158134 79937 158162 80036
rect 158226 79966 158254 80036
rect 158214 79960 158266 79966
rect 158030 79902 158082 79908
rect 158120 79928 158176 79937
rect 158214 79902 158266 79908
rect 158120 79863 158176 79872
rect 158168 79824 158220 79830
rect 157708 79756 157760 79762
rect 157248 79688 157300 79694
rect 157122 79614 157196 79642
rect 157248 79630 157300 79636
rect 157340 79688 157392 79694
rect 157340 79630 157392 79636
rect 157064 79484 157116 79490
rect 157064 79426 157116 79432
rect 157076 76498 157104 79426
rect 157168 78742 157196 79614
rect 157156 78736 157208 78742
rect 157156 78678 157208 78684
rect 157064 76492 157116 76498
rect 157064 76434 157116 76440
rect 156972 75200 157024 75206
rect 156972 75142 157024 75148
rect 156892 74310 157104 74338
rect 156972 74248 157024 74254
rect 156972 74190 157024 74196
rect 156788 74180 156840 74186
rect 156788 74122 156840 74128
rect 156696 73024 156748 73030
rect 156696 72966 156748 72972
rect 156420 72548 156472 72554
rect 156420 72490 156472 72496
rect 156800 70394 156828 74122
rect 156800 70366 156920 70394
rect 156892 64874 156920 70366
rect 156708 64846 156920 64874
rect 156144 62008 156196 62014
rect 156144 61950 156196 61956
rect 156052 55208 156104 55214
rect 156052 55150 156104 55156
rect 156708 41002 156736 64846
rect 156696 40996 156748 41002
rect 156696 40938 156748 40944
rect 156050 35184 156106 35193
rect 156050 35119 156106 35128
rect 156064 16574 156092 35119
rect 156984 29918 157012 74190
rect 157076 70922 157104 74310
rect 157156 73024 157208 73030
rect 157156 72966 157208 72972
rect 157168 72842 157196 72966
rect 157260 72962 157288 79630
rect 157248 72956 157300 72962
rect 157248 72898 157300 72904
rect 157168 72814 157288 72842
rect 157156 72548 157208 72554
rect 157156 72490 157208 72496
rect 157064 70916 157116 70922
rect 157064 70858 157116 70864
rect 156972 29912 157024 29918
rect 156972 29854 157024 29860
rect 157076 22982 157104 70858
rect 157064 22976 157116 22982
rect 157064 22918 157116 22924
rect 156064 16546 156184 16574
rect 155960 14680 156012 14686
rect 155960 14622 156012 14628
rect 148294 354 148406 480
rect 147876 326 148406 354
rect 148294 -960 148406 326
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156156 354 156184 16546
rect 157168 13326 157196 72490
rect 157156 13320 157208 13326
rect 157156 13262 157208 13268
rect 157260 9110 157288 72814
rect 157352 71534 157380 79630
rect 157432 78668 157484 78674
rect 157432 78610 157484 78616
rect 157340 71528 157392 71534
rect 157340 71470 157392 71476
rect 157340 71392 157392 71398
rect 157340 71334 157392 71340
rect 157352 18766 157380 71334
rect 157444 59294 157472 78610
rect 157536 77586 157564 79750
rect 157858 79750 157932 79778
rect 158318 79812 158346 80036
rect 158410 79966 158438 80036
rect 158502 79966 158530 80036
rect 158594 79971 158622 80036
rect 158398 79960 158450 79966
rect 158398 79902 158450 79908
rect 158490 79960 158542 79966
rect 158490 79902 158542 79908
rect 158580 79962 158636 79971
rect 158580 79897 158636 79906
rect 158220 79784 158346 79812
rect 158536 79824 158588 79830
rect 158168 79766 158220 79772
rect 158536 79766 158588 79772
rect 157708 79698 157760 79704
rect 157616 79688 157668 79694
rect 157616 79630 157668 79636
rect 157524 77580 157576 77586
rect 157524 77522 157576 77528
rect 157628 73154 157656 79630
rect 157536 73126 157656 73154
rect 157536 71670 157564 73126
rect 157720 72894 157748 79698
rect 157800 79552 157852 79558
rect 157800 79494 157852 79500
rect 157812 79257 157840 79494
rect 157798 79248 157854 79257
rect 157798 79183 157854 79192
rect 157800 79144 157852 79150
rect 157800 79086 157852 79092
rect 157708 72888 157760 72894
rect 157708 72830 157760 72836
rect 157524 71664 157576 71670
rect 157524 71606 157576 71612
rect 157812 71398 157840 79086
rect 157904 78674 157932 79750
rect 157984 79756 158036 79762
rect 157984 79698 158036 79704
rect 158076 79756 158128 79762
rect 158076 79698 158128 79704
rect 157892 78668 157944 78674
rect 157892 78610 157944 78616
rect 157996 73778 158024 79698
rect 158088 79150 158116 79698
rect 158168 79688 158220 79694
rect 158168 79630 158220 79636
rect 158260 79688 158312 79694
rect 158260 79630 158312 79636
rect 158442 79656 158498 79665
rect 158076 79144 158128 79150
rect 158076 79086 158128 79092
rect 158180 78674 158208 79630
rect 158168 78668 158220 78674
rect 158168 78610 158220 78616
rect 157984 73772 158036 73778
rect 157984 73714 158036 73720
rect 158272 72826 158300 79630
rect 158442 79591 158498 79600
rect 158548 79608 158576 79766
rect 158686 79676 158714 80036
rect 158778 79830 158806 80036
rect 158870 79898 158898 80036
rect 158962 79898 158990 80036
rect 158858 79892 158910 79898
rect 158858 79834 158910 79840
rect 158950 79892 159002 79898
rect 158950 79834 159002 79840
rect 158766 79824 158818 79830
rect 158766 79766 158818 79772
rect 158902 79792 158958 79801
rect 159054 79778 159082 80036
rect 158958 79750 159082 79778
rect 159146 79778 159174 80036
rect 159238 79966 159266 80036
rect 159330 79971 159358 80036
rect 159226 79960 159278 79966
rect 159226 79902 159278 79908
rect 159316 79962 159372 79971
rect 159316 79897 159372 79906
rect 159422 79830 159450 80036
rect 159514 79937 159542 80036
rect 159500 79928 159556 79937
rect 159500 79863 159556 79872
rect 159410 79824 159462 79830
rect 159146 79750 159220 79778
rect 159606 79812 159634 80036
rect 159698 79898 159726 80036
rect 159686 79892 159738 79898
rect 159686 79834 159738 79840
rect 159410 79766 159462 79772
rect 159560 79784 159634 79812
rect 159790 79801 159818 80036
rect 159882 79966 159910 80036
rect 159870 79960 159922 79966
rect 159974 79937 160002 80036
rect 159870 79902 159922 79908
rect 159960 79928 160016 79937
rect 159960 79863 160016 79872
rect 159776 79792 159832 79801
rect 158902 79727 158958 79736
rect 158686 79648 158944 79676
rect 158352 79484 158404 79490
rect 158352 79426 158404 79432
rect 158364 79354 158392 79426
rect 158352 79348 158404 79354
rect 158352 79290 158404 79296
rect 158352 78668 158404 78674
rect 158352 78610 158404 78616
rect 158260 72820 158312 72826
rect 158260 72762 158312 72768
rect 158272 72434 158300 72762
rect 158364 72622 158392 78610
rect 158456 78062 158484 79591
rect 158548 79580 158668 79608
rect 158536 79484 158588 79490
rect 158536 79426 158588 79432
rect 158444 78056 158496 78062
rect 158444 77998 158496 78004
rect 158548 73982 158576 79426
rect 158640 75614 158668 79580
rect 158810 79520 158866 79529
rect 158720 79484 158772 79490
rect 158810 79455 158866 79464
rect 158720 79426 158772 79432
rect 158732 76498 158760 79426
rect 158720 76492 158772 76498
rect 158720 76434 158772 76440
rect 158628 75608 158680 75614
rect 158628 75550 158680 75556
rect 158536 73976 158588 73982
rect 158536 73918 158588 73924
rect 158536 73772 158588 73778
rect 158536 73714 158588 73720
rect 158352 72616 158404 72622
rect 158352 72558 158404 72564
rect 158272 72406 158392 72434
rect 158260 71664 158312 71670
rect 158260 71606 158312 71612
rect 157800 71392 157852 71398
rect 157800 71334 157852 71340
rect 157432 59288 157484 59294
rect 157432 59230 157484 59236
rect 157432 51740 157484 51746
rect 157432 51682 157484 51688
rect 157340 18760 157392 18766
rect 157340 18702 157392 18708
rect 157444 16574 157472 51682
rect 158272 39574 158300 71606
rect 158364 40934 158392 72406
rect 158444 71528 158496 71534
rect 158444 71470 158496 71476
rect 158456 71398 158484 71470
rect 158444 71392 158496 71398
rect 158444 71334 158496 71340
rect 158352 40928 158404 40934
rect 158352 40870 158404 40876
rect 158260 39568 158312 39574
rect 158260 39510 158312 39516
rect 158456 35426 158484 71334
rect 158548 70854 158576 73714
rect 158536 70848 158588 70854
rect 158536 70790 158588 70796
rect 158444 35420 158496 35426
rect 158444 35362 158496 35368
rect 157444 16546 157840 16574
rect 157248 9104 157300 9110
rect 157248 9046 157300 9052
rect 157812 480 157840 16546
rect 158548 11966 158576 70790
rect 158536 11960 158588 11966
rect 158536 11902 158588 11908
rect 158640 10538 158668 75550
rect 158720 75132 158772 75138
rect 158720 75074 158772 75080
rect 158732 52426 158760 75074
rect 158824 57934 158852 79455
rect 158916 78713 158944 79648
rect 158996 79620 159048 79626
rect 158996 79562 159048 79568
rect 159088 79620 159140 79626
rect 159088 79562 159140 79568
rect 159008 79082 159036 79562
rect 158996 79076 159048 79082
rect 158996 79018 159048 79024
rect 158902 78704 158958 78713
rect 158902 78639 158958 78648
rect 159100 77294 159128 79562
rect 159008 77266 159128 77294
rect 158904 75064 158956 75070
rect 158904 75006 158956 75012
rect 158916 60654 158944 75006
rect 159008 64598 159036 77266
rect 159088 76492 159140 76498
rect 159088 76434 159140 76440
rect 159100 73098 159128 76434
rect 159088 73092 159140 73098
rect 159088 73034 159140 73040
rect 159192 72350 159220 79750
rect 159270 79656 159326 79665
rect 159560 79642 159588 79784
rect 159776 79727 159832 79736
rect 159914 79792 159970 79801
rect 160066 79778 160094 80036
rect 159914 79727 159970 79736
rect 160020 79750 160094 79778
rect 159270 79591 159326 79600
rect 159376 79614 159588 79642
rect 159284 78674 159312 79591
rect 159272 78668 159324 78674
rect 159272 78610 159324 78616
rect 159376 73846 159404 79614
rect 159456 79552 159508 79558
rect 159456 79494 159508 79500
rect 159468 78849 159496 79494
rect 159640 79484 159692 79490
rect 159640 79426 159692 79432
rect 159824 79484 159876 79490
rect 159824 79426 159876 79432
rect 159454 78840 159510 78849
rect 159454 78775 159510 78784
rect 159546 78704 159602 78713
rect 159456 78668 159508 78674
rect 159546 78639 159602 78648
rect 159456 78610 159508 78616
rect 159468 74254 159496 78610
rect 159560 75313 159588 78639
rect 159546 75304 159602 75313
rect 159546 75239 159602 75248
rect 159652 74458 159680 79426
rect 159730 79248 159786 79257
rect 159730 79183 159786 79192
rect 159640 74452 159692 74458
rect 159640 74394 159692 74400
rect 159456 74248 159508 74254
rect 159456 74190 159508 74196
rect 159364 73840 159416 73846
rect 159364 73782 159416 73788
rect 159180 72344 159232 72350
rect 159180 72286 159232 72292
rect 159468 70394 159496 74190
rect 159744 74050 159772 79183
rect 159836 76702 159864 79426
rect 159824 76696 159876 76702
rect 159824 76638 159876 76644
rect 159928 75070 159956 79727
rect 160020 75138 160048 79750
rect 160158 79744 160186 80036
rect 160250 79812 160278 80036
rect 160342 79937 160370 80036
rect 160434 79966 160462 80036
rect 160526 79966 160554 80036
rect 160618 79966 160646 80036
rect 160422 79960 160474 79966
rect 160328 79928 160384 79937
rect 160422 79902 160474 79908
rect 160514 79960 160566 79966
rect 160514 79902 160566 79908
rect 160606 79960 160658 79966
rect 160606 79902 160658 79908
rect 160710 79898 160738 80036
rect 160328 79863 160384 79872
rect 160698 79892 160750 79898
rect 160698 79834 160750 79840
rect 160376 79824 160428 79830
rect 160250 79784 160324 79812
rect 160158 79716 160232 79744
rect 160100 79620 160152 79626
rect 160100 79562 160152 79568
rect 160008 75132 160060 75138
rect 160008 75074 160060 75080
rect 159916 75064 159968 75070
rect 159916 75006 159968 75012
rect 159732 74044 159784 74050
rect 159732 73986 159784 73992
rect 159916 74044 159968 74050
rect 159916 73986 159968 73992
rect 159824 73976 159876 73982
rect 159824 73918 159876 73924
rect 159836 71466 159864 73918
rect 159928 71670 159956 73986
rect 160008 73840 160060 73846
rect 160008 73782 160060 73788
rect 159916 71664 159968 71670
rect 159916 71606 159968 71612
rect 159824 71460 159876 71466
rect 159824 71402 159876 71408
rect 159468 70366 159772 70394
rect 158996 64592 159048 64598
rect 158996 64534 159048 64540
rect 158904 60648 158956 60654
rect 158904 60590 158956 60596
rect 158812 57928 158864 57934
rect 158812 57870 158864 57876
rect 158720 52420 158772 52426
rect 158720 52362 158772 52368
rect 159744 32570 159772 70366
rect 159732 32564 159784 32570
rect 159732 32506 159784 32512
rect 159836 28490 159864 71402
rect 159824 28484 159876 28490
rect 159824 28426 159876 28432
rect 158628 10532 158680 10538
rect 158628 10474 158680 10480
rect 159928 7818 159956 71606
rect 160020 70990 160048 73782
rect 160008 70984 160060 70990
rect 160008 70926 160060 70932
rect 159916 7812 159968 7818
rect 159916 7754 159968 7760
rect 160020 6526 160048 70926
rect 160112 68921 160140 79562
rect 160204 76906 160232 79716
rect 160192 76900 160244 76906
rect 160192 76842 160244 76848
rect 160192 76696 160244 76702
rect 160192 76638 160244 76644
rect 160098 68912 160154 68921
rect 160098 68847 160154 68856
rect 160204 68542 160232 76638
rect 160192 68536 160244 68542
rect 160192 68478 160244 68484
rect 160296 68338 160324 79784
rect 160428 79801 160508 79812
rect 160428 79792 160522 79801
rect 160428 79784 160466 79792
rect 160376 79766 160428 79772
rect 160466 79727 160522 79736
rect 160802 79744 160830 80036
rect 160894 79937 160922 80036
rect 160880 79928 160936 79937
rect 160880 79863 160936 79872
rect 160986 79744 161014 80036
rect 161078 79898 161106 80036
rect 161170 79966 161198 80036
rect 161158 79960 161210 79966
rect 161158 79902 161210 79908
rect 161262 79898 161290 80036
rect 161354 79898 161382 80036
rect 161066 79892 161118 79898
rect 161066 79834 161118 79840
rect 161250 79892 161302 79898
rect 161250 79834 161302 79840
rect 161342 79892 161394 79898
rect 161342 79834 161394 79840
rect 161446 79801 161474 80036
rect 161538 79966 161566 80036
rect 161630 79966 161658 80036
rect 161722 79966 161750 80036
rect 161814 79971 161842 80036
rect 161526 79960 161578 79966
rect 161526 79902 161578 79908
rect 161618 79960 161670 79966
rect 161618 79902 161670 79908
rect 161710 79960 161762 79966
rect 161710 79902 161762 79908
rect 161800 79962 161856 79971
rect 161800 79897 161856 79906
rect 161906 79898 161934 80036
rect 161998 79898 162026 80036
rect 161894 79892 161946 79898
rect 161894 79834 161946 79840
rect 161986 79892 162038 79898
rect 161986 79834 162038 79840
rect 161432 79792 161488 79801
rect 160802 79716 160876 79744
rect 160986 79716 161060 79744
rect 161664 79756 161716 79762
rect 161432 79727 161488 79736
rect 160374 79656 160430 79665
rect 160374 79591 160430 79600
rect 160388 76702 160416 79591
rect 160560 79552 160612 79558
rect 160560 79494 160612 79500
rect 160468 79484 160520 79490
rect 160468 79426 160520 79432
rect 160376 76696 160428 76702
rect 160376 76638 160428 76644
rect 160480 73154 160508 79426
rect 160388 73126 160508 73154
rect 160388 69834 160416 73126
rect 160572 70394 160600 79494
rect 160744 78736 160796 78742
rect 160744 78678 160796 78684
rect 160756 78266 160784 78678
rect 160744 78260 160796 78266
rect 160744 78202 160796 78208
rect 160744 76900 160796 76906
rect 160744 76842 160796 76848
rect 160756 71534 160784 76842
rect 160848 76702 160876 79716
rect 160928 79484 160980 79490
rect 160928 79426 160980 79432
rect 160836 76696 160888 76702
rect 160836 76638 160888 76644
rect 160744 71528 160796 71534
rect 160744 71470 160796 71476
rect 160480 70366 160600 70394
rect 160756 70394 160784 71470
rect 160940 71262 160968 79426
rect 161032 76362 161060 79716
rect 161584 79716 161664 79744
rect 161112 79688 161164 79694
rect 161388 79688 161440 79694
rect 161112 79630 161164 79636
rect 161308 79648 161388 79676
rect 161020 76356 161072 76362
rect 161020 76298 161072 76304
rect 161124 73166 161152 79630
rect 161204 79552 161256 79558
rect 161204 79494 161256 79500
rect 161216 76809 161244 79494
rect 161308 76945 161336 79648
rect 161388 79630 161440 79636
rect 161480 79620 161532 79626
rect 161480 79562 161532 79568
rect 161492 78690 161520 79562
rect 161400 78662 161520 78690
rect 161294 76936 161350 76945
rect 161294 76871 161350 76880
rect 161202 76800 161258 76809
rect 161202 76735 161258 76744
rect 161296 76696 161348 76702
rect 161296 76638 161348 76644
rect 161112 73160 161164 73166
rect 161112 73102 161164 73108
rect 161112 71732 161164 71738
rect 161112 71674 161164 71680
rect 161124 71398 161152 71674
rect 161112 71392 161164 71398
rect 161308 71369 161336 76638
rect 161400 72418 161428 78662
rect 161480 78600 161532 78606
rect 161480 78542 161532 78548
rect 161388 72412 161440 72418
rect 161388 72354 161440 72360
rect 161112 71334 161164 71340
rect 161294 71360 161350 71369
rect 161294 71295 161350 71304
rect 160928 71256 160980 71262
rect 160928 71198 160980 71204
rect 160756 70366 160876 70394
rect 160480 70106 160508 70366
rect 160468 70100 160520 70106
rect 160468 70042 160520 70048
rect 160376 69828 160428 69834
rect 160376 69770 160428 69776
rect 160284 68332 160336 68338
rect 160284 68274 160336 68280
rect 160848 33998 160876 70366
rect 160836 33992 160888 33998
rect 160836 33934 160888 33940
rect 160100 33788 160152 33794
rect 160100 33730 160152 33736
rect 160008 6520 160060 6526
rect 160008 6462 160060 6468
rect 158902 6216 158958 6225
rect 158902 6151 158958 6160
rect 158916 480 158944 6151
rect 160112 3806 160140 33730
rect 160940 31278 160968 71198
rect 161204 70100 161256 70106
rect 161204 70042 161256 70048
rect 161018 68912 161074 68921
rect 161018 68847 161074 68856
rect 160928 31272 160980 31278
rect 160928 31214 160980 31220
rect 161032 28422 161060 68847
rect 161112 68332 161164 68338
rect 161112 68274 161164 68280
rect 161020 28416 161072 28422
rect 161020 28358 161072 28364
rect 161124 19990 161152 68274
rect 161112 19984 161164 19990
rect 161112 19926 161164 19932
rect 161216 16046 161244 70042
rect 161204 16040 161256 16046
rect 161204 15982 161256 15988
rect 160190 8936 160246 8945
rect 160190 8871 160246 8880
rect 160100 3800 160152 3806
rect 160100 3742 160152 3748
rect 160204 3482 160232 8871
rect 161308 7750 161336 71295
rect 161296 7744 161348 7750
rect 161296 7686 161348 7692
rect 161400 4962 161428 72354
rect 161492 59362 161520 78542
rect 161584 76906 161612 79716
rect 161664 79698 161716 79704
rect 161848 79756 161900 79762
rect 162090 79744 162118 80036
rect 161900 79716 161980 79744
rect 161848 79698 161900 79704
rect 161846 79656 161902 79665
rect 161664 79620 161716 79626
rect 161846 79591 161902 79600
rect 161664 79562 161716 79568
rect 161676 78606 161704 79562
rect 161756 79552 161808 79558
rect 161756 79494 161808 79500
rect 161664 78600 161716 78606
rect 161664 78542 161716 78548
rect 161664 78464 161716 78470
rect 161664 78406 161716 78412
rect 161572 76900 161624 76906
rect 161572 76842 161624 76848
rect 161572 76696 161624 76702
rect 161572 76638 161624 76644
rect 161584 65754 161612 76638
rect 161676 66094 161704 78406
rect 161768 77294 161796 79494
rect 161860 77518 161888 79591
rect 161848 77512 161900 77518
rect 161848 77454 161900 77460
rect 161768 77266 161888 77294
rect 161756 74792 161808 74798
rect 161756 74734 161808 74740
rect 161768 66230 161796 74734
rect 161860 70242 161888 77266
rect 161952 76702 161980 79716
rect 162044 79716 162118 79744
rect 161940 76696 161992 76702
rect 161940 76638 161992 76644
rect 162044 70394 162072 79716
rect 162182 79676 162210 80036
rect 162274 79744 162302 80036
rect 162366 79812 162394 80036
rect 162458 79966 162486 80036
rect 162446 79960 162498 79966
rect 162446 79902 162498 79908
rect 162366 79784 162440 79812
rect 162550 79801 162578 80036
rect 162274 79716 162348 79744
rect 162182 79648 162256 79676
rect 162124 79416 162176 79422
rect 162122 79384 162124 79393
rect 162176 79384 162178 79393
rect 162122 79319 162178 79328
rect 162124 79144 162176 79150
rect 162122 79112 162124 79121
rect 162176 79112 162178 79121
rect 162122 79047 162178 79056
rect 162228 78690 162256 79648
rect 162136 78662 162256 78690
rect 162136 73642 162164 78662
rect 162216 78056 162268 78062
rect 162216 77998 162268 78004
rect 162228 73846 162256 77998
rect 162320 76809 162348 79716
rect 162412 77790 162440 79784
rect 162536 79792 162592 79801
rect 162536 79727 162592 79736
rect 162492 79688 162544 79694
rect 162642 79676 162670 80036
rect 162734 79744 162762 80036
rect 162826 79937 162854 80036
rect 162812 79928 162868 79937
rect 162812 79863 162868 79872
rect 162918 79801 162946 80036
rect 163010 79812 163038 80036
rect 163102 79937 163130 80036
rect 163088 79928 163144 79937
rect 163194 79898 163222 80036
rect 163286 79898 163314 80036
rect 163378 79966 163406 80036
rect 163366 79960 163418 79966
rect 163366 79902 163418 79908
rect 163088 79863 163144 79872
rect 163182 79892 163234 79898
rect 163182 79834 163234 79840
rect 163274 79892 163326 79898
rect 163274 79834 163326 79840
rect 162904 79792 162960 79801
rect 162734 79716 162808 79744
rect 163010 79784 163084 79812
rect 163056 79778 163084 79784
rect 163056 79750 163130 79778
rect 162904 79727 162960 79736
rect 162492 79630 162544 79636
rect 162596 79648 162670 79676
rect 162504 78470 162532 79630
rect 162492 78464 162544 78470
rect 162492 78406 162544 78412
rect 162492 78260 162544 78266
rect 162492 78202 162544 78208
rect 162400 77784 162452 77790
rect 162400 77726 162452 77732
rect 162400 77512 162452 77518
rect 162400 77454 162452 77460
rect 162306 76800 162362 76809
rect 162306 76735 162362 76744
rect 162216 73840 162268 73846
rect 162216 73782 162268 73788
rect 162124 73636 162176 73642
rect 162124 73578 162176 73584
rect 162412 73154 162440 77454
rect 161952 70366 162072 70394
rect 162320 73126 162440 73154
rect 162504 73154 162532 78202
rect 162596 77217 162624 79648
rect 162676 79552 162728 79558
rect 162676 79494 162728 79500
rect 162688 79014 162716 79494
rect 162676 79008 162728 79014
rect 162676 78950 162728 78956
rect 162780 77874 162808 79716
rect 162950 79656 163006 79665
rect 162860 79620 162912 79626
rect 163102 79642 163130 79750
rect 163470 79744 163498 80036
rect 163562 79830 163590 80036
rect 163550 79824 163602 79830
rect 163550 79766 163602 79772
rect 163332 79716 163498 79744
rect 163102 79614 163176 79642
rect 162950 79591 163006 79600
rect 162860 79562 162912 79568
rect 162872 79354 162900 79562
rect 162860 79348 162912 79354
rect 162860 79290 162912 79296
rect 162688 77846 162808 77874
rect 162582 77208 162638 77217
rect 162582 77143 162638 77152
rect 162688 74798 162716 77846
rect 162768 77784 162820 77790
rect 162768 77726 162820 77732
rect 162676 74792 162728 74798
rect 162676 74734 162728 74740
rect 162504 73126 162624 73154
rect 161848 70236 161900 70242
rect 161848 70178 161900 70184
rect 161756 66224 161808 66230
rect 161756 66166 161808 66172
rect 161664 66088 161716 66094
rect 161664 66030 161716 66036
rect 161860 66042 161888 70178
rect 161952 69630 161980 70366
rect 162320 70174 162348 73126
rect 162596 70394 162624 73126
rect 162780 71398 162808 77726
rect 162860 76764 162912 76770
rect 162860 76706 162912 76712
rect 162768 71392 162820 71398
rect 162768 71334 162820 71340
rect 162504 70366 162624 70394
rect 162308 70168 162360 70174
rect 162308 70110 162360 70116
rect 161940 69624 161992 69630
rect 161940 69566 161992 69572
rect 162320 66722 162348 70110
rect 162504 67046 162532 70366
rect 162676 69624 162728 69630
rect 162676 69566 162728 69572
rect 162492 67040 162544 67046
rect 162492 66982 162544 66988
rect 162320 66694 162440 66722
rect 161860 66014 162348 66042
rect 161572 65748 161624 65754
rect 161572 65690 161624 65696
rect 162124 65748 162176 65754
rect 162124 65690 162176 65696
rect 161480 59356 161532 59362
rect 161480 59298 161532 59304
rect 162136 33930 162164 65690
rect 162124 33924 162176 33930
rect 162124 33866 162176 33872
rect 162320 27062 162348 66014
rect 162308 27056 162360 27062
rect 162308 26998 162360 27004
rect 162412 25702 162440 66694
rect 162492 66224 162544 66230
rect 162492 66166 162544 66172
rect 162400 25696 162452 25702
rect 162400 25638 162452 25644
rect 162504 13190 162532 66166
rect 162584 66088 162636 66094
rect 162584 66030 162636 66036
rect 162596 65890 162624 66030
rect 162584 65884 162636 65890
rect 162584 65826 162636 65832
rect 162492 13184 162544 13190
rect 162492 13126 162544 13132
rect 162596 10470 162624 65826
rect 162688 13258 162716 69566
rect 162780 14618 162808 71334
rect 162872 52358 162900 76706
rect 162964 53786 162992 79591
rect 163044 79552 163096 79558
rect 163044 79494 163096 79500
rect 163056 61946 163084 79494
rect 163148 78402 163176 79614
rect 163228 79552 163280 79558
rect 163228 79494 163280 79500
rect 163136 78396 163188 78402
rect 163136 78338 163188 78344
rect 163240 76702 163268 79494
rect 163228 76696 163280 76702
rect 163228 76638 163280 76644
rect 163228 76492 163280 76498
rect 163228 76434 163280 76440
rect 163136 74112 163188 74118
rect 163136 74054 163188 74060
rect 163148 64569 163176 74054
rect 163240 68950 163268 76434
rect 163332 69970 163360 79716
rect 163654 79676 163682 80036
rect 163746 79744 163774 80036
rect 163838 79812 163866 80036
rect 163930 79937 163958 80036
rect 163916 79928 163972 79937
rect 163916 79863 163972 79872
rect 163838 79784 163912 79812
rect 163746 79716 163820 79744
rect 163654 79648 163728 79676
rect 163504 79620 163556 79626
rect 163504 79562 163556 79568
rect 163412 76696 163464 76702
rect 163412 76638 163464 76644
rect 163320 69964 163372 69970
rect 163320 69906 163372 69912
rect 163424 69766 163452 76638
rect 163516 73982 163544 79562
rect 163700 76770 163728 79648
rect 163688 76764 163740 76770
rect 163688 76706 163740 76712
rect 163792 76430 163820 79716
rect 163780 76424 163832 76430
rect 163780 76366 163832 76372
rect 163884 74118 163912 79784
rect 164022 79744 164050 80036
rect 163976 79716 164050 79744
rect 164114 79744 164142 80036
rect 164206 79903 164234 80036
rect 164298 79966 164326 80036
rect 164286 79960 164338 79966
rect 164192 79894 164248 79903
rect 164286 79902 164338 79908
rect 164192 79829 164248 79838
rect 164286 79824 164338 79830
rect 164286 79766 164338 79772
rect 164114 79716 164188 79744
rect 163976 76498 164004 79716
rect 164056 79620 164108 79626
rect 164056 79562 164108 79568
rect 164068 78062 164096 79562
rect 164160 78198 164188 79716
rect 164298 79642 164326 79766
rect 164390 79744 164418 80036
rect 164482 79812 164510 80036
rect 164574 79937 164602 80036
rect 164666 79966 164694 80036
rect 164654 79960 164706 79966
rect 164560 79928 164616 79937
rect 164758 79937 164786 80036
rect 164850 79966 164878 80036
rect 164838 79960 164890 79966
rect 164654 79902 164706 79908
rect 164744 79928 164800 79937
rect 164560 79863 164616 79872
rect 164838 79902 164890 79908
rect 164744 79863 164800 79872
rect 164482 79784 164556 79812
rect 164390 79716 164464 79744
rect 164298 79614 164372 79642
rect 164240 79552 164292 79558
rect 164240 79494 164292 79500
rect 164252 78266 164280 79494
rect 164240 78260 164292 78266
rect 164240 78202 164292 78208
rect 164148 78192 164200 78198
rect 164148 78134 164200 78140
rect 164240 78124 164292 78130
rect 164240 78066 164292 78072
rect 164056 78056 164108 78062
rect 164056 77998 164108 78004
rect 164148 76900 164200 76906
rect 164148 76842 164200 76848
rect 163964 76492 164016 76498
rect 163964 76434 164016 76440
rect 163872 74112 163924 74118
rect 163872 74054 163924 74060
rect 164160 74050 164188 76842
rect 164148 74044 164200 74050
rect 164148 73986 164200 73992
rect 163504 73976 163556 73982
rect 163504 73918 163556 73924
rect 164056 70304 164108 70310
rect 164056 70246 164108 70252
rect 163964 70032 164016 70038
rect 163964 69974 164016 69980
rect 163976 69766 164004 69974
rect 164068 69970 164096 70246
rect 164056 69964 164108 69970
rect 164056 69906 164108 69912
rect 163412 69760 163464 69766
rect 163412 69702 163464 69708
rect 163964 69760 164016 69766
rect 163964 69702 164016 69708
rect 163228 68944 163280 68950
rect 163228 68886 163280 68892
rect 163872 68944 163924 68950
rect 163872 68886 163924 68892
rect 163884 68610 163912 68886
rect 163872 68604 163924 68610
rect 163872 68546 163924 68552
rect 163134 64560 163190 64569
rect 163134 64495 163190 64504
rect 163148 63617 163176 64495
rect 163134 63608 163190 63617
rect 163134 63543 163190 63552
rect 163778 63608 163834 63617
rect 163778 63543 163834 63552
rect 163044 61940 163096 61946
rect 163044 61882 163096 61888
rect 162952 53780 163004 53786
rect 162952 53722 163004 53728
rect 163504 53100 163556 53106
rect 163504 53042 163556 53048
rect 162860 52352 162912 52358
rect 162860 52294 162912 52300
rect 162768 14612 162820 14618
rect 162768 14554 162820 14560
rect 162676 13252 162728 13258
rect 162676 13194 162728 13200
rect 162584 10464 162636 10470
rect 162584 10406 162636 10412
rect 161388 4956 161440 4962
rect 161388 4898 161440 4904
rect 161388 3936 161440 3942
rect 161388 3878 161440 3884
rect 161400 3806 161428 3878
rect 161296 3800 161348 3806
rect 161296 3742 161348 3748
rect 161388 3800 161440 3806
rect 161388 3742 161440 3748
rect 160112 3454 160232 3482
rect 160112 480 160140 3454
rect 161308 480 161336 3742
rect 162492 3732 162544 3738
rect 162492 3674 162544 3680
rect 162504 480 162532 3674
rect 163516 3602 163544 53042
rect 163792 32502 163820 63543
rect 163780 32496 163832 32502
rect 163780 32438 163832 32444
rect 163884 31210 163912 68546
rect 163872 31204 163924 31210
rect 163872 31146 163924 31152
rect 163976 24342 164004 69702
rect 163964 24336 164016 24342
rect 163964 24278 164016 24284
rect 164068 22914 164096 69906
rect 164056 22908 164108 22914
rect 164056 22850 164108 22856
rect 164160 11898 164188 73986
rect 164148 11892 164200 11898
rect 164148 11834 164200 11840
rect 164252 11830 164280 78066
rect 164344 76770 164372 79614
rect 164332 76764 164384 76770
rect 164332 76706 164384 76712
rect 164332 76492 164384 76498
rect 164332 76434 164384 76440
rect 164344 63510 164372 76434
rect 164436 63918 164464 79716
rect 164528 76498 164556 79784
rect 164850 79744 164878 79902
rect 164804 79716 164878 79744
rect 164942 79744 164970 80036
rect 165034 79937 165062 80036
rect 165020 79928 165076 79937
rect 165020 79863 165076 79872
rect 165126 79744 165154 80036
rect 164942 79716 165016 79744
rect 164608 79688 164660 79694
rect 164608 79630 164660 79636
rect 164516 76492 164568 76498
rect 164516 76434 164568 76440
rect 164516 76288 164568 76294
rect 164516 76230 164568 76236
rect 164528 66230 164556 76230
rect 164620 68406 164648 79630
rect 164804 78130 164832 79716
rect 164792 78124 164844 78130
rect 164792 78066 164844 78072
rect 164884 77308 164936 77314
rect 164884 77250 164936 77256
rect 164896 77110 164924 77250
rect 164884 77104 164936 77110
rect 164884 77046 164936 77052
rect 164988 76809 165016 79716
rect 165080 79716 165154 79744
rect 164974 76800 165030 76809
rect 164792 76764 164844 76770
rect 164974 76735 165030 76744
rect 164792 76706 164844 76712
rect 164700 76696 164752 76702
rect 164700 76638 164752 76644
rect 164712 68950 164740 76638
rect 164804 69766 164832 76706
rect 165080 76702 165108 79716
rect 165218 79642 165246 80036
rect 165310 79744 165338 80036
rect 165402 79898 165430 80036
rect 165494 79903 165522 80036
rect 165390 79892 165442 79898
rect 165390 79834 165442 79840
rect 165480 79894 165536 79903
rect 165586 79898 165614 80036
rect 165678 79971 165706 80036
rect 165664 79962 165720 79971
rect 165770 79966 165798 80036
rect 165862 79966 165890 80036
rect 165954 79966 165982 80036
rect 166046 79971 166074 80036
rect 165480 79829 165536 79838
rect 165574 79892 165626 79898
rect 165664 79897 165720 79906
rect 165758 79960 165810 79966
rect 165758 79902 165810 79908
rect 165850 79960 165902 79966
rect 165850 79902 165902 79908
rect 165942 79960 165994 79966
rect 165942 79902 165994 79908
rect 166032 79962 166088 79971
rect 166032 79897 166088 79906
rect 165574 79834 165626 79840
rect 165804 79756 165856 79762
rect 165310 79716 165384 79744
rect 165172 79614 165246 79642
rect 165172 78470 165200 79614
rect 165252 79484 165304 79490
rect 165252 79426 165304 79432
rect 165264 79354 165292 79426
rect 165252 79348 165304 79354
rect 165252 79290 165304 79296
rect 165160 78464 165212 78470
rect 165160 78406 165212 78412
rect 165356 77353 165384 79716
rect 166138 79744 166166 80036
rect 166230 79966 166258 80036
rect 166322 79966 166350 80036
rect 166414 79966 166442 80036
rect 166506 79966 166534 80036
rect 166598 79966 166626 80036
rect 166218 79960 166270 79966
rect 166218 79902 166270 79908
rect 166310 79960 166362 79966
rect 166310 79902 166362 79908
rect 166402 79960 166454 79966
rect 166402 79902 166454 79908
rect 166494 79960 166546 79966
rect 166494 79902 166546 79908
rect 166586 79960 166638 79966
rect 166586 79902 166638 79908
rect 165804 79698 165856 79704
rect 166092 79716 166166 79744
rect 166264 79756 166316 79762
rect 165434 79656 165490 79665
rect 165434 79591 165490 79600
rect 165712 79620 165764 79626
rect 165342 77344 165398 77353
rect 165342 77279 165398 77288
rect 165356 76974 165384 77005
rect 165344 76968 165396 76974
rect 165342 76936 165344 76945
rect 165396 76936 165398 76945
rect 165342 76871 165398 76880
rect 165068 76696 165120 76702
rect 165068 76638 165120 76644
rect 165068 74316 165120 74322
rect 165068 74258 165120 74264
rect 164792 69760 164844 69766
rect 164792 69702 164844 69708
rect 164700 68944 164752 68950
rect 164700 68886 164752 68892
rect 164608 68400 164660 68406
rect 164608 68342 164660 68348
rect 164516 66224 164568 66230
rect 164516 66166 164568 66172
rect 164424 63912 164476 63918
rect 164424 63854 164476 63860
rect 164332 63504 164384 63510
rect 164332 63446 164384 63452
rect 165080 42226 165108 74258
rect 165356 70394 165384 76871
rect 165448 76294 165476 79591
rect 165712 79562 165764 79568
rect 165620 79484 165672 79490
rect 165620 79426 165672 79432
rect 165436 76288 165488 76294
rect 165436 76230 165488 76236
rect 165356 70366 165568 70394
rect 165160 69964 165212 69970
rect 165160 69906 165212 69912
rect 165172 69766 165200 69906
rect 165160 69760 165212 69766
rect 165160 69702 165212 69708
rect 165068 42220 165120 42226
rect 165068 42162 165120 42168
rect 165172 29850 165200 69702
rect 165436 68944 165488 68950
rect 165436 68886 165488 68892
rect 165448 68474 165476 68886
rect 165436 68468 165488 68474
rect 165436 68410 165488 68416
rect 165252 66224 165304 66230
rect 165252 66166 165304 66172
rect 165264 66094 165292 66166
rect 165252 66088 165304 66094
rect 165252 66030 165304 66036
rect 165160 29844 165212 29850
rect 165160 29786 165212 29792
rect 165264 24274 165292 66030
rect 165344 64728 165396 64734
rect 165344 64670 165396 64676
rect 165356 63918 165384 64670
rect 165344 63912 165396 63918
rect 165344 63854 165396 63860
rect 165252 24268 165304 24274
rect 165252 24210 165304 24216
rect 165356 14550 165384 63854
rect 165448 15978 165476 68410
rect 165436 15972 165488 15978
rect 165436 15914 165488 15920
rect 165344 14544 165396 14550
rect 165344 14486 165396 14492
rect 164240 11824 164292 11830
rect 164240 11766 164292 11772
rect 165540 9042 165568 70366
rect 165632 53650 165660 79426
rect 165724 75138 165752 79562
rect 165816 76906 165844 79698
rect 165988 79620 166040 79626
rect 165988 79562 166040 79568
rect 165804 76900 165856 76906
rect 165804 76842 165856 76848
rect 165802 76800 165858 76809
rect 165802 76735 165858 76744
rect 165712 75132 165764 75138
rect 165712 75074 165764 75080
rect 165724 74322 165752 75074
rect 165712 74316 165764 74322
rect 165712 74258 165764 74264
rect 165712 74112 165764 74118
rect 165712 74054 165764 74060
rect 165724 64870 165752 74054
rect 165712 64864 165764 64870
rect 165712 64806 165764 64812
rect 165724 63578 165752 64806
rect 165816 64054 165844 76735
rect 165896 76696 165948 76702
rect 165896 76638 165948 76644
rect 165908 66026 165936 76638
rect 166000 68950 166028 79562
rect 166092 76702 166120 79716
rect 166264 79698 166316 79704
rect 166540 79756 166592 79762
rect 166690 79744 166718 80036
rect 166782 79830 166810 80036
rect 166770 79824 166822 79830
rect 166770 79766 166822 79772
rect 166874 79778 166902 80036
rect 166966 79937 166994 80036
rect 167058 79966 167086 80036
rect 167046 79960 167098 79966
rect 166952 79928 167008 79937
rect 167046 79902 167098 79908
rect 166952 79863 167008 79872
rect 166998 79792 167054 79801
rect 166874 79762 166948 79778
rect 166874 79756 166960 79762
rect 166874 79750 166908 79756
rect 166540 79698 166592 79704
rect 166644 79716 166718 79744
rect 166172 79552 166224 79558
rect 166172 79494 166224 79500
rect 166184 79150 166212 79494
rect 166172 79144 166224 79150
rect 166172 79086 166224 79092
rect 166172 76900 166224 76906
rect 166172 76842 166224 76848
rect 166080 76696 166132 76702
rect 166080 76638 166132 76644
rect 166080 76288 166132 76294
rect 166080 76230 166132 76236
rect 166092 69630 166120 76230
rect 166184 69766 166212 76842
rect 166276 71330 166304 79698
rect 166356 76424 166408 76430
rect 166356 76366 166408 76372
rect 166264 71324 166316 71330
rect 166264 71266 166316 71272
rect 166172 69760 166224 69766
rect 166172 69702 166224 69708
rect 166080 69624 166132 69630
rect 166080 69566 166132 69572
rect 165988 68944 166040 68950
rect 165988 68886 166040 68892
rect 165896 66020 165948 66026
rect 165896 65962 165948 65968
rect 165804 64048 165856 64054
rect 165804 63990 165856 63996
rect 165712 63572 165764 63578
rect 165712 63514 165764 63520
rect 166368 60586 166396 76366
rect 166552 74118 166580 79698
rect 166644 79665 166672 79716
rect 167150 79778 167178 80036
rect 167242 79812 167270 80036
rect 167334 79937 167362 80036
rect 167426 79966 167454 80036
rect 167414 79960 167466 79966
rect 167320 79928 167376 79937
rect 167414 79902 167466 79908
rect 167320 79863 167376 79872
rect 167518 79812 167546 80036
rect 167242 79784 167316 79812
rect 166998 79727 167054 79736
rect 167104 79750 167178 79778
rect 166908 79698 166960 79704
rect 166630 79656 166686 79665
rect 166630 79591 166686 79600
rect 166632 79552 166684 79558
rect 166632 79494 166684 79500
rect 166816 79552 166868 79558
rect 166816 79494 166868 79500
rect 166908 79552 166960 79558
rect 166908 79494 166960 79500
rect 166644 75886 166672 79494
rect 166828 76294 166856 79494
rect 166920 77994 166948 79494
rect 166908 77988 166960 77994
rect 166908 77930 166960 77936
rect 166816 76288 166868 76294
rect 166816 76230 166868 76236
rect 166632 75880 166684 75886
rect 166632 75822 166684 75828
rect 166540 74112 166592 74118
rect 166540 74054 166592 74060
rect 166540 64660 166592 64666
rect 166540 64602 166592 64608
rect 166552 64054 166580 64602
rect 166540 64048 166592 64054
rect 166540 63990 166592 63996
rect 166448 63572 166500 63578
rect 166448 63514 166500 63520
rect 166356 60580 166408 60586
rect 166356 60522 166408 60528
rect 165620 53644 165672 53650
rect 165620 53586 165672 53592
rect 166460 35358 166488 63514
rect 166448 35352 166500 35358
rect 166448 35294 166500 35300
rect 166552 21418 166580 63990
rect 166644 28354 166672 75822
rect 166908 71324 166960 71330
rect 166908 71266 166960 71272
rect 166724 69624 166776 69630
rect 166724 69566 166776 69572
rect 166736 69494 166764 69566
rect 166724 69488 166776 69494
rect 166724 69430 166776 69436
rect 166632 28348 166684 28354
rect 166632 28290 166684 28296
rect 166540 21412 166592 21418
rect 166540 21354 166592 21360
rect 166736 15910 166764 69430
rect 166816 68944 166868 68950
rect 166816 68886 166868 68892
rect 166828 68814 166856 68886
rect 166816 68808 166868 68814
rect 166816 68750 166868 68756
rect 166724 15904 166776 15910
rect 166724 15846 166776 15852
rect 166828 10402 166856 68750
rect 166816 10396 166868 10402
rect 166816 10338 166868 10344
rect 165528 9036 165580 9042
rect 165528 8978 165580 8984
rect 166920 7682 166948 71266
rect 167012 49706 167040 79727
rect 167104 79642 167132 79750
rect 167104 79614 167224 79642
rect 167196 77790 167224 79614
rect 167288 78878 167316 79784
rect 167472 79784 167546 79812
rect 167368 79688 167420 79694
rect 167368 79630 167420 79636
rect 167276 78872 167328 78878
rect 167276 78814 167328 78820
rect 167184 77784 167236 77790
rect 167184 77726 167236 77732
rect 167380 77518 167408 79630
rect 167368 77512 167420 77518
rect 167368 77454 167420 77460
rect 167368 76764 167420 76770
rect 167368 76706 167420 76712
rect 167184 76696 167236 76702
rect 167184 76638 167236 76644
rect 167092 74588 167144 74594
rect 167092 74530 167144 74536
rect 167000 49700 167052 49706
rect 167000 49642 167052 49648
rect 167000 46232 167052 46238
rect 167000 46174 167052 46180
rect 167012 16574 167040 46174
rect 167104 39438 167132 74530
rect 167196 56574 167224 76638
rect 167276 74112 167328 74118
rect 167276 74054 167328 74060
rect 167288 62082 167316 74054
rect 167380 68950 167408 76706
rect 167472 76702 167500 79784
rect 167610 79744 167638 80036
rect 167702 79801 167730 80036
rect 167564 79716 167638 79744
rect 167688 79792 167744 79801
rect 167688 79727 167744 79736
rect 167794 79744 167822 80036
rect 167886 79937 167914 80036
rect 167872 79928 167928 79937
rect 167872 79863 167928 79872
rect 167978 79744 168006 80036
rect 168070 79801 168098 80036
rect 167794 79716 167868 79744
rect 167564 76770 167592 79716
rect 167644 79620 167696 79626
rect 167644 79562 167696 79568
rect 167552 76764 167604 76770
rect 167552 76706 167604 76712
rect 167460 76696 167512 76702
rect 167460 76638 167512 76644
rect 167656 73154 167684 79562
rect 167736 79484 167788 79490
rect 167736 79426 167788 79432
rect 167748 79014 167776 79426
rect 167736 79008 167788 79014
rect 167736 78950 167788 78956
rect 167748 74594 167776 78950
rect 167840 76809 167868 79716
rect 167932 79716 168006 79744
rect 168056 79792 168112 79801
rect 168056 79727 168112 79736
rect 168162 79744 168190 80036
rect 168254 79971 168282 80036
rect 168240 79962 168296 79971
rect 168346 79966 168374 80036
rect 168438 79966 168466 80036
rect 168530 79966 168558 80036
rect 168240 79897 168296 79906
rect 168334 79960 168386 79966
rect 168334 79902 168386 79908
rect 168426 79960 168478 79966
rect 168426 79902 168478 79908
rect 168518 79960 168570 79966
rect 168622 79937 168650 80036
rect 168518 79902 168570 79908
rect 168608 79928 168664 79937
rect 168608 79863 168664 79872
rect 168714 79801 168742 80036
rect 168806 79830 168834 80036
rect 168794 79824 168846 79830
rect 168378 79792 168434 79801
rect 168288 79756 168340 79762
rect 168162 79716 168236 79744
rect 167932 78305 167960 79716
rect 167918 78296 167974 78305
rect 167918 78231 167974 78240
rect 167826 76800 167882 76809
rect 167826 76735 167882 76744
rect 167736 74588 167788 74594
rect 167736 74530 167788 74536
rect 168208 74118 168236 79716
rect 168378 79727 168434 79736
rect 168700 79792 168756 79801
rect 168898 79812 168926 80036
rect 168990 79937 169018 80036
rect 168976 79928 169032 79937
rect 169082 79898 169110 80036
rect 168976 79863 169032 79872
rect 169070 79892 169122 79898
rect 169070 79834 169122 79840
rect 168898 79784 168972 79812
rect 168794 79766 168846 79772
rect 168944 79778 168972 79784
rect 168944 79750 169064 79778
rect 168700 79727 168756 79736
rect 168288 79698 168340 79704
rect 168300 77926 168328 79698
rect 168288 77920 168340 77926
rect 168288 77862 168340 77868
rect 168286 76936 168342 76945
rect 168286 76871 168342 76880
rect 168300 74322 168328 76871
rect 168288 74316 168340 74322
rect 168288 74258 168340 74264
rect 168196 74112 168248 74118
rect 168196 74054 168248 74060
rect 168196 73976 168248 73982
rect 168196 73918 168248 73924
rect 167920 73636 167972 73642
rect 167920 73578 167972 73584
rect 167472 73126 167684 73154
rect 167368 68944 167420 68950
rect 167368 68886 167420 68892
rect 167472 68882 167500 73126
rect 167460 68876 167512 68882
rect 167460 68818 167512 68824
rect 167276 62076 167328 62082
rect 167276 62018 167328 62024
rect 167184 56568 167236 56574
rect 167184 56510 167236 56516
rect 167932 55078 167960 73578
rect 168208 70394 168236 73918
rect 168024 70378 168236 70394
rect 168012 70372 168236 70378
rect 168064 70366 168236 70372
rect 168012 70314 168064 70320
rect 168196 68944 168248 68950
rect 168196 68886 168248 68892
rect 168104 68876 168156 68882
rect 168104 68818 168156 68824
rect 167920 55072 167972 55078
rect 167920 55014 167972 55020
rect 167092 39432 167144 39438
rect 167092 39374 167144 39380
rect 168116 17406 168144 68818
rect 168104 17400 168156 17406
rect 168104 17342 168156 17348
rect 167012 16546 167224 16574
rect 166908 7676 166960 7682
rect 166908 7618 166960 7624
rect 163688 3868 163740 3874
rect 163688 3810 163740 3816
rect 163504 3596 163556 3602
rect 163504 3538 163556 3544
rect 163700 480 163728 3810
rect 166080 3664 166132 3670
rect 166080 3606 166132 3612
rect 164884 3596 164936 3602
rect 164884 3538 164936 3544
rect 164896 480 164924 3538
rect 166092 480 166120 3606
rect 167196 480 167224 16546
rect 168208 6322 168236 68886
rect 168196 6316 168248 6322
rect 168196 6258 168248 6264
rect 168300 4894 168328 74258
rect 168392 52290 168420 79727
rect 168472 79688 168524 79694
rect 168472 79630 168524 79636
rect 168564 79688 168616 79694
rect 168564 79630 168616 79636
rect 168932 79688 168984 79694
rect 168932 79630 168984 79636
rect 168484 79529 168512 79630
rect 168470 79520 168526 79529
rect 168470 79455 168526 79464
rect 168470 79248 168526 79257
rect 168470 79183 168526 79192
rect 168380 52284 168432 52290
rect 168380 52226 168432 52232
rect 168380 49020 168432 49026
rect 168380 48962 168432 48968
rect 168288 4888 168340 4894
rect 168288 4830 168340 4836
rect 168392 3602 168420 48962
rect 168484 38010 168512 79183
rect 168576 78441 168604 79630
rect 168656 79620 168708 79626
rect 168656 79562 168708 79568
rect 168562 78432 168618 78441
rect 168562 78367 168618 78376
rect 168564 76696 168616 76702
rect 168564 76638 168616 76644
rect 168576 64530 168604 76638
rect 168668 66230 168696 79562
rect 168746 79520 168802 79529
rect 168746 79455 168802 79464
rect 168760 68746 168788 79455
rect 168944 75313 168972 79630
rect 169036 76401 169064 79750
rect 169174 79744 169202 80036
rect 169128 79716 169202 79744
rect 169266 79744 169294 80036
rect 169358 79966 169386 80036
rect 169346 79960 169398 79966
rect 169346 79902 169398 79908
rect 169450 79778 169478 80036
rect 169404 79762 169478 79778
rect 169392 79756 169478 79762
rect 169266 79716 169340 79744
rect 169128 76702 169156 79716
rect 169208 79620 169260 79626
rect 169208 79562 169260 79568
rect 169220 79257 169248 79562
rect 169206 79248 169262 79257
rect 169206 79183 169262 79192
rect 169312 76809 169340 79716
rect 169444 79750 169478 79756
rect 169542 79778 169570 80036
rect 169634 79937 169662 80036
rect 169620 79928 169676 79937
rect 169620 79863 169676 79872
rect 169542 79750 169616 79778
rect 169392 79698 169444 79704
rect 169482 79656 169538 79665
rect 169482 79591 169538 79600
rect 169392 78124 169444 78130
rect 169392 78066 169444 78072
rect 169298 76800 169354 76809
rect 169298 76735 169354 76744
rect 169116 76696 169168 76702
rect 169116 76638 169168 76644
rect 169022 76392 169078 76401
rect 169022 76327 169078 76336
rect 168930 75304 168986 75313
rect 168930 75239 168986 75248
rect 169036 73154 169064 76327
rect 169036 73126 169156 73154
rect 169128 71774 169156 73126
rect 169128 71746 169340 71774
rect 169208 70780 169260 70786
rect 169208 70722 169260 70728
rect 168748 68740 168800 68746
rect 168748 68682 168800 68688
rect 168656 66224 168708 66230
rect 168656 66166 168708 66172
rect 168564 64524 168616 64530
rect 168564 64466 168616 64472
rect 168564 38208 168616 38214
rect 168564 38150 168616 38156
rect 168472 38004 168524 38010
rect 168472 37946 168524 37952
rect 168576 6914 168604 38150
rect 169220 17338 169248 70722
rect 169312 47598 169340 71746
rect 169404 70786 169432 78066
rect 169496 73137 169524 79591
rect 169588 78130 169616 79750
rect 169726 79744 169754 80036
rect 169818 79971 169846 80036
rect 169804 79962 169860 79971
rect 169910 79966 169938 80036
rect 170002 79966 170030 80036
rect 170094 79966 170122 80036
rect 169804 79897 169860 79906
rect 169898 79960 169950 79966
rect 169898 79902 169950 79908
rect 169990 79960 170042 79966
rect 169990 79902 170042 79908
rect 170082 79960 170134 79966
rect 170082 79902 170134 79908
rect 170036 79824 170088 79830
rect 170186 79778 170214 80036
rect 170278 79830 170306 80036
rect 170370 79937 170398 80036
rect 170462 79966 170490 80036
rect 170450 79960 170502 79966
rect 170356 79928 170412 79937
rect 170554 79937 170582 80036
rect 170450 79902 170502 79908
rect 170540 79928 170596 79937
rect 170356 79863 170412 79872
rect 170540 79863 170596 79872
rect 170036 79766 170088 79772
rect 169680 79716 169754 79744
rect 169944 79756 169996 79762
rect 169576 78124 169628 78130
rect 169576 78066 169628 78072
rect 169680 77489 169708 79716
rect 169944 79698 169996 79704
rect 169850 79520 169906 79529
rect 169850 79455 169906 79464
rect 169864 79404 169892 79455
rect 169772 79376 169892 79404
rect 169772 78946 169800 79376
rect 169760 78940 169812 78946
rect 169760 78882 169812 78888
rect 169666 77480 169722 77489
rect 169666 77415 169722 77424
rect 169482 73128 169538 73137
rect 169482 73063 169538 73072
rect 169392 70780 169444 70786
rect 169392 70722 169444 70728
rect 169392 68740 169444 68746
rect 169392 68682 169444 68688
rect 169300 47592 169352 47598
rect 169300 47534 169352 47540
rect 169404 39506 169432 68682
rect 169392 39500 169444 39506
rect 169392 39442 169444 39448
rect 169496 38078 169524 73063
rect 169576 66224 169628 66230
rect 169576 66166 169628 66172
rect 169588 65754 169616 66166
rect 169576 65748 169628 65754
rect 169576 65690 169628 65696
rect 169484 38072 169536 38078
rect 169484 38014 169536 38020
rect 169588 29782 169616 65690
rect 169576 29776 169628 29782
rect 169576 29718 169628 29724
rect 169208 17332 169260 17338
rect 169208 17274 169260 17280
rect 169772 14482 169800 78882
rect 169956 78674 169984 79698
rect 170048 79540 170076 79766
rect 170140 79750 170214 79778
rect 170266 79824 170318 79830
rect 170266 79766 170318 79772
rect 170140 79665 170168 79750
rect 170220 79688 170272 79694
rect 170126 79656 170182 79665
rect 170370 79676 170398 79863
rect 170646 79812 170674 80036
rect 170738 79971 170766 80036
rect 170724 79962 170780 79971
rect 170724 79897 170780 79906
rect 170830 79898 170858 80036
rect 170922 79966 170950 80036
rect 171014 79966 171042 80036
rect 170910 79960 170962 79966
rect 170910 79902 170962 79908
rect 171002 79960 171054 79966
rect 171002 79902 171054 79908
rect 170818 79892 170870 79898
rect 170818 79834 170870 79840
rect 170646 79784 170720 79812
rect 170496 79756 170548 79762
rect 170496 79698 170548 79704
rect 170220 79630 170272 79636
rect 170324 79648 170398 79676
rect 170126 79591 170182 79600
rect 170048 79512 170168 79540
rect 169944 78668 169996 78674
rect 169944 78610 169996 78616
rect 169944 78532 169996 78538
rect 169944 78474 169996 78480
rect 169956 77654 169984 78474
rect 169944 77648 169996 77654
rect 169944 77590 169996 77596
rect 169944 77444 169996 77450
rect 169944 77386 169996 77392
rect 169852 76900 169904 76906
rect 169852 76842 169904 76848
rect 169864 33862 169892 76842
rect 169956 40866 169984 77386
rect 170036 77036 170088 77042
rect 170036 76978 170088 76984
rect 170048 42158 170076 76978
rect 170140 57866 170168 79512
rect 170232 73982 170260 79630
rect 170324 76906 170352 79648
rect 170508 78577 170536 79698
rect 170588 79552 170640 79558
rect 170692 79529 170720 79784
rect 171106 79744 171134 80036
rect 171060 79716 171134 79744
rect 171198 79744 171226 80036
rect 171290 79937 171318 80036
rect 171382 79966 171410 80036
rect 171370 79960 171422 79966
rect 171276 79928 171332 79937
rect 171370 79902 171422 79908
rect 171276 79863 171332 79872
rect 171324 79824 171376 79830
rect 171324 79766 171376 79772
rect 171198 79716 171272 79744
rect 170956 79688 171008 79694
rect 170956 79630 171008 79636
rect 170772 79620 170824 79626
rect 170772 79562 170824 79568
rect 170588 79494 170640 79500
rect 170678 79520 170734 79529
rect 170494 78568 170550 78577
rect 170494 78503 170550 78512
rect 170496 77988 170548 77994
rect 170496 77930 170548 77936
rect 170508 77858 170536 77930
rect 170496 77852 170548 77858
rect 170496 77794 170548 77800
rect 170312 76900 170364 76906
rect 170312 76842 170364 76848
rect 170600 75682 170628 79494
rect 170678 79455 170734 79464
rect 170692 77450 170720 79455
rect 170784 79393 170812 79562
rect 170770 79384 170826 79393
rect 170770 79319 170826 79328
rect 170680 77444 170732 77450
rect 170680 77386 170732 77392
rect 170784 77042 170812 79319
rect 170864 79280 170916 79286
rect 170864 79222 170916 79228
rect 170876 77586 170904 79222
rect 170864 77580 170916 77586
rect 170864 77522 170916 77528
rect 170772 77036 170824 77042
rect 170772 76978 170824 76984
rect 170862 76800 170918 76809
rect 170862 76735 170918 76744
rect 170588 75676 170640 75682
rect 170588 75618 170640 75624
rect 170220 73976 170272 73982
rect 170220 73918 170272 73924
rect 170220 66156 170272 66162
rect 170220 66098 170272 66104
rect 170232 65890 170260 66098
rect 170220 65884 170272 65890
rect 170220 65826 170272 65832
rect 170128 57860 170180 57866
rect 170128 57802 170180 57808
rect 170404 55888 170456 55894
rect 170404 55830 170456 55836
rect 170036 42152 170088 42158
rect 170036 42094 170088 42100
rect 169944 40860 169996 40866
rect 169944 40802 169996 40808
rect 169852 33856 169904 33862
rect 169852 33798 169904 33804
rect 169760 14476 169812 14482
rect 169760 14418 169812 14424
rect 168484 6886 168604 6914
rect 168380 3596 168432 3602
rect 168380 3538 168432 3544
rect 168484 3482 168512 6886
rect 170416 3874 170444 55830
rect 170876 36650 170904 76735
rect 170968 75993 170996 79630
rect 171060 78742 171088 79716
rect 171140 79620 171192 79626
rect 171140 79562 171192 79568
rect 171152 78849 171180 79562
rect 171244 79218 171272 79716
rect 171232 79212 171284 79218
rect 171232 79154 171284 79160
rect 171138 78840 171194 78849
rect 171138 78775 171194 78784
rect 171048 78736 171100 78742
rect 171048 78678 171100 78684
rect 171046 78568 171102 78577
rect 171046 78503 171102 78512
rect 170954 75984 171010 75993
rect 170954 75919 171010 75928
rect 171060 75800 171088 78503
rect 171140 78328 171192 78334
rect 171140 78270 171192 78276
rect 171152 78130 171180 78270
rect 171140 78124 171192 78130
rect 171140 78066 171192 78072
rect 171244 77194 171272 79154
rect 171336 78130 171364 79766
rect 171474 79642 171502 80036
rect 171566 79744 171594 80036
rect 171658 79966 171686 80036
rect 171750 79966 171778 80036
rect 171646 79960 171698 79966
rect 171646 79902 171698 79908
rect 171738 79960 171790 79966
rect 171738 79902 171790 79908
rect 171842 79812 171870 80036
rect 171934 79966 171962 80036
rect 171922 79960 171974 79966
rect 171922 79902 171974 79908
rect 172026 79898 172054 80036
rect 172014 79892 172066 79898
rect 172014 79834 172066 79840
rect 171704 79784 171870 79812
rect 171566 79716 171640 79744
rect 171428 79614 171502 79642
rect 171428 79121 171456 79614
rect 171414 79112 171470 79121
rect 171414 79047 171470 79056
rect 171324 78124 171376 78130
rect 171324 78066 171376 78072
rect 171244 77166 171364 77194
rect 171232 77036 171284 77042
rect 171232 76978 171284 76984
rect 171140 76696 171192 76702
rect 171140 76638 171192 76644
rect 170968 75772 171088 75800
rect 170968 73001 170996 75772
rect 171048 75676 171100 75682
rect 171048 75618 171100 75624
rect 170954 72992 171010 73001
rect 170954 72927 171010 72936
rect 170864 36644 170916 36650
rect 170864 36586 170916 36592
rect 170968 32434 170996 72927
rect 170956 32428 171008 32434
rect 170956 32370 171008 32376
rect 171060 13122 171088 75618
rect 171152 26994 171180 76638
rect 171244 29714 171272 76978
rect 171336 40798 171364 77166
rect 171428 77042 171456 79047
rect 171508 78600 171560 78606
rect 171508 78542 171560 78548
rect 171416 77036 171468 77042
rect 171416 76978 171468 76984
rect 171520 75290 171548 78542
rect 171428 75262 171548 75290
rect 171428 64462 171456 75262
rect 171612 71774 171640 79716
rect 171704 75585 171732 79784
rect 172118 79744 172146 80036
rect 172072 79716 172146 79744
rect 171966 79656 172022 79665
rect 171784 79620 171836 79626
rect 171966 79591 171968 79600
rect 171784 79562 171836 79568
rect 172020 79591 172022 79600
rect 171968 79562 172020 79568
rect 171796 76158 171824 79562
rect 171876 79484 171928 79490
rect 171876 79426 171928 79432
rect 171888 78169 171916 79426
rect 171874 78160 171930 78169
rect 171874 78095 171930 78104
rect 171980 76702 172008 79562
rect 171968 76696 172020 76702
rect 171968 76638 172020 76644
rect 172072 76514 172100 79716
rect 172210 79676 172238 80036
rect 172302 79744 172330 80036
rect 172394 79966 172422 80036
rect 172382 79960 172434 79966
rect 172486 79937 172514 80036
rect 172578 79966 172606 80036
rect 172670 79966 172698 80036
rect 172762 79966 172790 80036
rect 172566 79960 172618 79966
rect 172382 79902 172434 79908
rect 172472 79928 172528 79937
rect 172566 79902 172618 79908
rect 172658 79960 172710 79966
rect 172658 79902 172710 79908
rect 172750 79960 172802 79966
rect 172750 79902 172802 79908
rect 172472 79863 172528 79872
rect 172520 79824 172572 79830
rect 172518 79792 172520 79801
rect 172854 79812 172882 80036
rect 172572 79792 172574 79801
rect 172808 79784 172882 79812
rect 172946 79812 172974 80036
rect 173038 79966 173066 80036
rect 173026 79960 173078 79966
rect 173026 79902 173078 79908
rect 173130 79812 173158 80036
rect 172946 79784 173020 79812
rect 173084 79801 173158 79812
rect 172808 79778 172836 79784
rect 172428 79756 172480 79762
rect 172302 79716 172376 79744
rect 172210 79648 172284 79676
rect 172152 79552 172204 79558
rect 172152 79494 172204 79500
rect 171980 76486 172100 76514
rect 171784 76152 171836 76158
rect 171784 76094 171836 76100
rect 171690 75576 171746 75585
rect 171690 75511 171746 75520
rect 171520 71746 171640 71774
rect 171520 70009 171548 71746
rect 171980 70394 172008 76486
rect 172164 75177 172192 79494
rect 172256 78606 172284 79648
rect 172244 78600 172296 78606
rect 172244 78542 172296 78548
rect 172150 75168 172206 75177
rect 172150 75103 172206 75112
rect 172164 71774 172192 75103
rect 172348 73953 172376 79716
rect 172518 79727 172574 79736
rect 172716 79750 172836 79778
rect 172428 79698 172480 79704
rect 172440 78266 172468 79698
rect 172520 79620 172572 79626
rect 172520 79562 172572 79568
rect 172428 78260 172480 78266
rect 172428 78202 172480 78208
rect 172428 76696 172480 76702
rect 172428 76638 172480 76644
rect 172440 76158 172468 76638
rect 172428 76152 172480 76158
rect 172428 76094 172480 76100
rect 172334 73944 172390 73953
rect 172334 73879 172390 73888
rect 171704 70366 172008 70394
rect 172072 71746 172192 71774
rect 171506 70000 171562 70009
rect 171506 69935 171562 69944
rect 171704 69873 171732 70366
rect 171690 69864 171746 69873
rect 171690 69799 171746 69808
rect 171416 64456 171468 64462
rect 171416 64398 171468 64404
rect 172072 49026 172100 71746
rect 172150 70000 172206 70009
rect 172150 69935 172206 69944
rect 172060 49020 172112 49026
rect 172060 48962 172112 48968
rect 172164 42090 172192 69935
rect 172242 69864 172298 69873
rect 172242 69799 172298 69808
rect 172152 42084 172204 42090
rect 172152 42026 172204 42032
rect 171324 40792 171376 40798
rect 171324 40734 171376 40740
rect 171232 29708 171284 29714
rect 171232 29650 171284 29656
rect 171140 26988 171192 26994
rect 171140 26930 171192 26936
rect 172256 26926 172284 69799
rect 172244 26920 172296 26926
rect 172244 26862 172296 26868
rect 172348 25634 172376 73879
rect 172440 28286 172468 76094
rect 172532 53718 172560 79562
rect 172612 79484 172664 79490
rect 172612 79426 172664 79432
rect 172624 67590 172652 79426
rect 172716 77024 172744 79750
rect 172716 76996 172836 77024
rect 172808 76945 172836 76996
rect 172794 76936 172850 76945
rect 172704 76900 172756 76906
rect 172794 76871 172850 76880
rect 172704 76842 172756 76848
rect 172612 67584 172664 67590
rect 172612 67526 172664 67532
rect 172716 67454 172744 76842
rect 172992 75750 173020 79784
rect 173070 79792 173158 79801
rect 173126 79784 173158 79792
rect 173070 79727 173126 79736
rect 173222 79744 173250 80036
rect 173314 79966 173342 80036
rect 173302 79960 173354 79966
rect 173302 79902 173354 79908
rect 173406 79830 173434 80036
rect 173394 79824 173446 79830
rect 173394 79766 173446 79772
rect 173498 79744 173526 80036
rect 173590 79966 173618 80036
rect 173578 79960 173630 79966
rect 173578 79902 173630 79908
rect 173682 79812 173710 80036
rect 173774 79898 173802 80036
rect 173866 79971 173894 80036
rect 173852 79962 173908 79971
rect 173958 79966 173986 80036
rect 173762 79892 173814 79898
rect 173852 79897 173908 79906
rect 173946 79960 173998 79966
rect 173946 79902 173998 79908
rect 173762 79834 173814 79840
rect 173636 79784 173710 79812
rect 173222 79716 173296 79744
rect 173498 79716 173572 79744
rect 173072 79688 173124 79694
rect 173072 79630 173124 79636
rect 172980 75744 173032 75750
rect 172980 75686 173032 75692
rect 173084 74866 173112 79630
rect 173164 79620 173216 79626
rect 173164 79562 173216 79568
rect 173176 75002 173204 79562
rect 173268 75857 173296 79716
rect 173440 79620 173492 79626
rect 173440 79562 173492 79568
rect 173348 75948 173400 75954
rect 173348 75890 173400 75896
rect 173254 75848 173310 75857
rect 173254 75783 173310 75792
rect 173164 74996 173216 75002
rect 173164 74938 173216 74944
rect 173072 74860 173124 74866
rect 173072 74802 173124 74808
rect 173360 71641 173388 75890
rect 173452 75449 173480 79562
rect 173544 76906 173572 79716
rect 173532 76900 173584 76906
rect 173532 76842 173584 76848
rect 173636 75954 173664 79784
rect 174050 79744 174078 80036
rect 174004 79716 174078 79744
rect 174142 79744 174170 80036
rect 174234 79937 174262 80036
rect 174220 79928 174276 79937
rect 174220 79863 174222 79872
rect 174274 79863 174276 79872
rect 174222 79834 174274 79840
rect 174234 79803 174262 79834
rect 174326 79744 174354 80036
rect 174142 79716 174216 79744
rect 173716 79688 173768 79694
rect 174004 79665 174032 79716
rect 173716 79630 173768 79636
rect 173990 79656 174046 79665
rect 173624 75948 173676 75954
rect 173624 75890 173676 75896
rect 173728 75562 173756 79630
rect 173990 79591 174046 79600
rect 173900 79552 173952 79558
rect 173900 79494 173952 79500
rect 173912 78985 173940 79494
rect 173992 79484 174044 79490
rect 173992 79426 174044 79432
rect 173898 78976 173954 78985
rect 173898 78911 173954 78920
rect 173806 76936 173862 76945
rect 173806 76871 173862 76880
rect 173544 75534 173756 75562
rect 173438 75440 173494 75449
rect 173438 75375 173494 75384
rect 173544 75290 173572 75534
rect 173714 75440 173770 75449
rect 173714 75375 173770 75384
rect 173452 75262 173572 75290
rect 173346 71632 173402 71641
rect 173346 71567 173402 71576
rect 173452 70394 173480 75262
rect 173532 74996 173584 75002
rect 173532 74938 173584 74944
rect 173544 73681 173572 74938
rect 173728 73914 173756 75375
rect 173716 73908 173768 73914
rect 173716 73850 173768 73856
rect 173530 73672 173586 73681
rect 173530 73607 173586 73616
rect 172808 70366 173480 70394
rect 172808 67522 172836 70366
rect 172796 67516 172848 67522
rect 172796 67458 172848 67464
rect 172704 67448 172756 67454
rect 172704 67390 172756 67396
rect 173440 67448 173492 67454
rect 173440 67390 173492 67396
rect 173452 66706 173480 67390
rect 173440 66700 173492 66706
rect 173440 66642 173492 66648
rect 172520 53712 172572 53718
rect 172520 53654 172572 53660
rect 173452 36582 173480 66642
rect 173544 39370 173572 73607
rect 173624 67516 173676 67522
rect 173624 67458 173676 67464
rect 173636 66774 173664 67458
rect 173624 66768 173676 66774
rect 173624 66710 173676 66716
rect 173532 39364 173584 39370
rect 173532 39306 173584 39312
rect 173440 36576 173492 36582
rect 173440 36518 173492 36524
rect 172428 28280 172480 28286
rect 172428 28222 172480 28228
rect 172336 25628 172388 25634
rect 172336 25570 172388 25576
rect 173636 25566 173664 66710
rect 171784 25560 171836 25566
rect 171784 25502 171836 25508
rect 173624 25560 173676 25566
rect 173624 25502 173676 25508
rect 171048 13116 171100 13122
rect 171048 13058 171100 13064
rect 170404 3868 170456 3874
rect 170404 3810 170456 3816
rect 170772 3732 170824 3738
rect 170772 3674 170824 3680
rect 169576 3596 169628 3602
rect 169576 3538 169628 3544
rect 168392 3454 168512 3482
rect 168392 480 168420 3454
rect 169588 480 169616 3538
rect 170784 480 170812 3674
rect 171796 2922 171824 25502
rect 173728 22846 173756 73850
rect 173820 24206 173848 76871
rect 173808 24200 173860 24206
rect 173808 24142 173860 24148
rect 173716 22840 173768 22846
rect 173716 22782 173768 22788
rect 171874 22672 171930 22681
rect 171874 22607 171930 22616
rect 171888 3126 171916 22607
rect 173912 4826 173940 78911
rect 174004 7614 174032 79426
rect 174188 77314 174216 79716
rect 174280 79716 174354 79744
rect 174418 79744 174446 80036
rect 174510 79898 174538 80036
rect 174498 79892 174550 79898
rect 174498 79834 174550 79840
rect 174602 79744 174630 80036
rect 174694 79812 174722 80036
rect 174786 79966 174814 80036
rect 174878 79971 174906 80036
rect 174774 79960 174826 79966
rect 174774 79902 174826 79908
rect 174864 79962 174920 79971
rect 174864 79897 174920 79906
rect 174970 79898 174998 80036
rect 175062 79966 175090 80036
rect 175154 79966 175182 80036
rect 175246 79966 175274 80036
rect 175050 79960 175102 79966
rect 175050 79902 175102 79908
rect 175142 79960 175194 79966
rect 175142 79902 175194 79908
rect 175234 79960 175286 79966
rect 175338 79937 175366 80036
rect 175430 79966 175458 80036
rect 175522 79966 175550 80036
rect 175418 79960 175470 79966
rect 175234 79902 175286 79908
rect 175324 79928 175380 79937
rect 174958 79892 175010 79898
rect 175418 79902 175470 79908
rect 175510 79960 175562 79966
rect 175510 79902 175562 79908
rect 175324 79863 175380 79872
rect 174958 79834 175010 79840
rect 174694 79801 174768 79812
rect 174694 79792 174782 79801
rect 174694 79784 174726 79792
rect 174418 79716 174492 79744
rect 174602 79716 174676 79744
rect 174910 79792 174966 79801
rect 174726 79727 174782 79736
rect 174820 79756 174872 79762
rect 174176 77308 174228 77314
rect 174176 77250 174228 77256
rect 174280 77194 174308 79716
rect 174360 79416 174412 79422
rect 174360 79358 174412 79364
rect 174372 77586 174400 79358
rect 174360 77580 174412 77586
rect 174360 77522 174412 77528
rect 174096 77166 174308 77194
rect 174096 67386 174124 77166
rect 174176 77036 174228 77042
rect 174176 76978 174228 76984
rect 174188 67454 174216 76978
rect 174268 76764 174320 76770
rect 174268 76706 174320 76712
rect 174280 67522 174308 76706
rect 174464 71505 174492 79716
rect 174544 79620 174596 79626
rect 174544 79562 174596 79568
rect 174556 75449 174584 79562
rect 174648 76265 174676 79716
rect 174910 79727 174966 79736
rect 175004 79756 175056 79762
rect 174820 79698 174872 79704
rect 174728 78736 174780 78742
rect 174728 78678 174780 78684
rect 174634 76256 174690 76265
rect 174634 76191 174690 76200
rect 174542 75440 174598 75449
rect 174542 75375 174598 75384
rect 174740 71777 174768 78678
rect 174832 77217 174860 79698
rect 174818 77208 174874 77217
rect 174818 77143 174874 77152
rect 174924 77042 174952 79727
rect 175004 79698 175056 79704
rect 175188 79756 175240 79762
rect 175614 79744 175642 80036
rect 175706 79778 175734 80036
rect 175798 79898 175826 80036
rect 175786 79892 175838 79898
rect 175786 79834 175838 79840
rect 175706 79750 175780 79778
rect 175188 79698 175240 79704
rect 175568 79716 175642 79744
rect 174912 77036 174964 77042
rect 174912 76978 174964 76984
rect 174910 75440 174966 75449
rect 174910 75375 174966 75384
rect 174726 71768 174782 71777
rect 174726 71703 174782 71712
rect 174450 71496 174506 71505
rect 174450 71431 174506 71440
rect 174268 67516 174320 67522
rect 174268 67458 174320 67464
rect 174728 67516 174780 67522
rect 174728 67458 174780 67464
rect 174176 67448 174228 67454
rect 174176 67390 174228 67396
rect 174084 67380 174136 67386
rect 174084 67322 174136 67328
rect 174740 66842 174768 67458
rect 174820 67380 174872 67386
rect 174820 67322 174872 67328
rect 174832 67250 174860 67322
rect 174820 67244 174872 67250
rect 174820 67186 174872 67192
rect 174728 66836 174780 66842
rect 174728 66778 174780 66784
rect 174740 40730 174768 66778
rect 174728 40724 174780 40730
rect 174728 40666 174780 40672
rect 174832 35290 174860 67186
rect 174924 37942 174952 75375
rect 175016 72865 175044 79698
rect 175094 78840 175150 78849
rect 175094 78775 175150 78784
rect 175108 75818 175136 78775
rect 175200 76770 175228 79698
rect 175568 79676 175596 79716
rect 175384 79665 175596 79676
rect 175384 79656 175610 79665
rect 175384 79648 175554 79656
rect 175280 79620 175332 79626
rect 175280 79562 175332 79568
rect 175188 76764 175240 76770
rect 175188 76706 175240 76712
rect 175096 75812 175148 75818
rect 175096 75754 175148 75760
rect 175292 74050 175320 79562
rect 175280 74044 175332 74050
rect 175280 73986 175332 73992
rect 175292 73154 175320 73986
rect 175108 73126 175320 73154
rect 175002 72856 175058 72865
rect 175002 72791 175058 72800
rect 175004 67448 175056 67454
rect 175004 67390 175056 67396
rect 175016 67318 175044 67390
rect 175004 67312 175056 67318
rect 175004 67254 175056 67260
rect 174912 37936 174964 37942
rect 174912 37878 174964 37884
rect 174820 35284 174872 35290
rect 174820 35226 174872 35232
rect 175016 24138 175044 67254
rect 175004 24132 175056 24138
rect 175004 24074 175056 24080
rect 175108 11762 175136 73126
rect 175186 72856 175242 72865
rect 175186 72791 175242 72800
rect 175096 11756 175148 11762
rect 175096 11698 175148 11704
rect 175200 10334 175228 72791
rect 175188 10328 175240 10334
rect 175188 10270 175240 10276
rect 175384 8974 175412 79648
rect 175554 79591 175610 79600
rect 175556 79552 175608 79558
rect 175556 79494 175608 79500
rect 175464 79484 175516 79490
rect 175464 79426 175516 79432
rect 175476 77042 175504 79426
rect 175568 78112 175596 79494
rect 175568 78084 175688 78112
rect 175556 77988 175608 77994
rect 175556 77930 175608 77936
rect 175464 77036 175516 77042
rect 175464 76978 175516 76984
rect 175464 76900 175516 76906
rect 175464 76842 175516 76848
rect 175476 61878 175504 76842
rect 175568 67386 175596 77930
rect 175660 67522 175688 78084
rect 175752 77761 175780 79750
rect 175890 79608 175918 80036
rect 175982 79966 176010 80036
rect 175970 79960 176022 79966
rect 175970 79902 176022 79908
rect 176074 79801 176102 80036
rect 176060 79792 176116 79801
rect 176166 79778 176194 80036
rect 176258 79898 176286 80036
rect 176350 79898 176378 80036
rect 176246 79892 176298 79898
rect 176246 79834 176298 79840
rect 176338 79892 176390 79898
rect 176338 79834 176390 79840
rect 176442 79778 176470 80036
rect 176534 79898 176562 80036
rect 176626 79903 176654 80036
rect 176522 79892 176574 79898
rect 176522 79834 176574 79840
rect 176612 79894 176668 79903
rect 176612 79829 176668 79838
rect 176166 79750 176332 79778
rect 176442 79750 176516 79778
rect 176060 79727 176116 79736
rect 176108 79688 176160 79694
rect 176108 79630 176160 79636
rect 176200 79688 176252 79694
rect 176200 79630 176252 79636
rect 175844 79580 175918 79608
rect 175738 77752 175794 77761
rect 175738 77687 175794 77696
rect 175740 77648 175792 77654
rect 175844 77625 175872 79580
rect 175924 79484 175976 79490
rect 175924 79426 175976 79432
rect 175740 77590 175792 77596
rect 175830 77616 175886 77625
rect 175648 67516 175700 67522
rect 175648 67458 175700 67464
rect 175752 67454 175780 77590
rect 175830 77551 175886 77560
rect 175832 77376 175884 77382
rect 175832 77318 175884 77324
rect 175844 68270 175872 77318
rect 175936 70009 175964 79426
rect 176120 77994 176148 79630
rect 176108 77988 176160 77994
rect 176108 77930 176160 77936
rect 176212 77654 176240 79630
rect 176304 78849 176332 79750
rect 176384 79688 176436 79694
rect 176384 79630 176436 79636
rect 176290 78840 176346 78849
rect 176290 78775 176346 78784
rect 176200 77648 176252 77654
rect 176014 77616 176070 77625
rect 176200 77590 176252 77596
rect 176014 77551 176070 77560
rect 176028 76770 176056 77551
rect 176304 77500 176332 78775
rect 176120 77472 176332 77500
rect 176016 76764 176068 76770
rect 176016 76706 176068 76712
rect 176120 70394 176148 77472
rect 176396 76906 176424 79630
rect 176488 78577 176516 79750
rect 176568 79688 176620 79694
rect 176718 79676 176746 80036
rect 176810 79971 176838 80036
rect 176796 79962 176852 79971
rect 176796 79897 176852 79906
rect 176902 79812 176930 80036
rect 176994 79966 177022 80036
rect 176982 79960 177034 79966
rect 176982 79902 177034 79908
rect 177086 79898 177114 80036
rect 177074 79892 177126 79898
rect 177074 79834 177126 79840
rect 176902 79784 176976 79812
rect 176844 79688 176896 79694
rect 176718 79648 176792 79676
rect 176568 79630 176620 79636
rect 176474 78568 176530 78577
rect 176474 78503 176530 78512
rect 176580 77382 176608 79630
rect 176660 77648 176712 77654
rect 176660 77590 176712 77596
rect 176568 77376 176620 77382
rect 176568 77318 176620 77324
rect 176384 76900 176436 76906
rect 176384 76842 176436 76848
rect 176200 76764 176252 76770
rect 176200 76706 176252 76712
rect 176212 72593 176240 76706
rect 176198 72584 176254 72593
rect 176198 72519 176254 72528
rect 176382 72584 176438 72593
rect 176382 72519 176438 72528
rect 176120 70366 176240 70394
rect 175922 70000 175978 70009
rect 175922 69935 175978 69944
rect 175924 68672 175976 68678
rect 175924 68614 175976 68620
rect 175936 68474 175964 68614
rect 175924 68468 175976 68474
rect 175924 68410 175976 68416
rect 175832 68264 175884 68270
rect 175832 68206 175884 68212
rect 175740 67448 175792 67454
rect 175740 67390 175792 67396
rect 175556 67380 175608 67386
rect 175556 67322 175608 67328
rect 175464 61872 175516 61878
rect 175464 61814 175516 61820
rect 175372 8968 175424 8974
rect 175372 8910 175424 8916
rect 173992 7608 174044 7614
rect 173992 7550 174044 7556
rect 176212 6254 176240 70366
rect 176292 67448 176344 67454
rect 176292 67390 176344 67396
rect 176304 66978 176332 67390
rect 176292 66972 176344 66978
rect 176292 66914 176344 66920
rect 176304 31074 176332 66914
rect 176396 35222 176424 72519
rect 176672 70394 176700 77590
rect 176764 77330 176792 79648
rect 176844 79630 176896 79636
rect 176856 77654 176884 79630
rect 176948 79608 176976 79784
rect 177178 79642 177206 80036
rect 177132 79614 177206 79642
rect 177270 79642 177298 80036
rect 177362 79778 177390 80036
rect 177454 79880 177482 80036
rect 177546 79948 177574 80036
rect 177652 80022 177988 80050
rect 178040 80038 178092 80044
rect 177546 79920 177620 79948
rect 177454 79852 177528 79880
rect 177362 79750 177436 79778
rect 177270 79614 177344 79642
rect 176948 79580 177068 79608
rect 176844 77648 176896 77654
rect 176844 77590 176896 77596
rect 176764 77302 176884 77330
rect 176752 75472 176804 75478
rect 176752 75414 176804 75420
rect 176764 75002 176792 75414
rect 176752 74996 176804 75002
rect 176752 74938 176804 74944
rect 176672 70366 176792 70394
rect 176568 68468 176620 68474
rect 176568 68410 176620 68416
rect 176580 68270 176608 68410
rect 176568 68264 176620 68270
rect 176568 68206 176620 68212
rect 176476 67380 176528 67386
rect 176476 67322 176528 67328
rect 176488 67182 176516 67322
rect 176476 67176 176528 67182
rect 176476 67118 176528 67124
rect 176384 35216 176436 35222
rect 176384 35158 176436 35164
rect 176292 31068 176344 31074
rect 176292 31010 176344 31016
rect 176488 22778 176516 67118
rect 176476 22772 176528 22778
rect 176476 22714 176528 22720
rect 176580 18698 176608 68206
rect 176764 46850 176792 70366
rect 176856 51066 176884 77302
rect 176936 75472 176988 75478
rect 176936 75414 176988 75420
rect 176948 55146 176976 75414
rect 177040 65822 177068 79580
rect 177132 75478 177160 79614
rect 177316 79540 177344 79614
rect 177224 79512 177344 79540
rect 177224 76770 177252 79512
rect 177212 76764 177264 76770
rect 177212 76706 177264 76712
rect 177224 75954 177252 76706
rect 177212 75948 177264 75954
rect 177212 75890 177264 75896
rect 177120 75472 177172 75478
rect 177120 75414 177172 75420
rect 177212 67380 177264 67386
rect 177212 67322 177264 67328
rect 177120 67244 177172 67250
rect 177120 67186 177172 67192
rect 177132 66774 177160 67186
rect 177120 66768 177172 66774
rect 177120 66710 177172 66716
rect 177224 66706 177252 67322
rect 177212 66700 177264 66706
rect 177212 66642 177264 66648
rect 177028 65816 177080 65822
rect 177028 65758 177080 65764
rect 176936 55140 176988 55146
rect 176936 55082 176988 55088
rect 176844 51060 176896 51066
rect 176844 51002 176896 51008
rect 176752 46844 176804 46850
rect 176752 46786 176804 46792
rect 177408 44130 177436 79750
rect 177500 78033 177528 79852
rect 177486 78024 177542 78033
rect 177486 77959 177542 77968
rect 177592 77897 177620 79920
rect 177854 79928 177910 79937
rect 177764 79892 177816 79898
rect 177854 79863 177910 79872
rect 177764 79834 177816 79840
rect 177670 79792 177726 79801
rect 177670 79727 177726 79736
rect 177684 79529 177712 79727
rect 177670 79520 177726 79529
rect 177670 79455 177726 79464
rect 177578 77888 177634 77897
rect 177578 77823 177634 77832
rect 177776 77654 177804 79834
rect 177764 77648 177816 77654
rect 177764 77590 177816 77596
rect 177580 77308 177632 77314
rect 177580 77250 177632 77256
rect 177592 68270 177620 77250
rect 177672 75948 177724 75954
rect 177672 75890 177724 75896
rect 177580 68264 177632 68270
rect 177580 68206 177632 68212
rect 177396 44124 177448 44130
rect 177396 44066 177448 44072
rect 177684 33794 177712 75890
rect 177672 33788 177724 33794
rect 177672 33730 177724 33736
rect 177776 29646 177804 77590
rect 177868 76906 177896 79863
rect 177960 77994 177988 80022
rect 178038 79656 178094 79665
rect 178144 79626 178172 80514
rect 182192 80442 182220 80566
rect 184388 80572 184440 80578
rect 184388 80514 184440 80520
rect 178592 80436 178644 80442
rect 178592 80378 178644 80384
rect 182180 80436 182232 80442
rect 182180 80378 182232 80384
rect 178314 80336 178370 80345
rect 178314 80271 178370 80280
rect 178224 80028 178276 80034
rect 178224 79970 178276 79976
rect 178038 79591 178094 79600
rect 178132 79620 178184 79626
rect 178052 78577 178080 79591
rect 178132 79562 178184 79568
rect 178236 79529 178264 79970
rect 178328 79558 178356 80271
rect 178316 79552 178368 79558
rect 178222 79520 178278 79529
rect 178316 79494 178368 79500
rect 178222 79455 178278 79464
rect 178038 78568 178094 78577
rect 178038 78503 178094 78512
rect 177948 77988 178000 77994
rect 177948 77930 178000 77936
rect 178500 77512 178552 77518
rect 178500 77454 178552 77460
rect 177856 76900 177908 76906
rect 177856 76842 177908 76848
rect 177764 29640 177816 29646
rect 177764 29582 177816 29588
rect 176568 18692 176620 18698
rect 176568 18634 176620 18640
rect 177868 18630 177896 76842
rect 178512 76673 178540 77454
rect 178038 76664 178094 76673
rect 178038 76599 178094 76608
rect 178498 76664 178554 76673
rect 178498 76599 178554 76608
rect 177948 74860 178000 74866
rect 177948 74802 178000 74808
rect 177856 18624 177908 18630
rect 177856 18566 177908 18572
rect 177960 17270 177988 74802
rect 177948 17264 178000 17270
rect 177948 17206 178000 17212
rect 178052 16574 178080 76599
rect 178604 76498 178632 80378
rect 183466 80336 183522 80345
rect 183466 80271 183522 80280
rect 179512 80232 179564 80238
rect 179512 80174 179564 80180
rect 178960 79484 179012 79490
rect 178960 79426 179012 79432
rect 178776 78192 178828 78198
rect 178776 78134 178828 78140
rect 178684 78056 178736 78062
rect 178684 77998 178736 78004
rect 178592 76492 178644 76498
rect 178592 76434 178644 76440
rect 178052 16546 178632 16574
rect 176200 6248 176252 6254
rect 176200 6190 176252 6196
rect 173900 4820 173952 4826
rect 173900 4762 173952 4768
rect 173164 3868 173216 3874
rect 173164 3810 173216 3816
rect 171968 3800 172020 3806
rect 171968 3742 172020 3748
rect 171876 3120 171928 3126
rect 171876 3062 171928 3068
rect 171784 2916 171836 2922
rect 171784 2858 171836 2864
rect 171980 480 172008 3742
rect 173176 480 173204 3810
rect 175464 3528 175516 3534
rect 175464 3470 175516 3476
rect 174268 3120 174320 3126
rect 174268 3062 174320 3068
rect 174280 480 174308 3062
rect 175476 480 175504 3470
rect 176660 3460 176712 3466
rect 176660 3402 176712 3408
rect 176672 480 176700 3402
rect 177856 2916 177908 2922
rect 177856 2858 177908 2864
rect 177868 480 177896 2858
rect 156574 354 156686 480
rect 156156 326 156686 354
rect 156574 -960 156686 326
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 178604 354 178632 16546
rect 178696 3942 178724 77998
rect 178684 3936 178736 3942
rect 178684 3878 178736 3884
rect 178788 3874 178816 78134
rect 178972 78062 179000 79426
rect 179144 79416 179196 79422
rect 179144 79358 179196 79364
rect 179052 79144 179104 79150
rect 179052 79086 179104 79092
rect 179064 78674 179092 79086
rect 179052 78668 179104 78674
rect 179052 78610 179104 78616
rect 179156 78198 179184 79358
rect 179236 78668 179288 78674
rect 179236 78610 179288 78616
rect 179144 78192 179196 78198
rect 179144 78134 179196 78140
rect 178960 78056 179012 78062
rect 178960 77998 179012 78004
rect 179144 77852 179196 77858
rect 179144 77794 179196 77800
rect 179052 77784 179104 77790
rect 179052 77726 179104 77732
rect 178868 77580 178920 77586
rect 178868 77522 178920 77528
rect 178880 69562 178908 77522
rect 179064 73710 179092 77726
rect 179052 73704 179104 73710
rect 179052 73646 179104 73652
rect 178868 69556 178920 69562
rect 178868 69498 178920 69504
rect 178776 3868 178828 3874
rect 178776 3810 178828 3816
rect 179064 3670 179092 73646
rect 179156 6458 179184 77794
rect 179248 76786 179276 78610
rect 179328 78192 179380 78198
rect 179328 78134 179380 78140
rect 179340 77858 179368 78134
rect 179328 77852 179380 77858
rect 179328 77794 179380 77800
rect 179248 76758 179368 76786
rect 179234 76664 179290 76673
rect 179234 76599 179290 76608
rect 179144 6452 179196 6458
rect 179144 6394 179196 6400
rect 179248 3738 179276 76599
rect 179340 3806 179368 76758
rect 179524 64874 179552 80174
rect 180982 79792 181038 79801
rect 180982 79727 181038 79736
rect 180996 79218 181024 79727
rect 180984 79212 181036 79218
rect 180984 79154 181036 79160
rect 183480 78577 183508 80271
rect 183466 78568 183522 78577
rect 183466 78503 183522 78512
rect 180064 78260 180116 78266
rect 180064 78202 180116 78208
rect 179972 77852 180024 77858
rect 179972 77794 180024 77800
rect 179984 75546 180012 77794
rect 180076 75721 180104 78202
rect 181996 77988 182048 77994
rect 181996 77930 182048 77936
rect 180616 77920 180668 77926
rect 180616 77862 180668 77868
rect 180062 75712 180118 75721
rect 180062 75647 180118 75656
rect 179972 75540 180024 75546
rect 179972 75482 180024 75488
rect 180524 73976 180576 73982
rect 180524 73918 180576 73924
rect 180536 73778 180564 73918
rect 180524 73772 180576 73778
rect 180524 73714 180576 73720
rect 179432 64846 179552 64874
rect 179432 16574 179460 64846
rect 179432 16546 180288 16574
rect 179328 3800 179380 3806
rect 179328 3742 179380 3748
rect 179236 3732 179288 3738
rect 179236 3674 179288 3680
rect 179052 3664 179104 3670
rect 179052 3606 179104 3612
rect 180260 480 180288 16546
rect 180536 3466 180564 73714
rect 180628 6390 180656 77862
rect 181444 76628 181496 76634
rect 181444 76570 181496 76576
rect 180800 75608 180852 75614
rect 180800 75550 180852 75556
rect 180708 75540 180760 75546
rect 180708 75482 180760 75488
rect 180720 75041 180748 75482
rect 180706 75032 180762 75041
rect 180706 74967 180762 74976
rect 180616 6384 180668 6390
rect 180616 6326 180668 6332
rect 180720 3534 180748 74967
rect 180812 16574 180840 75550
rect 180812 16546 181024 16574
rect 180708 3528 180760 3534
rect 180708 3470 180760 3476
rect 180524 3460 180576 3466
rect 180524 3402 180576 3408
rect 179022 354 179134 480
rect 178604 326 179134 354
rect 179022 -960 179134 326
rect 180218 -960 180330 480
rect 180996 354 181024 16546
rect 181456 4078 181484 76570
rect 182008 74934 182036 77930
rect 183480 77489 183508 78503
rect 183466 77480 183522 77489
rect 183466 77415 183522 77424
rect 184294 77480 184350 77489
rect 184294 77415 184350 77424
rect 181996 74928 182048 74934
rect 181996 74870 182048 74876
rect 181534 73808 181590 73817
rect 181534 73743 181590 73752
rect 181444 4072 181496 4078
rect 181444 4014 181496 4020
rect 181548 4010 181576 73743
rect 182008 70394 182036 74870
rect 182180 72480 182232 72486
rect 182180 72422 182232 72428
rect 182008 70366 182128 70394
rect 182100 6186 182128 70366
rect 182088 6180 182140 6186
rect 182088 6122 182140 6128
rect 181536 4004 181588 4010
rect 181536 3946 181588 3952
rect 181414 354 181526 480
rect 180996 326 181526 354
rect 182192 354 182220 72422
rect 184204 71120 184256 71126
rect 184204 71062 184256 71068
rect 182822 68368 182878 68377
rect 182822 68303 182878 68312
rect 182836 3398 182864 68303
rect 183560 64184 183612 64190
rect 183560 64126 183612 64132
rect 183572 16574 183600 64126
rect 183572 16546 183784 16574
rect 182824 3392 182876 3398
rect 182824 3334 182876 3340
rect 183756 480 183784 16546
rect 184216 3262 184244 71062
rect 184308 31142 184336 77415
rect 184400 68338 184428 80514
rect 186226 79520 186282 79529
rect 186226 79455 186282 79464
rect 185584 78804 185636 78810
rect 185584 78746 185636 78752
rect 184940 76560 184992 76566
rect 184940 76502 184992 76508
rect 184388 68332 184440 68338
rect 184388 68274 184440 68280
rect 184296 31136 184348 31142
rect 184296 31078 184348 31084
rect 184952 11694 184980 76502
rect 185032 74996 185084 75002
rect 185032 74938 185084 74944
rect 184940 11688 184992 11694
rect 184940 11630 184992 11636
rect 185044 6914 185072 74938
rect 185596 65890 185624 78746
rect 186240 78577 186268 79455
rect 186226 78568 186282 78577
rect 186226 78503 186282 78512
rect 186226 74488 186282 74497
rect 186226 74423 186282 74432
rect 185584 65884 185636 65890
rect 185584 65826 185636 65832
rect 186136 11688 186188 11694
rect 186136 11630 186188 11636
rect 184952 6886 185072 6914
rect 184204 3256 184256 3262
rect 184204 3198 184256 3204
rect 184952 480 184980 6886
rect 186148 480 186176 11630
rect 186240 3602 186268 74423
rect 186608 64802 186636 198902
rect 186700 81462 186728 200194
rect 187056 197940 187108 197946
rect 187056 197882 187108 197888
rect 186780 151632 186832 151638
rect 186780 151574 186832 151580
rect 186688 81456 186740 81462
rect 186688 81398 186740 81404
rect 186688 80912 186740 80918
rect 186688 80854 186740 80860
rect 186700 80646 186728 80854
rect 186688 80640 186740 80646
rect 186688 80582 186740 80588
rect 186792 65754 186820 151574
rect 186964 149048 187016 149054
rect 186964 148990 187016 148996
rect 186872 141976 186924 141982
rect 186872 141918 186924 141924
rect 186884 69494 186912 141918
rect 186976 81530 187004 148990
rect 187068 138145 187096 197882
rect 187424 189644 187476 189650
rect 187424 189586 187476 189592
rect 187240 151496 187292 151502
rect 187240 151438 187292 151444
rect 187148 141976 187200 141982
rect 187148 141918 187200 141924
rect 187160 141778 187188 141918
rect 187148 141772 187200 141778
rect 187148 141714 187200 141720
rect 187148 140276 187200 140282
rect 187148 140218 187200 140224
rect 187054 138136 187110 138145
rect 187054 138071 187110 138080
rect 187054 138000 187110 138009
rect 187054 137935 187110 137944
rect 186964 81524 187016 81530
rect 186964 81466 187016 81472
rect 186964 81116 187016 81122
rect 186964 81058 187016 81064
rect 186976 80714 187004 81058
rect 186964 80708 187016 80714
rect 186964 80650 187016 80656
rect 187068 71194 187096 137935
rect 187160 79490 187188 140218
rect 187252 99521 187280 151438
rect 187332 141636 187384 141642
rect 187332 141578 187384 141584
rect 187344 137193 187372 141578
rect 187436 137873 187464 189586
rect 187514 140584 187570 140593
rect 187514 140519 187570 140528
rect 187528 139505 187556 140519
rect 187514 139496 187570 139505
rect 187514 139431 187570 139440
rect 187422 137864 187478 137873
rect 187422 137799 187478 137808
rect 187330 137184 187386 137193
rect 187330 137119 187386 137128
rect 187238 99512 187294 99521
rect 187238 99447 187294 99456
rect 187238 98696 187294 98705
rect 187238 98631 187294 98640
rect 187148 79484 187200 79490
rect 187148 79426 187200 79432
rect 187252 72758 187280 98631
rect 187424 81524 187476 81530
rect 187424 81466 187476 81472
rect 187332 81116 187384 81122
rect 187332 81058 187384 81064
rect 187344 80578 187372 81058
rect 187332 80572 187384 80578
rect 187332 80514 187384 80520
rect 187436 76362 187464 81466
rect 187516 81456 187568 81462
rect 187516 81398 187568 81404
rect 187528 80850 187556 81398
rect 187516 80844 187568 80850
rect 187516 80786 187568 80792
rect 187528 80510 187556 80786
rect 187712 80782 187740 200262
rect 187884 199776 187936 199782
rect 187884 199718 187936 199724
rect 187792 195424 187844 195430
rect 187792 195366 187844 195372
rect 187700 80776 187752 80782
rect 187700 80718 187752 80724
rect 187516 80504 187568 80510
rect 187516 80446 187568 80452
rect 187606 78568 187662 78577
rect 187606 78503 187662 78512
rect 187424 76356 187476 76362
rect 187424 76298 187476 76304
rect 187240 72752 187292 72758
rect 187240 72694 187292 72700
rect 187056 71188 187108 71194
rect 187056 71130 187108 71136
rect 187620 71097 187648 78503
rect 187700 78124 187752 78130
rect 187700 78066 187752 78072
rect 187712 77761 187740 78066
rect 187698 77752 187754 77761
rect 187698 77687 187754 77696
rect 187712 77314 187740 77687
rect 187700 77308 187752 77314
rect 187700 77250 187752 77256
rect 187700 76492 187752 76498
rect 187700 76434 187752 76440
rect 187712 76265 187740 76434
rect 187698 76256 187754 76265
rect 187698 76191 187754 76200
rect 187700 75336 187752 75342
rect 187700 75278 187752 75284
rect 187606 71088 187662 71097
rect 187606 71023 187662 71032
rect 186872 69488 186924 69494
rect 186872 69430 186924 69436
rect 186780 65748 186832 65754
rect 186780 65690 186832 65696
rect 186596 64796 186648 64802
rect 186596 64738 186648 64744
rect 186608 64394 186636 64738
rect 187146 64560 187202 64569
rect 187146 64495 187202 64504
rect 187160 64462 187188 64495
rect 187148 64456 187200 64462
rect 187148 64398 187200 64404
rect 186596 64388 186648 64394
rect 186596 64330 186648 64336
rect 187160 63578 187188 64398
rect 187148 63572 187200 63578
rect 187148 63514 187200 63520
rect 186320 49224 186372 49230
rect 186320 49166 186372 49172
rect 186332 16574 186360 49166
rect 187712 16574 187740 75278
rect 187804 56273 187832 195366
rect 187896 60489 187924 199718
rect 187988 144498 188016 262375
rect 188160 148912 188212 148918
rect 188160 148854 188212 148860
rect 187976 144492 188028 144498
rect 187976 144434 188028 144440
rect 187976 143472 188028 143478
rect 187976 143414 188028 143420
rect 188068 143472 188120 143478
rect 188068 143414 188120 143420
rect 187988 73817 188016 143414
rect 188080 143138 188108 143414
rect 188068 143132 188120 143138
rect 188068 143074 188120 143080
rect 188068 142656 188120 142662
rect 188068 142598 188120 142604
rect 187974 73808 188030 73817
rect 187974 73743 188030 73752
rect 187988 73545 188016 73743
rect 187974 73536 188030 73545
rect 187974 73471 188030 73480
rect 188080 70854 188108 142598
rect 188172 72622 188200 148854
rect 188264 148617 188292 263638
rect 189092 200802 189120 277374
rect 199396 267034 199424 404330
rect 203536 287706 203564 630634
rect 203524 287700 203576 287706
rect 203524 287642 203576 287648
rect 204720 276684 204772 276690
rect 204720 276626 204772 276632
rect 204732 276078 204760 276626
rect 204444 276072 204496 276078
rect 204444 276014 204496 276020
rect 204720 276072 204772 276078
rect 204720 276014 204772 276020
rect 199384 267028 199436 267034
rect 199384 266970 199436 266976
rect 195980 265532 196032 265538
rect 195980 265474 196032 265480
rect 192116 265464 192168 265470
rect 192116 265406 192168 265412
rect 190644 263764 190696 263770
rect 190644 263706 190696 263712
rect 190000 263492 190052 263498
rect 190000 263434 190052 263440
rect 190012 262614 190040 263434
rect 189264 262608 189316 262614
rect 189264 262550 189316 262556
rect 190000 262608 190052 262614
rect 190000 262550 190052 262556
rect 189276 262313 189304 262550
rect 190460 262404 190512 262410
rect 190460 262346 190512 262352
rect 189262 262304 189318 262313
rect 189172 262268 189224 262274
rect 189262 262239 189318 262248
rect 189172 262210 189224 262216
rect 189080 200796 189132 200802
rect 189080 200738 189132 200744
rect 189184 198762 189212 262210
rect 189816 261588 189868 261594
rect 189816 261530 189868 261536
rect 189540 260568 189592 260574
rect 189540 260510 189592 260516
rect 189264 199164 189316 199170
rect 189264 199106 189316 199112
rect 189172 198756 189224 198762
rect 189172 198698 189224 198704
rect 188344 197600 188396 197606
rect 188344 197542 188396 197548
rect 188250 148608 188306 148617
rect 188250 148543 188306 148552
rect 188252 142996 188304 143002
rect 188252 142938 188304 142944
rect 188264 98705 188292 142938
rect 188356 100881 188384 197542
rect 189172 196920 189224 196926
rect 189172 196862 189224 196868
rect 188528 178084 188580 178090
rect 188528 178026 188580 178032
rect 188436 151836 188488 151842
rect 188436 151778 188488 151784
rect 188448 149025 188476 151778
rect 188434 149016 188490 149025
rect 188434 148951 188490 148960
rect 188436 146056 188488 146062
rect 188436 145998 188488 146004
rect 188448 113174 188476 145998
rect 188540 144294 188568 178026
rect 188712 151564 188764 151570
rect 188712 151506 188764 151512
rect 188620 148980 188672 148986
rect 188620 148922 188672 148928
rect 188528 144288 188580 144294
rect 188528 144230 188580 144236
rect 188632 139262 188660 148922
rect 188724 142662 188752 151506
rect 188712 142656 188764 142662
rect 188712 142598 188764 142604
rect 188620 139256 188672 139262
rect 188620 139198 188672 139204
rect 188448 113146 188936 113174
rect 188342 100872 188398 100881
rect 188342 100807 188398 100816
rect 188618 99512 188674 99521
rect 188618 99447 188674 99456
rect 188342 98832 188398 98841
rect 188342 98767 188398 98776
rect 188250 98696 188306 98705
rect 188250 98631 188306 98640
rect 188356 72690 188384 98767
rect 188526 93800 188582 93809
rect 188526 93735 188582 93744
rect 188540 74390 188568 93735
rect 188528 74384 188580 74390
rect 188528 74326 188580 74332
rect 188540 73982 188568 74326
rect 188528 73976 188580 73982
rect 188528 73918 188580 73924
rect 188344 72684 188396 72690
rect 188344 72626 188396 72632
rect 188160 72616 188212 72622
rect 188160 72558 188212 72564
rect 188632 70922 188660 99447
rect 188908 92546 188936 113146
rect 189078 100872 189134 100881
rect 189078 100807 189134 100816
rect 188988 99408 189040 99414
rect 188988 99350 189040 99356
rect 189000 98841 189028 99350
rect 188986 98832 189042 98841
rect 188986 98767 189042 98776
rect 188896 92540 188948 92546
rect 188896 92482 188948 92488
rect 189092 74186 189120 100807
rect 189080 74180 189132 74186
rect 189080 74122 189132 74128
rect 188620 70916 188672 70922
rect 188620 70858 188672 70864
rect 188068 70848 188120 70854
rect 188068 70790 188120 70796
rect 188434 68912 188490 68921
rect 188434 68847 188490 68856
rect 189078 68912 189134 68921
rect 189078 68847 189134 68856
rect 188448 67726 188476 68847
rect 189092 68406 189120 68847
rect 189080 68400 189132 68406
rect 189080 68342 189132 68348
rect 189092 67794 189120 68342
rect 189080 67788 189132 67794
rect 189080 67730 189132 67736
rect 188436 67720 188488 67726
rect 189184 67674 189212 196862
rect 189276 80714 189304 199106
rect 189448 145852 189500 145858
rect 189448 145794 189500 145800
rect 189356 143540 189408 143546
rect 189356 143482 189408 143488
rect 189264 80708 189316 80714
rect 189264 80650 189316 80656
rect 189264 76832 189316 76838
rect 189264 76774 189316 76780
rect 189276 76634 189304 76774
rect 189264 76628 189316 76634
rect 189264 76570 189316 76576
rect 188436 67662 188488 67668
rect 189092 67646 189212 67674
rect 189092 65958 189120 67646
rect 189080 65952 189132 65958
rect 189080 65894 189132 65900
rect 189092 65618 189120 65894
rect 189080 65612 189132 65618
rect 189080 65554 189132 65560
rect 189080 63436 189132 63442
rect 189080 63378 189132 63384
rect 189092 62898 189120 63378
rect 189080 62892 189132 62898
rect 189080 62834 189132 62840
rect 187882 60480 187938 60489
rect 187882 60415 187938 60424
rect 187790 56264 187846 56273
rect 187790 56199 187846 56208
rect 189368 55078 189396 143482
rect 189460 67046 189488 145794
rect 189552 142730 189580 260510
rect 189724 260160 189776 260166
rect 189724 260102 189776 260108
rect 189632 260092 189684 260098
rect 189632 260034 189684 260040
rect 189644 143041 189672 260034
rect 189736 158438 189764 260102
rect 189828 193186 189856 261530
rect 190090 259856 190146 259865
rect 190090 259791 190146 259800
rect 190000 199232 190052 199238
rect 190000 199174 190052 199180
rect 189816 193180 189868 193186
rect 189816 193122 189868 193128
rect 189816 165640 189868 165646
rect 189816 165582 189868 165588
rect 189724 158432 189776 158438
rect 189724 158374 189776 158380
rect 189828 144226 189856 165582
rect 189906 146976 189962 146985
rect 189906 146911 189962 146920
rect 189816 144220 189868 144226
rect 189816 144162 189868 144168
rect 189630 143032 189686 143041
rect 189630 142967 189686 142976
rect 189540 142724 189592 142730
rect 189540 142666 189592 142672
rect 189816 141228 189868 141234
rect 189816 141170 189868 141176
rect 189632 139528 189684 139534
rect 189632 139470 189684 139476
rect 189644 75138 189672 139470
rect 189724 139256 189776 139262
rect 189724 139198 189776 139204
rect 189736 76634 189764 139198
rect 189828 99414 189856 141170
rect 189920 138718 189948 146911
rect 189908 138712 189960 138718
rect 189908 138654 189960 138660
rect 189816 99408 189868 99414
rect 189816 99350 189868 99356
rect 189724 76628 189776 76634
rect 189724 76570 189776 76576
rect 189632 75132 189684 75138
rect 189632 75074 189684 75080
rect 189724 69692 189776 69698
rect 189724 69634 189776 69640
rect 189448 67040 189500 67046
rect 189448 66982 189500 66988
rect 189356 55072 189408 55078
rect 189356 55014 189408 55020
rect 189368 54534 189396 55014
rect 189356 54528 189408 54534
rect 189356 54470 189408 54476
rect 189736 16574 189764 69634
rect 190012 62898 190040 199174
rect 190104 142769 190132 259791
rect 190182 259720 190238 259729
rect 190182 259655 190238 259664
rect 190090 142760 190146 142769
rect 190090 142695 190146 142704
rect 190196 142089 190224 259655
rect 190472 199510 190500 262346
rect 190552 262336 190604 262342
rect 190552 262278 190604 262284
rect 190460 199504 190512 199510
rect 190460 199446 190512 199452
rect 190564 199442 190592 262278
rect 190552 199436 190604 199442
rect 190552 199378 190604 199384
rect 190552 199096 190604 199102
rect 190552 199038 190604 199044
rect 190460 195492 190512 195498
rect 190460 195434 190512 195440
rect 190276 143404 190328 143410
rect 190276 143346 190328 143352
rect 190182 142080 190238 142089
rect 190182 142015 190238 142024
rect 190288 72554 190316 143346
rect 190368 98252 190420 98258
rect 190368 98194 190420 98200
rect 190276 72548 190328 72554
rect 190276 72490 190328 72496
rect 190000 62892 190052 62898
rect 190000 62834 190052 62840
rect 190380 34513 190408 98194
rect 190472 55214 190500 195434
rect 190564 62014 190592 199038
rect 190656 143206 190684 263706
rect 191012 260228 191064 260234
rect 191012 260170 191064 260176
rect 190920 260092 190972 260098
rect 190920 260034 190972 260040
rect 190826 259992 190882 260001
rect 190826 259927 190882 259936
rect 190736 259480 190788 259486
rect 190736 259422 190788 259428
rect 190644 143200 190696 143206
rect 190644 143142 190696 143148
rect 190748 141409 190776 259422
rect 190840 142905 190868 259927
rect 190932 143070 190960 260034
rect 191024 155854 191052 260170
rect 191930 195664 191986 195673
rect 191930 195599 191986 195608
rect 191012 155848 191064 155854
rect 191012 155790 191064 155796
rect 191012 148572 191064 148578
rect 191012 148514 191064 148520
rect 190920 143064 190972 143070
rect 190920 143006 190972 143012
rect 190826 142896 190882 142905
rect 190826 142831 190882 142840
rect 190734 141400 190790 141409
rect 190734 141335 190790 141344
rect 190644 140480 190696 140486
rect 190644 140422 190696 140428
rect 190552 62008 190604 62014
rect 190552 61950 190604 61956
rect 190460 55208 190512 55214
rect 190460 55150 190512 55156
rect 190656 52329 190684 140422
rect 190828 140412 190880 140418
rect 190828 140354 190880 140360
rect 190736 140344 190788 140350
rect 190736 140286 190788 140292
rect 190748 53689 190776 140286
rect 190840 54641 190868 140354
rect 191024 72962 191052 148514
rect 191104 148300 191156 148306
rect 191104 148242 191156 148248
rect 191116 80442 191144 148242
rect 191196 145648 191248 145654
rect 191196 145590 191248 145596
rect 191104 80436 191156 80442
rect 191104 80378 191156 80384
rect 191208 79626 191236 145590
rect 191380 143472 191432 143478
rect 191380 143414 191432 143420
rect 191286 138952 191342 138961
rect 191286 138887 191342 138896
rect 191196 79620 191248 79626
rect 191196 79562 191248 79568
rect 191300 77858 191328 138887
rect 191288 77852 191340 77858
rect 191288 77794 191340 77800
rect 191392 75070 191420 143414
rect 191840 92540 191892 92546
rect 191840 92482 191892 92488
rect 191748 75336 191800 75342
rect 191748 75278 191800 75284
rect 191760 75070 191788 75278
rect 191380 75064 191432 75070
rect 191380 75006 191432 75012
rect 191748 75064 191800 75070
rect 191748 75006 191800 75012
rect 191012 72956 191064 72962
rect 191012 72898 191064 72904
rect 191852 72826 191880 92482
rect 191840 72820 191892 72826
rect 191840 72762 191892 72768
rect 191748 62008 191800 62014
rect 191748 61950 191800 61956
rect 191760 61606 191788 61950
rect 191748 61600 191800 61606
rect 191748 61542 191800 61548
rect 191944 60058 191972 195599
rect 192024 195356 192076 195362
rect 192024 195298 192076 195304
rect 192036 74534 192064 195298
rect 192128 141574 192156 265406
rect 195244 265192 195296 265198
rect 195244 265134 195296 265140
rect 194876 265056 194928 265062
rect 194876 264998 194928 265004
rect 193588 262812 193640 262818
rect 193588 262754 193640 262760
rect 192484 262744 192536 262750
rect 192484 262686 192536 262692
rect 192208 262676 192260 262682
rect 192208 262618 192260 262624
rect 192220 142118 192248 262618
rect 192392 262540 192444 262546
rect 192392 262482 192444 262488
rect 192300 260364 192352 260370
rect 192300 260306 192352 260312
rect 192208 142112 192260 142118
rect 192208 142054 192260 142060
rect 192312 141846 192340 260306
rect 192404 144430 192432 262482
rect 192496 144566 192524 262686
rect 192668 262472 192720 262478
rect 192668 262414 192720 262420
rect 192576 259956 192628 259962
rect 192576 259898 192628 259904
rect 192484 144560 192536 144566
rect 192484 144502 192536 144508
rect 192392 144424 192444 144430
rect 192392 144366 192444 144372
rect 192588 142254 192616 259898
rect 192680 145382 192708 262414
rect 193496 261384 193548 261390
rect 193496 261326 193548 261332
rect 193312 200388 193364 200394
rect 193312 200330 193364 200336
rect 193220 199300 193272 199306
rect 193220 199242 193272 199248
rect 192758 196616 192814 196625
rect 192758 196551 192814 196560
rect 192668 145376 192720 145382
rect 192668 145318 192720 145324
rect 192668 142792 192720 142798
rect 192668 142734 192720 142740
rect 192576 142248 192628 142254
rect 192576 142190 192628 142196
rect 192300 141840 192352 141846
rect 192300 141782 192352 141788
rect 192116 141568 192168 141574
rect 192116 141510 192168 141516
rect 192392 140684 192444 140690
rect 192392 140626 192444 140632
rect 192300 140616 192352 140622
rect 192300 140558 192352 140564
rect 192036 74506 192156 74534
rect 191944 60030 192064 60058
rect 191930 57216 191986 57225
rect 191930 57151 191986 57160
rect 191748 55208 191800 55214
rect 191748 55150 191800 55156
rect 190826 54632 190882 54641
rect 191760 54602 191788 55150
rect 190826 54567 190882 54576
rect 191748 54596 191800 54602
rect 191748 54538 191800 54544
rect 190734 53680 190790 53689
rect 190734 53615 190790 53624
rect 190642 52320 190698 52329
rect 190642 52255 190698 52264
rect 191746 52320 191802 52329
rect 191746 52255 191802 52264
rect 191760 51921 191788 52255
rect 191746 51912 191802 51921
rect 191746 51847 191802 51856
rect 191944 45554 191972 57151
rect 192036 50697 192064 60030
rect 192128 59294 192156 74506
rect 192312 71738 192340 140558
rect 192300 71732 192352 71738
rect 192300 71674 192352 71680
rect 192404 71602 192432 140626
rect 192576 140140 192628 140146
rect 192576 140082 192628 140088
rect 192482 138816 192538 138825
rect 192482 138751 192538 138760
rect 192496 72894 192524 138751
rect 192588 79558 192616 140082
rect 192680 98258 192708 142734
rect 192668 98252 192720 98258
rect 192668 98194 192720 98200
rect 192576 79552 192628 79558
rect 192576 79494 192628 79500
rect 192484 72888 192536 72894
rect 192484 72830 192536 72836
rect 192496 72690 192524 72830
rect 192484 72684 192536 72690
rect 192484 72626 192536 72632
rect 192392 71596 192444 71602
rect 192392 71538 192444 71544
rect 192116 59288 192168 59294
rect 192116 59230 192168 59236
rect 192772 56545 192800 196551
rect 192852 145988 192904 145994
rect 192852 145930 192904 145936
rect 192864 70990 192892 145930
rect 192944 144152 192996 144158
rect 192944 144094 192996 144100
rect 192956 73846 192984 144094
rect 193128 79280 193180 79286
rect 193128 79222 193180 79228
rect 193140 76838 193168 79222
rect 193128 76832 193180 76838
rect 193128 76774 193180 76780
rect 193126 76528 193182 76537
rect 193126 76463 193182 76472
rect 192944 73840 192996 73846
rect 192944 73782 192996 73788
rect 192852 70984 192904 70990
rect 192852 70926 192904 70932
rect 193036 59288 193088 59294
rect 193036 59230 193088 59236
rect 193048 58750 193076 59230
rect 193036 58744 193088 58750
rect 193036 58686 193088 58692
rect 192758 56536 192814 56545
rect 192758 56471 192814 56480
rect 193034 56536 193090 56545
rect 193034 56471 193090 56480
rect 193048 56137 193076 56471
rect 193034 56128 193090 56137
rect 193034 56063 193090 56072
rect 192022 50688 192078 50697
rect 192022 50623 192078 50632
rect 191852 45526 191972 45554
rect 189998 34504 190054 34513
rect 189998 34439 190054 34448
rect 190366 34504 190422 34513
rect 190366 34439 190422 34448
rect 190012 33833 190040 34439
rect 189998 33824 190054 33833
rect 189998 33759 190054 33768
rect 191852 16574 191880 45526
rect 186332 16546 186912 16574
rect 187712 16546 188568 16574
rect 189736 16546 189856 16574
rect 191852 16546 192064 16574
rect 186228 3596 186280 3602
rect 186228 3538 186280 3544
rect 182518 354 182630 480
rect 182192 326 182630 354
rect 181414 -960 181526 326
rect 182518 -960 182630 326
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 186884 354 186912 16546
rect 188540 480 188568 16546
rect 189828 4146 189856 16546
rect 189816 4140 189868 4146
rect 189816 4082 189868 4088
rect 190828 4072 190880 4078
rect 190828 4014 190880 4020
rect 189724 3256 189776 3262
rect 189724 3198 189776 3204
rect 189736 480 189764 3198
rect 190840 480 190868 4014
rect 192036 480 192064 16546
rect 193140 3330 193168 76463
rect 193232 57934 193260 199242
rect 193324 64598 193352 200330
rect 193404 195696 193456 195702
rect 193404 195638 193456 195644
rect 193312 64592 193364 64598
rect 193312 64534 193364 64540
rect 193324 64258 193352 64534
rect 193312 64252 193364 64258
rect 193312 64194 193364 64200
rect 193416 60654 193444 195638
rect 193508 143342 193536 261326
rect 193600 144634 193628 262754
rect 193680 261656 193732 261662
rect 193680 261598 193732 261604
rect 193588 144628 193640 144634
rect 193588 144570 193640 144576
rect 193692 144362 193720 261598
rect 193772 261316 193824 261322
rect 193772 261258 193824 261264
rect 193784 145450 193812 261258
rect 193864 260296 193916 260302
rect 193864 260238 193916 260244
rect 193876 155174 193904 260238
rect 194600 195832 194652 195838
rect 194600 195774 194652 195780
rect 193864 155168 193916 155174
rect 193864 155110 193916 155116
rect 193956 148164 194008 148170
rect 193956 148106 194008 148112
rect 193864 147008 193916 147014
rect 193864 146950 193916 146956
rect 193772 145444 193824 145450
rect 193772 145386 193824 145392
rect 193680 144356 193732 144362
rect 193680 144298 193732 144304
rect 193496 143336 193548 143342
rect 193496 143278 193548 143284
rect 193770 139360 193826 139369
rect 193770 139295 193826 139304
rect 193678 139224 193734 139233
rect 193678 139159 193734 139168
rect 193692 71466 193720 139159
rect 193784 71670 193812 139295
rect 193876 79082 193904 146950
rect 193968 81705 193996 148106
rect 194140 146260 194192 146266
rect 194140 146202 194192 146208
rect 194046 139088 194102 139097
rect 194046 139023 194102 139032
rect 193954 81696 194010 81705
rect 193954 81631 194010 81640
rect 193864 79076 193916 79082
rect 193864 79018 193916 79024
rect 193864 75268 193916 75274
rect 193864 75210 193916 75216
rect 193772 71664 193824 71670
rect 193772 71606 193824 71612
rect 193680 71460 193732 71466
rect 193680 71402 193732 71408
rect 193404 60648 193456 60654
rect 193404 60590 193456 60596
rect 193220 57928 193272 57934
rect 193220 57870 193272 57876
rect 193310 53136 193366 53145
rect 193310 53071 193366 53080
rect 193218 52456 193274 52465
rect 193218 52391 193220 52400
rect 193272 52391 193274 52400
rect 193220 52362 193272 52368
rect 193324 16574 193352 53071
rect 193324 16546 193812 16574
rect 193784 3482 193812 16546
rect 193876 4078 193904 75210
rect 194060 74254 194088 139023
rect 194048 74248 194100 74254
rect 194048 74190 194100 74196
rect 194152 73098 194180 146202
rect 194232 145920 194284 145926
rect 194232 145862 194284 145868
rect 194140 73092 194192 73098
rect 194140 73034 194192 73040
rect 194152 72554 194180 73034
rect 194140 72548 194192 72554
rect 194140 72490 194192 72496
rect 194244 72418 194272 145862
rect 194508 79484 194560 79490
rect 194508 79426 194560 79432
rect 194520 79082 194548 79426
rect 194508 79076 194560 79082
rect 194508 79018 194560 79024
rect 194232 72412 194284 72418
rect 194232 72354 194284 72360
rect 194612 68542 194640 195774
rect 194692 195764 194744 195770
rect 194692 195706 194744 195712
rect 194704 69834 194732 195706
rect 194784 148844 194836 148850
rect 194784 148786 194836 148792
rect 194692 69828 194744 69834
rect 194692 69770 194744 69776
rect 194796 69630 194824 148786
rect 194888 139670 194916 264998
rect 194968 263084 195020 263090
rect 194968 263026 195020 263032
rect 194980 141914 195008 263026
rect 195060 261180 195112 261186
rect 195060 261122 195112 261128
rect 195072 144838 195100 261122
rect 195152 190188 195204 190194
rect 195152 190130 195204 190136
rect 195060 144832 195112 144838
rect 195060 144774 195112 144780
rect 194968 141908 195020 141914
rect 194968 141850 195020 141856
rect 195060 141364 195112 141370
rect 195060 141306 195112 141312
rect 194968 141296 195020 141302
rect 194968 141238 195020 141244
rect 194876 139664 194928 139670
rect 194876 139606 194928 139612
rect 194980 70106 195008 141238
rect 195072 71534 195100 141306
rect 195164 81122 195192 190130
rect 195256 139913 195284 265134
rect 195520 145784 195572 145790
rect 195520 145726 195572 145732
rect 195336 140548 195388 140554
rect 195336 140490 195388 140496
rect 195242 139904 195298 139913
rect 195242 139839 195298 139848
rect 195244 138712 195296 138718
rect 195244 138654 195296 138660
rect 195152 81116 195204 81122
rect 195152 81058 195204 81064
rect 195256 73166 195284 138654
rect 195348 81841 195376 140490
rect 195426 90400 195482 90409
rect 195426 90335 195482 90344
rect 195334 81832 195390 81841
rect 195334 81767 195390 81776
rect 195244 73160 195296 73166
rect 195244 73102 195296 73108
rect 195256 72486 195284 73102
rect 195244 72480 195296 72486
rect 195244 72422 195296 72428
rect 195060 71528 195112 71534
rect 195060 71470 195112 71476
rect 194968 70100 195020 70106
rect 194968 70042 195020 70048
rect 194784 69624 194836 69630
rect 194784 69566 194836 69572
rect 194600 68536 194652 68542
rect 194600 68478 194652 68484
rect 195060 68536 195112 68542
rect 195060 68478 195112 68484
rect 195072 68338 195100 68478
rect 195060 68332 195112 68338
rect 195060 68274 195112 68280
rect 194508 60648 194560 60654
rect 194508 60590 194560 60596
rect 194520 60110 194548 60590
rect 194508 60104 194560 60110
rect 194508 60046 194560 60052
rect 194508 57928 194560 57934
rect 194508 57870 194560 57876
rect 194520 57254 194548 57870
rect 194508 57248 194560 57254
rect 194508 57190 194560 57196
rect 194508 52420 194560 52426
rect 194508 52362 194560 52368
rect 194520 51202 194548 52362
rect 194508 51196 194560 51202
rect 194508 51138 194560 51144
rect 195440 36689 195468 90335
rect 195532 71262 195560 145726
rect 195992 145518 196020 265474
rect 197636 265396 197688 265402
rect 197636 265338 197688 265344
rect 196624 263152 196676 263158
rect 196624 263094 196676 263100
rect 196440 261112 196492 261118
rect 196440 261054 196492 261060
rect 196348 196852 196400 196858
rect 196348 196794 196400 196800
rect 196254 196752 196310 196761
rect 196254 196687 196310 196696
rect 196070 195800 196126 195809
rect 196070 195735 196126 195744
rect 195980 145512 196032 145518
rect 195980 145454 196032 145460
rect 195520 71256 195572 71262
rect 195520 71198 195572 71204
rect 195978 68232 196034 68241
rect 195978 68167 196034 68176
rect 195426 36680 195482 36689
rect 195426 36615 195482 36624
rect 195992 16574 196020 68167
rect 196084 45257 196112 195735
rect 196162 195528 196218 195537
rect 196162 195463 196218 195472
rect 196176 49609 196204 195463
rect 196268 60874 196296 196687
rect 196360 64818 196388 196794
rect 196452 151814 196480 261054
rect 196452 151786 196572 151814
rect 196440 147620 196492 147626
rect 196440 147562 196492 147568
rect 196452 147529 196480 147562
rect 196438 147520 196494 147529
rect 196438 147455 196494 147464
rect 196544 145874 196572 151786
rect 196452 145846 196572 145874
rect 196452 143274 196480 145846
rect 196532 145716 196584 145722
rect 196532 145658 196584 145664
rect 196440 143268 196492 143274
rect 196440 143210 196492 143216
rect 196544 71398 196572 145658
rect 196636 144702 196664 263094
rect 197084 260976 197136 260982
rect 197084 260918 197136 260924
rect 196716 259616 196768 259622
rect 196716 259558 196768 259564
rect 196728 146198 196756 259558
rect 196992 148436 197044 148442
rect 196992 148378 197044 148384
rect 196716 146192 196768 146198
rect 196716 146134 196768 146140
rect 196898 145616 196954 145625
rect 196898 145551 196954 145560
rect 196808 144900 196860 144906
rect 196808 144842 196860 144848
rect 196624 144696 196676 144702
rect 196624 144638 196676 144644
rect 196624 142044 196676 142050
rect 196624 141986 196676 141992
rect 196532 71392 196584 71398
rect 196532 71334 196584 71340
rect 196636 70242 196664 141986
rect 196716 141976 196768 141982
rect 196716 141918 196768 141924
rect 196624 70236 196676 70242
rect 196624 70178 196676 70184
rect 196728 70174 196756 141918
rect 196820 82113 196848 144842
rect 196806 82104 196862 82113
rect 196806 82039 196862 82048
rect 196716 70168 196768 70174
rect 196716 70110 196768 70116
rect 196360 64790 196572 64818
rect 196268 60846 196480 60874
rect 196256 60580 196308 60586
rect 196256 60522 196308 60528
rect 196268 60042 196296 60522
rect 196256 60036 196308 60042
rect 196256 59978 196308 59984
rect 196256 59356 196308 59362
rect 196256 59298 196308 59304
rect 196268 58682 196296 59298
rect 196256 58676 196308 58682
rect 196256 58618 196308 58624
rect 196256 57860 196308 57866
rect 196256 57802 196308 57808
rect 196268 57361 196296 57802
rect 196254 57352 196310 57361
rect 196254 57287 196310 57296
rect 196268 56642 196296 57287
rect 196256 56636 196308 56642
rect 196256 56578 196308 56584
rect 196254 56400 196310 56409
rect 196452 56386 196480 60846
rect 196544 59362 196572 64790
rect 196912 60042 196940 145551
rect 197004 74118 197032 148378
rect 197096 143177 197124 260918
rect 197360 197192 197412 197198
rect 197360 197134 197412 197140
rect 197450 197160 197506 197169
rect 197082 143168 197138 143177
rect 197082 143103 197138 143112
rect 196992 74112 197044 74118
rect 196992 74054 197044 74060
rect 197372 61946 197400 197134
rect 197450 197095 197506 197104
rect 197360 61940 197412 61946
rect 197360 61882 197412 61888
rect 197372 61470 197400 61882
rect 197360 61464 197412 61470
rect 197360 61406 197412 61412
rect 196900 60036 196952 60042
rect 196900 59978 196952 59984
rect 196532 59356 196584 59362
rect 196532 59298 196584 59304
rect 196310 56358 196480 56386
rect 196254 56335 196310 56344
rect 196268 56001 196296 56335
rect 196254 55992 196310 56001
rect 196254 55927 196310 55936
rect 196162 49600 196218 49609
rect 196162 49535 196218 49544
rect 196714 49600 196770 49609
rect 196714 49535 196770 49544
rect 196728 49065 196756 49535
rect 196714 49056 196770 49065
rect 196714 48991 196770 49000
rect 197464 48113 197492 197095
rect 197544 196988 197596 196994
rect 197544 196930 197596 196936
rect 197556 52358 197584 196930
rect 197648 139738 197676 265338
rect 199200 265328 199252 265334
rect 199200 265270 199252 265276
rect 199108 265260 199160 265266
rect 199108 265202 199160 265208
rect 197728 263628 197780 263634
rect 197728 263570 197780 263576
rect 197740 147422 197768 263570
rect 197912 261248 197964 261254
rect 197912 261190 197964 261196
rect 197820 260908 197872 260914
rect 197820 260850 197872 260856
rect 197728 147416 197780 147422
rect 197728 147358 197780 147364
rect 197832 145586 197860 260850
rect 197924 147286 197952 261190
rect 198004 261044 198056 261050
rect 198004 260986 198056 260992
rect 198016 150074 198044 260986
rect 199016 200456 199068 200462
rect 199016 200398 199068 200404
rect 198830 197296 198886 197305
rect 198830 197231 198886 197240
rect 198464 151428 198516 151434
rect 198464 151370 198516 151376
rect 198004 150068 198056 150074
rect 198004 150010 198056 150016
rect 198372 148776 198424 148782
rect 198372 148718 198424 148724
rect 198280 148708 198332 148714
rect 198280 148650 198332 148656
rect 197912 147280 197964 147286
rect 197912 147222 197964 147228
rect 198096 147144 198148 147150
rect 198096 147086 198148 147092
rect 197820 145580 197872 145586
rect 197820 145522 197872 145528
rect 197912 140208 197964 140214
rect 197912 140150 197964 140156
rect 197820 140072 197872 140078
rect 197820 140014 197872 140020
rect 197636 139732 197688 139738
rect 197636 139674 197688 139680
rect 197636 78464 197688 78470
rect 197636 78406 197688 78412
rect 197648 78130 197676 78406
rect 197636 78124 197688 78130
rect 197636 78066 197688 78072
rect 197832 69018 197860 140014
rect 197924 70038 197952 140150
rect 198108 76702 198136 147086
rect 198188 147076 198240 147082
rect 198188 147018 198240 147024
rect 198200 79218 198228 147018
rect 198188 79212 198240 79218
rect 198188 79154 198240 79160
rect 198096 76696 198148 76702
rect 198096 76638 198148 76644
rect 197912 70032 197964 70038
rect 197912 69974 197964 69980
rect 197820 69012 197872 69018
rect 197820 68954 197872 68960
rect 198292 68610 198320 148650
rect 198280 68604 198332 68610
rect 198280 68546 198332 68552
rect 197636 61668 197688 61674
rect 197636 61610 197688 61616
rect 197544 52352 197596 52358
rect 197544 52294 197596 52300
rect 197450 48104 197506 48113
rect 197450 48039 197506 48048
rect 196070 45248 196126 45257
rect 196070 45183 196126 45192
rect 197648 16574 197676 61610
rect 198384 53786 198412 148718
rect 198476 78130 198504 151370
rect 198740 147552 198792 147558
rect 198740 147494 198792 147500
rect 198752 146849 198780 147494
rect 198738 146840 198794 146849
rect 198738 146775 198794 146784
rect 198740 78396 198792 78402
rect 198740 78338 198792 78344
rect 198464 78124 198516 78130
rect 198464 78066 198516 78072
rect 198752 78062 198780 78338
rect 198740 78056 198792 78062
rect 198740 77998 198792 78004
rect 198740 58948 198792 58954
rect 198740 58890 198792 58896
rect 198372 53780 198424 53786
rect 198372 53722 198424 53728
rect 198384 53242 198412 53722
rect 198372 53236 198424 53242
rect 198372 53178 198424 53184
rect 198096 52352 198148 52358
rect 198096 52294 198148 52300
rect 198108 51746 198136 52294
rect 198096 51740 198148 51746
rect 198096 51682 198148 51688
rect 198462 48104 198518 48113
rect 198462 48039 198518 48048
rect 198476 47841 198504 48039
rect 198462 47832 198518 47841
rect 198462 47767 198518 47776
rect 195992 16546 196848 16574
rect 197648 16546 197952 16574
rect 193864 4072 193916 4078
rect 193864 4014 193916 4020
rect 195612 4072 195664 4078
rect 195612 4014 195664 4020
rect 195704 4072 195756 4078
rect 195704 4014 195756 4020
rect 193784 3454 194456 3482
rect 193220 3392 193272 3398
rect 193220 3334 193272 3340
rect 193128 3324 193180 3330
rect 193128 3266 193180 3272
rect 193232 480 193260 3334
rect 194428 480 194456 3454
rect 195624 480 195652 4014
rect 195716 3330 195744 4014
rect 195704 3324 195756 3330
rect 195704 3266 195756 3272
rect 196820 480 196848 16546
rect 197924 480 197952 16546
rect 187302 354 187414 480
rect 186884 326 187414 354
rect 187302 -960 187414 326
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198752 354 198780 58890
rect 198844 50425 198872 197231
rect 198924 193112 198976 193118
rect 198924 193054 198976 193060
rect 198936 53650 198964 193054
rect 199028 63510 199056 200398
rect 199120 147218 199148 265202
rect 199212 147354 199240 265270
rect 203248 265124 203300 265130
rect 203248 265066 203300 265072
rect 203156 264988 203208 264994
rect 203156 264930 203208 264936
rect 199292 261520 199344 261526
rect 199292 261462 199344 261468
rect 199200 147348 199252 147354
rect 199200 147290 199252 147296
rect 199108 147212 199160 147218
rect 199108 147154 199160 147160
rect 199304 146130 199332 261462
rect 201868 259820 201920 259826
rect 201868 259762 201920 259768
rect 201590 200288 201646 200297
rect 201590 200223 201646 200232
rect 201130 200152 201186 200161
rect 201130 200087 201186 200096
rect 200304 199028 200356 199034
rect 200304 198970 200356 198976
rect 199660 197124 199712 197130
rect 199660 197066 199712 197072
rect 199384 148504 199436 148510
rect 199384 148446 199436 148452
rect 199292 146124 199344 146130
rect 199292 146066 199344 146072
rect 199292 141704 199344 141710
rect 199292 141646 199344 141652
rect 199108 78532 199160 78538
rect 199108 78474 199160 78480
rect 199120 77994 199148 78474
rect 199108 77988 199160 77994
rect 199108 77930 199160 77936
rect 199304 69970 199332 141646
rect 199396 76974 199424 148446
rect 199474 145752 199530 145761
rect 199474 145687 199530 145696
rect 199488 78062 199516 145687
rect 199566 137184 199622 137193
rect 199566 137119 199622 137128
rect 199580 78538 199608 137119
rect 199568 78532 199620 78538
rect 199568 78474 199620 78480
rect 199476 78056 199528 78062
rect 199476 77998 199528 78004
rect 199384 76968 199436 76974
rect 199384 76910 199436 76916
rect 199292 69964 199344 69970
rect 199292 69906 199344 69912
rect 199016 63504 199068 63510
rect 199016 63446 199068 63452
rect 199200 63504 199252 63510
rect 199200 63446 199252 63452
rect 199212 62830 199240 63446
rect 199200 62824 199252 62830
rect 199200 62766 199252 62772
rect 199106 61976 199162 61985
rect 199106 61911 199162 61920
rect 199120 61878 199148 61911
rect 199108 61872 199160 61878
rect 199108 61814 199160 61820
rect 199120 60790 199148 61814
rect 199108 60784 199160 60790
rect 199108 60726 199160 60732
rect 199672 57497 199700 197066
rect 200210 197024 200266 197033
rect 200210 196959 200266 196968
rect 199844 148640 199896 148646
rect 199844 148582 199896 148588
rect 199750 146296 199806 146305
rect 199750 146231 199806 146240
rect 199764 137329 199792 146231
rect 199750 137320 199806 137329
rect 199750 137255 199806 137264
rect 199856 68678 199884 148582
rect 199936 148232 199988 148238
rect 199936 148174 199988 148180
rect 199844 68672 199896 68678
rect 199844 68614 199896 68620
rect 199948 64734 199976 148174
rect 200120 71052 200172 71058
rect 200120 70994 200172 71000
rect 199936 64728 199988 64734
rect 199936 64670 199988 64676
rect 199658 57488 199714 57497
rect 199658 57423 199714 57432
rect 198924 53644 198976 53650
rect 198924 53586 198976 53592
rect 199108 53644 199160 53650
rect 199108 53586 199160 53592
rect 199120 53174 199148 53586
rect 199108 53168 199160 53174
rect 199108 53110 199160 53116
rect 198830 50416 198886 50425
rect 198830 50351 198886 50360
rect 200132 16574 200160 70994
rect 200224 55185 200252 196959
rect 200316 66026 200344 198970
rect 200396 187604 200448 187610
rect 200396 187546 200448 187552
rect 200304 66020 200356 66026
rect 200304 65962 200356 65968
rect 200408 64666 200436 187546
rect 200764 155644 200816 155650
rect 200764 155586 200816 155592
rect 200672 155576 200724 155582
rect 200672 155518 200724 155524
rect 200580 152584 200632 152590
rect 200580 152526 200632 152532
rect 200486 148336 200542 148345
rect 200486 148271 200542 148280
rect 200396 64660 200448 64666
rect 200396 64602 200448 64608
rect 200210 55176 200266 55185
rect 200210 55111 200266 55120
rect 200500 44033 200528 148271
rect 200592 68814 200620 152526
rect 200684 71330 200712 155518
rect 200776 75886 200804 155586
rect 200946 151192 201002 151201
rect 200946 151127 201002 151136
rect 200854 138680 200910 138689
rect 200854 138615 200910 138624
rect 200764 75880 200816 75886
rect 200764 75822 200816 75828
rect 200672 71324 200724 71330
rect 200672 71266 200724 71272
rect 200762 68912 200818 68921
rect 200762 68847 200818 68856
rect 200580 68808 200632 68814
rect 200580 68750 200632 68756
rect 200776 68270 200804 68847
rect 200764 68264 200816 68270
rect 200764 68206 200816 68212
rect 200868 64870 200896 138615
rect 200960 78674 200988 151127
rect 200948 78668 201000 78674
rect 200948 78610 201000 78616
rect 201144 69698 201172 200087
rect 201500 191412 201552 191418
rect 201500 191354 201552 191360
rect 201222 81424 201278 81433
rect 201222 81359 201278 81368
rect 201236 80102 201264 81359
rect 201224 80096 201276 80102
rect 201224 80038 201276 80044
rect 201512 73710 201540 191354
rect 201500 73704 201552 73710
rect 201500 73646 201552 73652
rect 201132 69692 201184 69698
rect 201132 69634 201184 69640
rect 201408 68264 201460 68270
rect 201408 68206 201460 68212
rect 201420 67658 201448 68206
rect 201408 67652 201460 67658
rect 201408 67594 201460 67600
rect 201408 66020 201460 66026
rect 201408 65962 201460 65968
rect 201420 65550 201448 65962
rect 201408 65544 201460 65550
rect 201408 65486 201460 65492
rect 200856 64864 200908 64870
rect 200856 64806 200908 64812
rect 201604 56574 201632 200223
rect 201684 197056 201736 197062
rect 201684 196998 201736 197004
rect 201696 79014 201724 196998
rect 201776 191344 201828 191350
rect 201776 191286 201828 191292
rect 201684 79008 201736 79014
rect 201684 78950 201736 78956
rect 201788 77926 201816 191286
rect 201880 155922 201908 259762
rect 201960 259548 202012 259554
rect 201960 259490 202012 259496
rect 201972 158370 202000 259490
rect 203064 194132 203116 194138
rect 203064 194074 203116 194080
rect 202878 192808 202934 192817
rect 202878 192743 202934 192752
rect 201960 158364 202012 158370
rect 201960 158306 202012 158312
rect 201868 155916 201920 155922
rect 201868 155858 201920 155864
rect 201868 155780 201920 155786
rect 201868 155722 201920 155728
rect 201776 77920 201828 77926
rect 201776 77862 201828 77868
rect 201684 75200 201736 75206
rect 201684 75142 201736 75148
rect 201592 56568 201644 56574
rect 201592 56510 201644 56516
rect 201406 55176 201462 55185
rect 201406 55111 201462 55120
rect 201420 54505 201448 55111
rect 201406 54496 201462 54505
rect 201406 54431 201462 54440
rect 201592 49088 201644 49094
rect 201592 49030 201644 49036
rect 200486 44024 200542 44033
rect 200486 43959 200542 43968
rect 201406 44024 201462 44033
rect 201406 43959 201462 43968
rect 201420 43625 201448 43959
rect 201406 43616 201462 43625
rect 201406 43551 201462 43560
rect 200132 16546 200344 16574
rect 200316 480 200344 16546
rect 201604 6914 201632 49030
rect 201696 16574 201724 75142
rect 201880 49706 201908 155722
rect 202236 155712 202288 155718
rect 202236 155654 202288 155660
rect 202144 155508 202196 155514
rect 202144 155450 202196 155456
rect 202050 148472 202106 148481
rect 202050 148407 202106 148416
rect 201958 136096 202014 136105
rect 201958 136031 202014 136040
rect 201972 55214 202000 136031
rect 202064 62082 202092 148407
rect 202156 68882 202184 155450
rect 202248 68950 202276 155654
rect 202328 155236 202380 155242
rect 202328 155178 202380 155184
rect 202340 74322 202368 155178
rect 202328 74316 202380 74322
rect 202328 74258 202380 74264
rect 202236 68944 202288 68950
rect 202236 68886 202288 68892
rect 202144 68876 202196 68882
rect 202144 68818 202196 68824
rect 202892 64530 202920 192743
rect 202972 191276 203024 191282
rect 202972 191218 203024 191224
rect 202984 78441 203012 191218
rect 203076 81977 203104 194074
rect 203168 158234 203196 264930
rect 203260 158302 203288 265066
rect 203616 195628 203668 195634
rect 203616 195570 203668 195576
rect 203248 158296 203300 158302
rect 203248 158238 203300 158244
rect 203156 158228 203208 158234
rect 203156 158170 203208 158176
rect 203246 155680 203302 155689
rect 203246 155615 203302 155624
rect 203154 155544 203210 155553
rect 203154 155479 203210 155488
rect 203062 81968 203118 81977
rect 203062 81903 203118 81912
rect 202970 78432 203026 78441
rect 202970 78367 203026 78376
rect 202880 64524 202932 64530
rect 202880 64466 202932 64472
rect 202892 64190 202920 64466
rect 202880 64184 202932 64190
rect 202880 64126 202932 64132
rect 202052 62076 202104 62082
rect 202052 62018 202104 62024
rect 202788 62076 202840 62082
rect 202788 62018 202840 62024
rect 202800 61402 202828 62018
rect 202788 61396 202840 61402
rect 202788 61338 202840 61344
rect 202788 56568 202840 56574
rect 202788 56510 202840 56516
rect 202800 55894 202828 56510
rect 202788 55888 202840 55894
rect 202788 55830 202840 55836
rect 201972 55186 202092 55214
rect 201958 52456 202014 52465
rect 201958 52391 202014 52400
rect 201972 52290 202000 52391
rect 201960 52284 202012 52290
rect 201960 52226 202012 52232
rect 201868 49700 201920 49706
rect 201868 49642 201920 49648
rect 202064 46345 202092 55186
rect 202788 52284 202840 52290
rect 202788 52226 202840 52232
rect 202800 51134 202828 52226
rect 202788 51128 202840 51134
rect 202788 51070 202840 51076
rect 202788 49700 202840 49706
rect 202788 49642 202840 49648
rect 202800 49094 202828 49642
rect 202788 49088 202840 49094
rect 202788 49030 202840 49036
rect 203168 47977 203196 155479
rect 203260 57633 203288 155615
rect 203432 155372 203484 155378
rect 203432 155314 203484 155320
rect 203338 155272 203394 155281
rect 203338 155207 203394 155216
rect 203352 68746 203380 155207
rect 203444 73137 203472 155314
rect 203524 155304 203576 155310
rect 203524 155246 203576 155252
rect 203536 78334 203564 155246
rect 203628 149161 203656 195570
rect 203708 195560 203760 195566
rect 203708 195502 203760 195508
rect 203614 149152 203670 149161
rect 203614 149087 203670 149096
rect 203616 149048 203668 149054
rect 203616 148990 203668 148996
rect 203524 78328 203576 78334
rect 203524 78270 203576 78276
rect 203628 73914 203656 148990
rect 203720 136649 203748 195502
rect 204352 192024 204404 192030
rect 204352 191966 204404 191972
rect 204258 187096 204314 187105
rect 204258 187031 204314 187040
rect 203800 150000 203852 150006
rect 203800 149942 203852 149948
rect 203812 149054 203840 149942
rect 203800 149048 203852 149054
rect 203800 148990 203852 148996
rect 203706 136640 203762 136649
rect 203706 136575 203762 136584
rect 203706 135960 203762 135969
rect 203706 135895 203762 135904
rect 203720 78169 203748 135895
rect 203706 78160 203762 78169
rect 203706 78095 203762 78104
rect 203616 73908 203668 73914
rect 203616 73850 203668 73856
rect 203430 73128 203486 73137
rect 203430 73063 203486 73072
rect 203340 68740 203392 68746
rect 203340 68682 203392 68688
rect 203524 66904 203576 66910
rect 203524 66846 203576 66852
rect 203246 57624 203302 57633
rect 203246 57559 203302 57568
rect 203340 55140 203392 55146
rect 203340 55082 203392 55088
rect 203352 54777 203380 55082
rect 203338 54768 203394 54777
rect 203338 54703 203394 54712
rect 203154 47968 203210 47977
rect 203154 47903 203210 47912
rect 202050 46336 202106 46345
rect 202050 46271 202106 46280
rect 201696 16546 202736 16574
rect 201512 6886 201632 6914
rect 201512 480 201540 6886
rect 202708 480 202736 16546
rect 203536 2990 203564 66846
rect 203614 66056 203670 66065
rect 203614 65991 203670 66000
rect 203628 65822 203656 65991
rect 203616 65816 203668 65822
rect 203616 65758 203668 65764
rect 204168 65816 204220 65822
rect 204168 65758 204220 65764
rect 204180 64938 204208 65758
rect 204168 64932 204220 64938
rect 204168 64874 204220 64880
rect 204166 57624 204222 57633
rect 204166 57559 204222 57568
rect 204180 57361 204208 57559
rect 204166 57352 204222 57361
rect 204166 57287 204222 57296
rect 203982 54768 204038 54777
rect 203982 54703 204038 54712
rect 203996 53854 204024 54703
rect 203984 53848 204036 53854
rect 203984 53790 204036 53796
rect 204166 47968 204222 47977
rect 204166 47903 204222 47912
rect 204180 47705 204208 47903
rect 204166 47696 204222 47705
rect 204166 47631 204222 47640
rect 204272 35873 204300 187031
rect 204364 66201 204392 191966
rect 204456 151230 204484 276014
rect 218072 262886 218100 703582
rect 218808 703474 218836 703582
rect 218950 703520 219062 704960
rect 234632 703582 235028 703610
rect 218992 703474 219020 703520
rect 218808 703446 219020 703474
rect 234632 278050 234660 703582
rect 235000 703474 235028 703582
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 267660 700670 267688 703520
rect 283852 702434 283880 703520
rect 282932 702406 283880 702434
rect 267648 700664 267700 700670
rect 267648 700606 267700 700612
rect 234620 278044 234672 278050
rect 234620 277986 234672 277992
rect 282932 263498 282960 702406
rect 299492 276690 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 332520 700466 332548 703520
rect 348804 702434 348832 703520
rect 364996 702434 365024 703520
rect 347792 702406 348832 702434
rect 364352 702406 365024 702434
rect 332508 700460 332560 700466
rect 332508 700402 332560 700408
rect 299480 276684 299532 276690
rect 299480 276626 299532 276632
rect 282920 263492 282972 263498
rect 282920 263434 282972 263440
rect 347792 262993 347820 702406
rect 364352 275233 364380 702406
rect 397472 699718 397500 703520
rect 413664 700398 413692 703520
rect 413652 700392 413704 700398
rect 413652 700334 413704 700340
rect 429856 699718 429884 703520
rect 396724 699712 396776 699718
rect 396724 699654 396776 699660
rect 397460 699712 397512 699718
rect 397460 699654 397512 699660
rect 428464 699712 428516 699718
rect 428464 699654 428516 699660
rect 429844 699712 429896 699718
rect 429844 699654 429896 699660
rect 396736 284986 396764 699654
rect 396724 284980 396776 284986
rect 396724 284922 396776 284928
rect 364338 275224 364394 275233
rect 364338 275159 364394 275168
rect 428476 273970 428504 699654
rect 462332 660346 462360 703520
rect 478524 702434 478552 703520
rect 477512 702406 478552 702434
rect 462320 660340 462372 660346
rect 462320 660282 462372 660288
rect 428464 273964 428516 273970
rect 428464 273906 428516 273912
rect 347778 262984 347834 262993
rect 347778 262919 347834 262928
rect 218060 262880 218112 262886
rect 477512 262857 477540 702406
rect 494072 271182 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 527192 283626 527220 703520
rect 543476 700330 543504 703520
rect 559668 700330 559696 703520
rect 543464 700324 543516 700330
rect 543464 700266 543516 700272
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 543004 700256 543056 700262
rect 543004 700198 543056 700204
rect 527180 283620 527232 283626
rect 527180 283562 527232 283568
rect 494060 271176 494112 271182
rect 494060 271118 494112 271124
rect 543016 269822 543044 700198
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 579802 564360 579858 564369
rect 579802 564295 579858 564304
rect 579816 563106 579844 564295
rect 579804 563100 579856 563106
rect 579804 563042 579856 563048
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580184 430642 580212 431559
rect 580172 430636 580224 430642
rect 580172 430578 580224 430584
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580184 418198 580212 418231
rect 580172 418192 580224 418198
rect 580172 418134 580224 418140
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 580262 365120 580318 365129
rect 580262 365055 580318 365064
rect 580172 351960 580224 351966
rect 580170 351928 580172 351937
rect 580224 351928 580226 351937
rect 580170 351863 580226 351872
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580184 324358 580212 325207
rect 580172 324352 580224 324358
rect 580172 324294 580224 324300
rect 579986 312080 580042 312089
rect 579986 312015 580042 312024
rect 580000 311914 580028 312015
rect 579988 311908 580040 311914
rect 579988 311850 580040 311856
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580184 298178 580212 298687
rect 580172 298172 580224 298178
rect 580172 298114 580224 298120
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580184 271930 580212 272167
rect 580172 271924 580224 271930
rect 580172 271866 580224 271872
rect 543004 269816 543056 269822
rect 543004 269758 543056 269764
rect 580276 263566 580304 365055
rect 580264 263560 580316 263566
rect 580264 263502 580316 263508
rect 580356 263016 580408 263022
rect 580356 262958 580408 262964
rect 218060 262822 218112 262828
rect 477498 262848 477554 262857
rect 477498 262783 477554 262792
rect 471244 261452 471296 261458
rect 471244 261394 471296 261400
rect 471256 206990 471284 261394
rect 485044 260432 485096 260438
rect 485044 260374 485096 260380
rect 485056 245614 485084 260374
rect 580172 259412 580224 259418
rect 580172 259354 580224 259360
rect 580184 258913 580212 259354
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 485044 245608 485096 245614
rect 580172 245608 580224 245614
rect 485044 245550 485096 245556
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 580368 219065 580396 262958
rect 580448 262948 580500 262954
rect 580448 262890 580500 262896
rect 580460 232393 580488 262890
rect 580446 232384 580502 232393
rect 580446 232319 580502 232328
rect 580354 219056 580410 219065
rect 580354 218991 580410 219000
rect 471244 206984 471296 206990
rect 471244 206926 471296 206932
rect 579804 206984 579856 206990
rect 579804 206926 579856 206932
rect 579816 205737 579844 206926
rect 579802 205728 579858 205737
rect 579802 205663 579858 205672
rect 208674 200424 208730 200433
rect 208674 200359 208730 200368
rect 204626 199336 204682 199345
rect 204626 199271 204682 199280
rect 204536 192908 204588 192914
rect 204536 192850 204588 192856
rect 204444 151224 204496 151230
rect 204444 151166 204496 151172
rect 204442 150240 204498 150249
rect 204442 150175 204498 150184
rect 204350 66192 204406 66201
rect 204350 66127 204406 66136
rect 204456 49473 204484 150175
rect 204548 73001 204576 192850
rect 204640 79150 204668 199271
rect 208582 194440 208638 194449
rect 208582 194375 208638 194384
rect 208490 194304 208546 194313
rect 208490 194239 208546 194248
rect 207296 194200 207348 194206
rect 207202 194168 207258 194177
rect 207296 194142 207348 194148
rect 207202 194103 207258 194112
rect 204720 193044 204772 193050
rect 204720 192986 204772 192992
rect 204628 79144 204680 79150
rect 204628 79086 204680 79092
rect 204732 75682 204760 192986
rect 205916 192976 205968 192982
rect 205916 192918 205968 192924
rect 204904 192704 204956 192710
rect 204904 192646 204956 192652
rect 204812 191888 204864 191894
rect 204812 191830 204864 191836
rect 204824 78418 204852 191830
rect 204916 78946 204944 192646
rect 205732 192092 205784 192098
rect 205732 192034 205784 192040
rect 205638 191040 205694 191049
rect 205638 190975 205694 190984
rect 204996 151360 205048 151366
rect 204996 151302 205048 151308
rect 204904 78940 204956 78946
rect 204904 78882 204956 78888
rect 204824 78390 204944 78418
rect 204916 75818 204944 78390
rect 204904 75812 204956 75818
rect 204904 75754 204956 75760
rect 204720 75676 204772 75682
rect 204720 75618 204772 75624
rect 204916 75274 204944 75754
rect 204904 75268 204956 75274
rect 204904 75210 204956 75216
rect 204534 72992 204590 73001
rect 204534 72927 204590 72936
rect 205008 70310 205036 151302
rect 205088 149728 205140 149734
rect 205088 149670 205140 149676
rect 205100 71641 205128 149670
rect 205086 71632 205142 71641
rect 205086 71567 205142 71576
rect 205100 71233 205128 71567
rect 205086 71224 205142 71233
rect 205086 71159 205142 71168
rect 204996 70304 205048 70310
rect 204996 70246 205048 70252
rect 204718 66192 204774 66201
rect 204718 66127 204774 66136
rect 204732 65521 204760 66127
rect 204718 65512 204774 65521
rect 204718 65447 204774 65456
rect 204442 49464 204498 49473
rect 204442 49399 204498 49408
rect 204718 49464 204774 49473
rect 204718 49399 204774 49408
rect 204732 48929 204760 49399
rect 204718 48920 204774 48929
rect 204718 48855 204774 48864
rect 204352 41064 204404 41070
rect 204352 41006 204404 41012
rect 204258 35864 204314 35873
rect 204258 35799 204314 35808
rect 204272 35193 204300 35799
rect 204258 35184 204314 35193
rect 204258 35119 204314 35128
rect 204364 16574 204392 41006
rect 205652 26217 205680 190975
rect 205744 55865 205772 192034
rect 205824 190052 205876 190058
rect 205824 189994 205876 190000
rect 205836 66094 205864 189994
rect 205928 70281 205956 192918
rect 206008 192840 206060 192846
rect 206008 192782 206060 192788
rect 205914 70272 205970 70281
rect 205914 70207 205970 70216
rect 206020 70145 206048 192782
rect 206100 191956 206152 191962
rect 206100 191898 206152 191904
rect 206112 79098 206140 191898
rect 206190 190088 206246 190097
rect 206190 190023 206246 190032
rect 206204 79218 206232 190023
rect 207020 187468 207072 187474
rect 207020 187410 207072 187416
rect 206468 149932 206520 149938
rect 206468 149874 206520 149880
rect 206284 149864 206336 149870
rect 206284 149806 206336 149812
rect 206192 79212 206244 79218
rect 206192 79154 206244 79160
rect 206112 79070 206232 79098
rect 206204 75449 206232 79070
rect 206190 75440 206246 75449
rect 206190 75375 206246 75384
rect 206296 72865 206324 149806
rect 206376 149796 206428 149802
rect 206376 149738 206428 149744
rect 206388 74050 206416 149738
rect 206480 78849 206508 149874
rect 206650 80064 206706 80073
rect 206650 79999 206706 80008
rect 206560 79212 206612 79218
rect 206560 79154 206612 79160
rect 206466 78840 206522 78849
rect 206466 78775 206522 78784
rect 206572 75721 206600 79154
rect 206664 76770 206692 79999
rect 206652 76764 206704 76770
rect 206652 76706 206704 76712
rect 206558 75712 206614 75721
rect 206558 75647 206614 75656
rect 206926 75712 206982 75721
rect 206926 75647 206982 75656
rect 206940 75313 206968 75647
rect 206926 75304 206982 75313
rect 206926 75239 206982 75248
rect 206376 74044 206428 74050
rect 206376 73986 206428 73992
rect 206282 72856 206338 72865
rect 206282 72791 206338 72800
rect 206006 70136 206062 70145
rect 206006 70071 206062 70080
rect 205824 66088 205876 66094
rect 205824 66030 205876 66036
rect 205730 55856 205786 55865
rect 205730 55791 205786 55800
rect 205732 32700 205784 32706
rect 205732 32642 205784 32648
rect 205638 26208 205694 26217
rect 205638 26143 205694 26152
rect 205652 25537 205680 26143
rect 205638 25528 205694 25537
rect 205638 25463 205694 25472
rect 205744 16574 205772 32642
rect 207032 21865 207060 187410
rect 207112 187400 207164 187406
rect 207112 187342 207164 187348
rect 207018 21856 207074 21865
rect 207018 21791 207074 21800
rect 207124 21321 207152 187342
rect 207216 53718 207244 194103
rect 207308 67250 207336 194142
rect 207572 193996 207624 194002
rect 207572 193938 207624 193944
rect 207480 190256 207532 190262
rect 207480 190198 207532 190204
rect 207388 189712 207440 189718
rect 207388 189654 207440 189660
rect 207296 67244 207348 67250
rect 207296 67186 207348 67192
rect 207400 66842 207428 189654
rect 207492 67386 207520 190198
rect 207584 75750 207612 193938
rect 207664 193928 207716 193934
rect 207664 193870 207716 193876
rect 207676 75857 207704 193870
rect 207848 151292 207900 151298
rect 207848 151234 207900 151240
rect 207756 150408 207808 150414
rect 207754 150376 207756 150385
rect 207808 150376 207810 150385
rect 207754 150311 207810 150320
rect 207860 150226 207888 151234
rect 207768 150198 207888 150226
rect 207768 79422 207796 150198
rect 207848 142860 207900 142866
rect 207848 142802 207900 142808
rect 207756 79416 207808 79422
rect 207756 79358 207808 79364
rect 207860 77722 207888 142802
rect 207848 77716 207900 77722
rect 207848 77658 207900 77664
rect 207662 75848 207718 75857
rect 207662 75783 207718 75792
rect 207572 75744 207624 75750
rect 207572 75686 207624 75692
rect 207860 70394 207888 77658
rect 208214 75848 208270 75857
rect 208214 75783 208270 75792
rect 208228 75177 208256 75783
rect 208308 75744 208360 75750
rect 208308 75686 208360 75692
rect 208320 75206 208348 75686
rect 208308 75200 208360 75206
rect 208214 75168 208270 75177
rect 208308 75142 208360 75148
rect 208214 75103 208270 75112
rect 207768 70366 207888 70394
rect 207480 67380 207532 67386
rect 207480 67322 207532 67328
rect 207388 66836 207440 66842
rect 207388 66778 207440 66784
rect 207204 53712 207256 53718
rect 207204 53654 207256 53660
rect 207216 53106 207244 53654
rect 207204 53100 207256 53106
rect 207204 53042 207256 53048
rect 207204 51060 207256 51066
rect 207204 51002 207256 51008
rect 207216 50969 207244 51002
rect 207202 50960 207258 50969
rect 207202 50895 207258 50904
rect 207216 49774 207244 50895
rect 207204 49768 207256 49774
rect 207204 49710 207256 49716
rect 207204 46844 207256 46850
rect 207204 46786 207256 46792
rect 207216 46753 207244 46786
rect 207202 46744 207258 46753
rect 207202 46679 207258 46688
rect 207110 21312 207166 21321
rect 207110 21247 207166 21256
rect 204364 16546 205128 16574
rect 205744 16546 206232 16574
rect 203892 4140 203944 4146
rect 203892 4082 203944 4088
rect 203524 2984 203576 2990
rect 203524 2926 203576 2932
rect 203904 480 203932 4082
rect 205100 480 205128 16546
rect 206204 480 206232 16546
rect 207768 3330 207796 70366
rect 208400 47728 208452 47734
rect 208400 47670 208452 47676
rect 207938 45656 207994 45665
rect 207938 45591 207940 45600
rect 207992 45591 207994 45600
rect 207940 45562 207992 45568
rect 208412 16574 208440 47670
rect 208504 45529 208532 194239
rect 208596 52193 208624 194375
rect 208688 70009 208716 200359
rect 213920 200184 213972 200190
rect 213920 200126 213972 200132
rect 211344 198620 211396 198626
rect 211344 198562 211396 198568
rect 208860 198484 208912 198490
rect 208860 198426 208912 198432
rect 208768 194064 208820 194070
rect 208768 194006 208820 194012
rect 208674 70000 208730 70009
rect 208674 69935 208730 69944
rect 208780 67318 208808 194006
rect 208872 73778 208900 198426
rect 209870 198248 209926 198257
rect 209870 198183 209926 198192
rect 209780 192568 209832 192574
rect 209318 192536 209374 192545
rect 209780 192510 209832 192516
rect 209318 192471 209374 192480
rect 208952 190120 209004 190126
rect 208952 190062 209004 190068
rect 208860 73772 208912 73778
rect 208860 73714 208912 73720
rect 208964 67454 208992 190062
rect 209044 187536 209096 187542
rect 209044 187478 209096 187484
rect 208952 67448 209004 67454
rect 208952 67390 209004 67396
rect 208768 67312 208820 67318
rect 208768 67254 208820 67260
rect 209056 66162 209084 187478
rect 209136 151156 209188 151162
rect 209136 151098 209188 151104
rect 209148 76537 209176 151098
rect 209228 142928 209280 142934
rect 209228 142870 209280 142876
rect 209240 78810 209268 142870
rect 209228 78804 209280 78810
rect 209228 78746 209280 78752
rect 209240 77353 209268 78746
rect 209226 77344 209282 77353
rect 209226 77279 209282 77288
rect 209134 76528 209190 76537
rect 209134 76463 209190 76472
rect 209044 66156 209096 66162
rect 209044 66098 209096 66104
rect 208582 52184 208638 52193
rect 208582 52119 208638 52128
rect 208766 52184 208822 52193
rect 208766 52119 208822 52128
rect 208780 51785 208808 52119
rect 208766 51776 208822 51785
rect 208766 51711 208822 51720
rect 208490 45520 208546 45529
rect 208490 45455 208546 45464
rect 208504 44849 208532 45455
rect 208490 44840 208546 44849
rect 208490 44775 208546 44784
rect 209332 44169 209360 192471
rect 209318 44160 209374 44169
rect 209318 44095 209374 44104
rect 209792 17921 209820 192510
rect 209884 48249 209912 198183
rect 209964 194268 210016 194274
rect 209964 194210 210016 194216
rect 209976 66978 210004 194210
rect 210332 192636 210384 192642
rect 210332 192578 210384 192584
rect 210056 190324 210108 190330
rect 210056 190266 210108 190272
rect 210068 67182 210096 190266
rect 210238 189816 210294 189825
rect 210238 189751 210294 189760
rect 210148 187332 210200 187338
rect 210148 187274 210200 187280
rect 210056 67176 210108 67182
rect 210056 67118 210108 67124
rect 209964 66972 210016 66978
rect 209964 66914 210016 66920
rect 210160 66230 210188 187274
rect 210252 70394 210280 189751
rect 210344 73030 210372 192578
rect 211160 192500 211212 192506
rect 211160 192442 211212 192448
rect 210424 190460 210476 190466
rect 210424 190402 210476 190408
rect 210436 76906 210464 190402
rect 210516 152720 210568 152726
rect 210516 152662 210568 152668
rect 210528 84130 210556 152662
rect 210608 152652 210660 152658
rect 210608 152594 210660 152600
rect 210620 93854 210648 152594
rect 210620 93826 210832 93854
rect 210528 84102 210740 84130
rect 210514 77208 210570 77217
rect 210514 77143 210570 77152
rect 210528 77042 210556 77143
rect 210516 77036 210568 77042
rect 210516 76978 210568 76984
rect 210424 76900 210476 76906
rect 210424 76842 210476 76848
rect 210528 75954 210556 76978
rect 210516 75948 210568 75954
rect 210516 75890 210568 75896
rect 210332 73024 210384 73030
rect 210332 72966 210384 72972
rect 210252 70366 210464 70394
rect 210332 69556 210384 69562
rect 210332 69498 210384 69504
rect 210148 66224 210200 66230
rect 210148 66166 210200 66172
rect 210344 64874 210372 69498
rect 210436 68474 210464 70366
rect 210712 69562 210740 84102
rect 210804 75002 210832 93826
rect 210792 74996 210844 75002
rect 210792 74938 210844 74944
rect 210700 69556 210752 69562
rect 210700 69498 210752 69504
rect 210424 68468 210476 68474
rect 210424 68410 210476 68416
rect 210344 64846 210464 64874
rect 209870 48240 209926 48249
rect 209870 48175 209926 48184
rect 209870 45384 209926 45393
rect 209870 45319 209926 45328
rect 209778 17912 209834 17921
rect 209778 17847 209834 17856
rect 208412 16546 208624 16574
rect 207756 3324 207808 3330
rect 207756 3266 207808 3272
rect 207388 2984 207440 2990
rect 207388 2926 207440 2932
rect 207400 480 207428 2926
rect 208596 480 208624 16546
rect 209884 6914 209912 45319
rect 209792 6886 209912 6914
rect 209792 480 209820 6886
rect 210436 3398 210464 64846
rect 211066 48240 211122 48249
rect 211066 48175 211122 48184
rect 211080 47569 211108 48175
rect 211066 47560 211122 47569
rect 211066 47495 211122 47504
rect 211172 38593 211200 192442
rect 211250 189952 211306 189961
rect 211250 189887 211306 189896
rect 211264 44130 211292 189887
rect 211356 74934 211384 198562
rect 211528 198552 211580 198558
rect 211528 198494 211580 198500
rect 211436 198008 211488 198014
rect 211436 197950 211488 197956
rect 211448 79354 211476 197950
rect 211540 80753 211568 198494
rect 212724 198416 212776 198422
rect 212724 198358 212776 198364
rect 212632 198280 212684 198286
rect 212632 198222 212684 198228
rect 211804 198144 211856 198150
rect 211804 198086 211856 198092
rect 211712 190392 211764 190398
rect 211712 190334 211764 190340
rect 211620 187128 211672 187134
rect 211620 187070 211672 187076
rect 211526 80744 211582 80753
rect 211526 80679 211582 80688
rect 211436 79348 211488 79354
rect 211436 79290 211488 79296
rect 211344 74928 211396 74934
rect 211344 74870 211396 74876
rect 211632 74225 211660 187070
rect 211724 77654 211752 190334
rect 211816 78742 211844 198086
rect 212538 189680 212594 189689
rect 212538 189615 212594 189624
rect 211896 155440 211948 155446
rect 211896 155382 211948 155388
rect 211804 78736 211856 78742
rect 211804 78678 211856 78684
rect 211816 78606 211844 78678
rect 211804 78600 211856 78606
rect 211804 78542 211856 78548
rect 211908 77897 211936 155382
rect 211988 152516 212040 152522
rect 211988 152458 212040 152464
rect 212000 78033 212028 152458
rect 211986 78024 212042 78033
rect 211986 77959 212042 77968
rect 211894 77888 211950 77897
rect 211894 77823 211950 77832
rect 211712 77648 211764 77654
rect 211712 77590 211764 77596
rect 211618 74216 211674 74225
rect 211618 74151 211674 74160
rect 211632 70394 211660 74151
rect 211632 70366 211844 70394
rect 211252 44124 211304 44130
rect 211252 44066 211304 44072
rect 211158 38584 211214 38593
rect 211158 38519 211214 38528
rect 211066 17912 211122 17921
rect 211066 17847 211122 17856
rect 211080 17241 211108 17847
rect 211066 17232 211122 17241
rect 211066 17167 211122 17176
rect 211816 4146 211844 70366
rect 212448 44124 212500 44130
rect 212448 44066 212500 44072
rect 212460 43450 212488 44066
rect 212448 43444 212500 43450
rect 212448 43386 212500 43392
rect 212446 38584 212502 38593
rect 212446 38519 212502 38528
rect 212460 37913 212488 38519
rect 212446 37904 212502 37913
rect 212446 37839 212502 37848
rect 212552 21593 212580 189615
rect 212644 59265 212672 198222
rect 212736 62121 212764 198358
rect 212908 198348 212960 198354
rect 212908 198290 212960 198296
rect 212814 198112 212870 198121
rect 212814 198047 212870 198056
rect 212828 66881 212856 198047
rect 212920 67590 212948 198290
rect 212998 197976 213054 197985
rect 212998 197911 213054 197920
rect 213012 71777 213040 197911
rect 213092 193860 213144 193866
rect 213092 193802 213144 193808
rect 213104 78198 213132 193802
rect 213184 158092 213236 158098
rect 213184 158034 213236 158040
rect 213092 78192 213144 78198
rect 213092 78134 213144 78140
rect 213196 77178 213224 158034
rect 213184 77172 213236 77178
rect 213184 77114 213236 77120
rect 212998 71768 213054 71777
rect 212998 71703 213054 71712
rect 212908 67584 212960 67590
rect 212908 67526 212960 67532
rect 213828 67584 213880 67590
rect 213828 67526 213880 67532
rect 213840 66978 213868 67526
rect 213828 66972 213880 66978
rect 213828 66914 213880 66920
rect 212814 66872 212870 66881
rect 212814 66807 212870 66816
rect 213932 64297 213960 200126
rect 214012 199708 214064 199714
rect 214012 199650 214064 199656
rect 213918 64288 213974 64297
rect 213918 64223 213974 64232
rect 213918 62792 213974 62801
rect 213918 62727 213974 62736
rect 212722 62112 212778 62121
rect 212722 62047 212778 62056
rect 213826 62112 213882 62121
rect 213826 62047 213882 62056
rect 213840 61441 213868 62047
rect 213826 61432 213882 61441
rect 213826 61367 213882 61376
rect 212630 59256 212686 59265
rect 212630 59191 212686 59200
rect 213826 59256 213882 59265
rect 213826 59191 213882 59200
rect 213840 58585 213868 59191
rect 213826 58576 213882 58585
rect 213826 58511 213882 58520
rect 212630 30968 212686 30977
rect 212630 30903 212686 30912
rect 212538 21584 212594 21593
rect 212538 21519 212594 21528
rect 212644 16574 212672 30903
rect 213932 16574 213960 62727
rect 214024 52057 214052 199650
rect 215852 199640 215904 199646
rect 215852 199582 215904 199588
rect 215576 199368 215628 199374
rect 215576 199310 215628 199316
rect 215484 198212 215536 198218
rect 215484 198154 215536 198160
rect 214380 198076 214432 198082
rect 214380 198018 214432 198024
rect 214288 189984 214340 189990
rect 214288 189926 214340 189932
rect 214196 187264 214248 187270
rect 214196 187206 214248 187212
rect 214104 187196 214156 187202
rect 214104 187138 214156 187144
rect 214116 57905 214144 187138
rect 214208 60722 214236 187206
rect 214300 70378 214328 189926
rect 214392 80730 214420 198018
rect 215300 196784 215352 196790
rect 215300 196726 215352 196732
rect 214472 158160 214524 158166
rect 214472 158102 214524 158108
rect 214484 80866 214512 158102
rect 214654 151056 214710 151065
rect 214654 150991 214710 151000
rect 214564 141432 214616 141438
rect 214564 141374 214616 141380
rect 214576 81122 214604 141374
rect 214668 93854 214696 150991
rect 214668 93826 214788 93854
rect 214564 81116 214616 81122
rect 214564 81058 214616 81064
rect 214484 80838 214604 80866
rect 214392 80702 214512 80730
rect 214484 80054 214512 80702
rect 214392 80026 214512 80054
rect 214392 79354 214420 80026
rect 214380 79348 214432 79354
rect 214380 79290 214432 79296
rect 214392 78878 214420 79290
rect 214380 78872 214432 78878
rect 214380 78814 214432 78820
rect 214576 76838 214604 80838
rect 214760 77081 214788 93826
rect 214840 81116 214892 81122
rect 214840 81058 214892 81064
rect 214746 77072 214802 77081
rect 214746 77007 214802 77016
rect 214564 76832 214616 76838
rect 214564 76774 214616 76780
rect 214288 70372 214340 70378
rect 214288 70314 214340 70320
rect 214300 69766 214328 70314
rect 214288 69760 214340 69766
rect 214288 69702 214340 69708
rect 214852 65890 214880 81058
rect 214840 65884 214892 65890
rect 214840 65826 214892 65832
rect 214196 60716 214248 60722
rect 214196 60658 214248 60664
rect 214472 60716 214524 60722
rect 214472 60658 214524 60664
rect 214484 60178 214512 60658
rect 214472 60172 214524 60178
rect 214472 60114 214524 60120
rect 214102 57896 214158 57905
rect 214102 57831 214158 57840
rect 215312 57769 215340 196726
rect 215390 195256 215446 195265
rect 215390 195191 215446 195200
rect 215404 60625 215432 195191
rect 215496 63345 215524 198154
rect 215588 68513 215616 199310
rect 215668 196716 215720 196722
rect 215668 196658 215720 196664
rect 215574 68504 215630 68513
rect 215574 68439 215630 68448
rect 215680 68354 215708 196658
rect 215760 187060 215812 187066
rect 215760 187002 215812 187008
rect 215588 68326 215708 68354
rect 215588 67522 215616 68326
rect 215772 67561 215800 187002
rect 215864 80918 215892 199582
rect 216680 196648 216732 196654
rect 216680 196590 216732 196596
rect 215852 80912 215904 80918
rect 215852 80854 215904 80860
rect 216692 75546 216720 196590
rect 218152 195288 218204 195294
rect 218152 195230 218204 195236
rect 216772 191208 216824 191214
rect 216772 191150 216824 191156
rect 216680 75540 216732 75546
rect 216680 75482 216732 75488
rect 216680 75404 216732 75410
rect 216680 75346 216732 75352
rect 215758 67552 215814 67561
rect 215576 67516 215628 67522
rect 215758 67487 215814 67496
rect 215576 67458 215628 67464
rect 215588 66910 215616 67458
rect 215576 66904 215628 66910
rect 215576 66846 215628 66852
rect 215482 63336 215538 63345
rect 215482 63271 215538 63280
rect 215496 62801 215524 63271
rect 215482 62792 215538 62801
rect 215482 62727 215538 62736
rect 215390 60616 215446 60625
rect 215390 60551 215446 60560
rect 215404 60081 215432 60551
rect 215390 60072 215446 60081
rect 215390 60007 215446 60016
rect 215298 57760 215354 57769
rect 215298 57695 215354 57704
rect 215312 57225 215340 57695
rect 215298 57216 215354 57225
rect 215298 57151 215354 57160
rect 214010 52048 214066 52057
rect 214010 51983 214066 51992
rect 215300 47660 215352 47666
rect 215300 47602 215352 47608
rect 212644 16546 213408 16574
rect 213932 16546 214512 16574
rect 211804 4140 211856 4146
rect 211804 4082 211856 4088
rect 212172 4004 212224 4010
rect 212172 3946 212224 3952
rect 210424 3392 210476 3398
rect 210424 3334 210476 3340
rect 210976 3324 211028 3330
rect 210976 3266 211028 3272
rect 210988 480 211016 3266
rect 212184 480 212212 3946
rect 213380 480 213408 16546
rect 214484 480 214512 16546
rect 199078 354 199190 480
rect 198752 326 199190 354
rect 199078 -960 199190 326
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215312 354 215340 47602
rect 216692 16574 216720 75346
rect 216784 63481 216812 191150
rect 216956 189916 217008 189922
rect 216956 189858 217008 189864
rect 216862 155408 216918 155417
rect 216862 155343 216918 155352
rect 216770 63472 216826 63481
rect 216770 63407 216826 63416
rect 216772 46912 216824 46918
rect 216772 46854 216824 46860
rect 216784 46238 216812 46854
rect 216772 46232 216824 46238
rect 216772 46174 216824 46180
rect 216876 37233 216904 155343
rect 216968 72826 216996 189858
rect 218058 186960 218114 186969
rect 218058 186895 218114 186904
rect 217140 158024 217192 158030
rect 217140 157966 217192 157972
rect 217048 148368 217100 148374
rect 217048 148310 217100 148316
rect 216956 72820 217008 72826
rect 216956 72762 217008 72768
rect 216968 72350 216996 72762
rect 216956 72344 217008 72350
rect 216956 72286 217008 72292
rect 217060 46918 217088 148310
rect 217152 79558 217180 157966
rect 217232 151088 217284 151094
rect 217232 151030 217284 151036
rect 217140 79552 217192 79558
rect 217140 79494 217192 79500
rect 217244 79370 217272 151030
rect 217324 141500 217376 141506
rect 217324 141442 217376 141448
rect 217152 79342 217272 79370
rect 217152 77246 217180 79342
rect 217140 77240 217192 77246
rect 217140 77182 217192 77188
rect 217152 76770 217180 77182
rect 217336 76838 217364 141442
rect 217416 79552 217468 79558
rect 217416 79494 217468 79500
rect 217324 76832 217376 76838
rect 217324 76774 217376 76780
rect 217140 76764 217192 76770
rect 217140 76706 217192 76712
rect 217428 76673 217456 79494
rect 217138 76664 217194 76673
rect 217138 76599 217194 76608
rect 217414 76664 217470 76673
rect 217414 76599 217470 76608
rect 217152 76129 217180 76599
rect 217138 76120 217194 76129
rect 217138 76055 217194 76064
rect 217048 46912 217100 46918
rect 218072 46889 218100 186895
rect 218164 74458 218192 195230
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 218336 191140 218388 191146
rect 218336 191082 218388 191088
rect 218244 189848 218296 189854
rect 218244 189790 218296 189796
rect 218152 74452 218204 74458
rect 218152 74394 218204 74400
rect 218164 73914 218192 74394
rect 218256 74186 218284 189790
rect 218348 74526 218376 191082
rect 218428 189780 218480 189786
rect 218428 189722 218480 189728
rect 218336 74520 218388 74526
rect 218336 74462 218388 74468
rect 218244 74180 218296 74186
rect 218244 74122 218296 74128
rect 218242 74080 218298 74089
rect 218348 74050 218376 74462
rect 218440 74361 218468 189722
rect 218520 186992 218572 186998
rect 218520 186934 218572 186940
rect 218426 74352 218482 74361
rect 218426 74287 218482 74296
rect 218242 74015 218298 74024
rect 218336 74044 218388 74050
rect 218152 73908 218204 73914
rect 218152 73850 218204 73856
rect 218256 73409 218284 74015
rect 218336 73986 218388 73992
rect 218440 73953 218468 74287
rect 218532 74089 218560 186934
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580184 178090 580212 179143
rect 580172 178084 580224 178090
rect 580172 178026 580224 178032
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580184 165646 580212 165815
rect 580172 165640 580224 165646
rect 580172 165582 580224 165588
rect 579986 152688 580042 152697
rect 579986 152623 580042 152632
rect 580000 151842 580028 152623
rect 579988 151836 580040 151842
rect 579988 151778 580040 151784
rect 580448 150476 580500 150482
rect 580448 150418 580500 150424
rect 580264 149116 580316 149122
rect 580264 149058 580316 149064
rect 467102 142352 467158 142361
rect 467102 142287 467158 142296
rect 464342 141264 464398 141273
rect 464342 141199 464398 141208
rect 327724 139460 327776 139466
rect 327724 139402 327776 139408
rect 234620 80912 234672 80918
rect 234620 80854 234672 80860
rect 218612 74180 218664 74186
rect 218612 74122 218664 74128
rect 218518 74080 218574 74089
rect 218518 74015 218574 74024
rect 218426 73944 218482 73953
rect 218426 73879 218482 73888
rect 218242 73400 218298 73409
rect 218242 73335 218298 73344
rect 218624 72894 218652 74122
rect 218152 72888 218204 72894
rect 218152 72830 218204 72836
rect 218612 72888 218664 72894
rect 218612 72830 218664 72836
rect 229744 72888 229796 72894
rect 229744 72830 229796 72836
rect 218164 72282 218192 72830
rect 218152 72276 218204 72282
rect 218152 72218 218204 72224
rect 220818 68504 220874 68513
rect 220818 68439 220874 68448
rect 220084 64320 220136 64326
rect 220084 64262 220136 64268
rect 217048 46854 217100 46860
rect 218058 46880 218114 46889
rect 218058 46815 218114 46824
rect 218152 42356 218204 42362
rect 218152 42298 218204 42304
rect 216862 37224 216918 37233
rect 216862 37159 216918 37168
rect 217230 37224 217286 37233
rect 217230 37159 217286 37168
rect 217244 36553 217272 37159
rect 217230 36544 217286 36553
rect 217230 36479 217286 36488
rect 218164 16574 218192 42298
rect 219440 17468 219492 17474
rect 219440 17410 219492 17416
rect 219452 16574 219480 17410
rect 216692 16546 216904 16574
rect 218164 16546 219296 16574
rect 219452 16546 220032 16574
rect 216496 4072 216548 4078
rect 216680 4072 216732 4078
rect 216548 4020 216680 4026
rect 216496 4014 216732 4020
rect 216508 3998 216720 4014
rect 216876 480 216904 16546
rect 217324 4140 217376 4146
rect 217324 4082 217376 4088
rect 217336 4010 217364 4082
rect 217324 4004 217376 4010
rect 217324 3946 217376 3952
rect 218060 3392 218112 3398
rect 218060 3334 218112 3340
rect 218072 480 218100 3334
rect 219268 480 219296 16546
rect 215638 354 215750 480
rect 215312 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220004 354 220032 16546
rect 220096 2990 220124 64262
rect 220832 16574 220860 68439
rect 227718 67552 227774 67561
rect 227718 67487 227774 67496
rect 223580 65680 223632 65686
rect 223580 65622 223632 65628
rect 222200 49156 222252 49162
rect 222200 49098 222252 49104
rect 222212 16574 222240 49098
rect 220832 16546 221136 16574
rect 222212 16546 222792 16574
rect 220084 2984 220136 2990
rect 220084 2926 220136 2932
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 221108 354 221136 16546
rect 222764 480 222792 16546
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 220422 -960 220534 326
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223592 354 223620 65622
rect 225604 50380 225656 50386
rect 225604 50322 225656 50328
rect 225616 3398 225644 50322
rect 227732 16574 227760 67487
rect 229100 29980 229152 29986
rect 229100 29922 229152 29928
rect 229112 16574 229140 29922
rect 227732 16546 228312 16574
rect 229112 16546 229416 16574
rect 227536 7880 227588 7886
rect 227536 7822 227588 7828
rect 225604 3392 225656 3398
rect 225604 3334 225656 3340
rect 226340 3392 226392 3398
rect 226340 3334 226392 3340
rect 225144 2984 225196 2990
rect 225144 2926 225196 2932
rect 225156 480 225184 2926
rect 226352 480 226380 3334
rect 227548 480 227576 7822
rect 223918 354 224030 480
rect 223592 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228284 354 228312 16546
rect 228702 354 228814 480
rect 228284 326 228814 354
rect 229388 354 229416 16546
rect 229756 4146 229784 72830
rect 231858 60208 231914 60217
rect 231858 60143 231914 60152
rect 230952 4146 231164 4162
rect 229744 4140 229796 4146
rect 229744 4082 229796 4088
rect 230940 4140 231164 4146
rect 230992 4134 231164 4140
rect 230940 4082 230992 4088
rect 231136 4010 231164 4134
rect 231032 4004 231084 4010
rect 231032 3946 231084 3952
rect 231124 4004 231176 4010
rect 231124 3946 231176 3952
rect 231044 480 231072 3946
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 228702 -960 228814 326
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 231872 354 231900 60143
rect 233240 43512 233292 43518
rect 233240 43454 233292 43460
rect 233252 16574 233280 43454
rect 233252 16546 233464 16574
rect 233436 480 233464 16546
rect 234632 11694 234660 80854
rect 252560 80844 252612 80850
rect 252560 80786 252612 80792
rect 247684 76900 247736 76906
rect 247684 76842 247736 76848
rect 237378 74080 237434 74089
rect 237378 74015 237434 74024
rect 236000 39636 236052 39642
rect 236000 39578 236052 39584
rect 234710 33824 234766 33833
rect 234710 33759 234766 33768
rect 234620 11688 234672 11694
rect 234620 11630 234672 11636
rect 234724 6914 234752 33759
rect 236012 16574 236040 39578
rect 237392 16574 237420 74015
rect 242164 69896 242216 69902
rect 242164 69838 242216 69844
rect 238760 65748 238812 65754
rect 238760 65690 238812 65696
rect 238772 16574 238800 65690
rect 239404 54664 239456 54670
rect 239404 54606 239456 54612
rect 236012 16546 236592 16574
rect 237392 16546 237696 16574
rect 238772 16546 239352 16574
rect 235816 11688 235868 11694
rect 235816 11630 235868 11636
rect 234632 6886 234752 6914
rect 234632 480 234660 6886
rect 235828 480 235856 11630
rect 232198 354 232310 480
rect 231872 326 232310 354
rect 232198 -960 232310 326
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 16546
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 237668 354 237696 16546
rect 239324 480 239352 16546
rect 239416 3398 239444 54606
rect 241704 10600 241756 10606
rect 241704 10542 241756 10548
rect 239404 3392 239456 3398
rect 239404 3334 239456 3340
rect 240508 3392 240560 3398
rect 240508 3334 240560 3340
rect 240520 480 240548 3334
rect 241716 480 241744 10542
rect 242176 3398 242204 69838
rect 245660 62960 245712 62966
rect 245660 62902 245712 62908
rect 242992 28552 243044 28558
rect 242992 28494 243044 28500
rect 243004 16574 243032 28494
rect 245672 16574 245700 62902
rect 243004 16546 244136 16574
rect 245672 16546 245976 16574
rect 242164 3392 242216 3398
rect 242164 3334 242216 3340
rect 242900 3392 242952 3398
rect 242900 3334 242952 3340
rect 242912 480 242940 3334
rect 244108 480 244136 16546
rect 245200 12028 245252 12034
rect 245200 11970 245252 11976
rect 245212 480 245240 11970
rect 238086 354 238198 480
rect 237668 326 238198 354
rect 236982 -960 237094 326
rect 238086 -960 238198 326
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 245948 354 245976 16546
rect 247696 4146 247724 76842
rect 249800 58880 249852 58886
rect 249800 58822 249852 58828
rect 249812 16574 249840 58822
rect 251178 46472 251234 46481
rect 251178 46407 251234 46416
rect 249812 16546 250024 16574
rect 248420 16108 248472 16114
rect 248420 16050 248472 16056
rect 247592 4140 247644 4146
rect 247592 4082 247644 4088
rect 247684 4140 247736 4146
rect 247684 4082 247736 4088
rect 247604 480 247632 4082
rect 246366 354 246478 480
rect 245948 326 246478 354
rect 246366 -960 246478 326
rect 247562 -960 247674 480
rect 248432 354 248460 16050
rect 249996 480 250024 16546
rect 251192 4078 251220 46407
rect 251272 38140 251324 38146
rect 251272 38082 251324 38088
rect 251180 4072 251232 4078
rect 251180 4014 251232 4020
rect 251284 3482 251312 38082
rect 252572 16574 252600 80786
rect 270500 80776 270552 80782
rect 270500 80718 270552 80724
rect 260102 76664 260158 76673
rect 260102 76599 260158 76608
rect 255320 74044 255372 74050
rect 255320 73986 255372 73992
rect 255332 16574 255360 73986
rect 256700 64388 256752 64394
rect 256700 64330 256752 64336
rect 252572 16546 253520 16574
rect 255332 16546 255912 16574
rect 252376 4072 252428 4078
rect 252376 4014 252428 4020
rect 251192 3454 251312 3482
rect 251192 480 251220 3454
rect 252388 480 252416 4014
rect 253492 480 253520 16546
rect 254676 4140 254728 4146
rect 254676 4082 254728 4088
rect 254688 480 254716 4082
rect 255884 480 255912 16546
rect 248758 354 248870 480
rect 248432 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 256712 354 256740 64330
rect 259458 52048 259514 52057
rect 259458 51983 259514 51992
rect 258264 13388 258316 13394
rect 258264 13330 258316 13336
rect 258276 480 258304 13330
rect 259472 3398 259500 51983
rect 259552 6588 259604 6594
rect 259552 6530 259604 6536
rect 259460 3392 259512 3398
rect 259460 3334 259512 3340
rect 259564 3210 259592 6530
rect 259472 3182 259592 3210
rect 259472 480 259500 3182
rect 260116 2922 260144 76599
rect 261484 73976 261536 73982
rect 261484 73918 261536 73924
rect 261496 3398 261524 73918
rect 269118 73808 269174 73817
rect 269118 73743 269174 73752
rect 263598 57624 263654 57633
rect 263598 57559 263654 57568
rect 263612 16574 263640 57559
rect 267740 44872 267792 44878
rect 267740 44814 267792 44820
rect 264980 32632 265032 32638
rect 264980 32574 265032 32580
rect 263612 16546 264192 16574
rect 260656 3392 260708 3398
rect 260656 3334 260708 3340
rect 261484 3392 261536 3398
rect 261484 3334 261536 3340
rect 262956 3392 263008 3398
rect 262956 3334 263008 3340
rect 260104 2916 260156 2922
rect 260104 2858 260156 2864
rect 260668 480 260696 3334
rect 261760 2916 261812 2922
rect 261760 2858 261812 2864
rect 261772 480 261800 2858
rect 262968 480 262996 3334
rect 264164 480 264192 16546
rect 257038 354 257150 480
rect 256712 326 257150 354
rect 257038 -960 257150 326
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 264992 354 265020 32574
rect 266360 18828 266412 18834
rect 266360 18770 266412 18776
rect 266372 16574 266400 18770
rect 266372 16546 266584 16574
rect 266556 480 266584 16546
rect 267752 480 267780 44814
rect 267832 36712 267884 36718
rect 267832 36654 267884 36660
rect 267844 16574 267872 36654
rect 269132 16574 269160 73743
rect 270512 16574 270540 80718
rect 288440 80708 288492 80714
rect 288440 80650 288492 80656
rect 284298 73944 284354 73953
rect 284298 73879 284354 73888
rect 274640 67108 274692 67114
rect 274640 67050 274692 67056
rect 274652 16574 274680 67050
rect 277400 61532 277452 61538
rect 277400 61474 277452 61480
rect 276110 43888 276166 43897
rect 276110 43823 276166 43832
rect 275284 27124 275336 27130
rect 275284 27066 275336 27072
rect 267844 16546 268424 16574
rect 269132 16546 270080 16574
rect 270512 16546 270816 16574
rect 274652 16546 274864 16574
rect 265318 354 265430 480
rect 264992 326 265430 354
rect 265318 -960 265430 326
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268396 354 268424 16546
rect 270052 480 270080 16546
rect 268814 354 268926 480
rect 268396 326 268926 354
rect 268814 -960 268926 326
rect 270010 -960 270122 480
rect 270788 354 270816 16546
rect 272432 14748 272484 14754
rect 272432 14690 272484 14696
rect 272444 480 272472 14690
rect 273628 5024 273680 5030
rect 273628 4966 273680 4972
rect 273640 480 273668 4966
rect 274836 480 274864 16546
rect 275296 3398 275324 27066
rect 276124 16574 276152 43823
rect 277412 16574 277440 61474
rect 281540 58812 281592 58818
rect 281540 58754 281592 58760
rect 278780 25764 278832 25770
rect 278780 25706 278832 25712
rect 278792 16574 278820 25706
rect 280160 20188 280212 20194
rect 280160 20130 280212 20136
rect 280172 16574 280200 20130
rect 276124 16546 276704 16574
rect 277412 16546 278360 16574
rect 278792 16546 279096 16574
rect 280172 16546 280752 16574
rect 275284 3392 275336 3398
rect 275284 3334 275336 3340
rect 276020 3392 276072 3398
rect 276020 3334 276072 3340
rect 276032 480 276060 3334
rect 271206 354 271318 480
rect 270788 326 271318 354
rect 271206 -960 271318 326
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 276676 354 276704 16546
rect 278332 480 278360 16546
rect 277094 354 277206 480
rect 276676 326 277206 354
rect 277094 -960 277206 326
rect 278290 -960 278402 480
rect 279068 354 279096 16546
rect 280724 480 280752 16546
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281552 354 281580 58754
rect 282920 24404 282972 24410
rect 282920 24346 282972 24352
rect 282932 16574 282960 24346
rect 282932 16546 283144 16574
rect 283116 480 283144 16546
rect 284312 480 284340 73879
rect 284390 56264 284446 56273
rect 284390 56199 284446 56208
rect 284404 16574 284432 56199
rect 285680 42288 285732 42294
rect 285680 42230 285732 42236
rect 285692 16574 285720 42230
rect 287060 20120 287112 20126
rect 287060 20062 287112 20068
rect 287072 16574 287100 20062
rect 288452 16574 288480 80650
rect 302238 78704 302294 78713
rect 302238 78639 302294 78648
rect 289820 76832 289872 76838
rect 289820 76774 289872 76780
rect 284404 16546 284984 16574
rect 285692 16546 286640 16574
rect 287072 16546 287376 16574
rect 288452 16546 289032 16574
rect 281878 354 281990 480
rect 281552 326 281990 354
rect 281878 -960 281990 326
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 284956 354 284984 16546
rect 286612 480 286640 16546
rect 285374 354 285486 480
rect 284956 326 285486 354
rect 285374 -960 285486 326
rect 286570 -960 286682 480
rect 287348 354 287376 16546
rect 289004 480 289032 16546
rect 287766 354 287878 480
rect 287348 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 289832 354 289860 76774
rect 296720 76764 296772 76770
rect 296720 76706 296772 76712
rect 295340 65612 295392 65618
rect 295340 65554 295392 65560
rect 292580 62892 292632 62898
rect 292580 62834 292632 62840
rect 291200 20052 291252 20058
rect 291200 19994 291252 20000
rect 291212 16574 291240 19994
rect 291212 16546 291424 16574
rect 291396 480 291424 16546
rect 292592 480 292620 62834
rect 292672 46232 292724 46238
rect 292672 46174 292724 46180
rect 292684 16574 292712 46174
rect 293958 37904 294014 37913
rect 293958 37839 294014 37848
rect 293972 16574 294000 37839
rect 295352 16574 295380 65554
rect 296732 16574 296760 76706
rect 299480 60172 299532 60178
rect 299480 60114 299532 60120
rect 292684 16546 293264 16574
rect 293972 16546 294920 16574
rect 295352 16546 295656 16574
rect 296732 16546 297312 16574
rect 290158 354 290270 480
rect 289832 326 290270 354
rect 290158 -960 290270 326
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 354 293264 16546
rect 294892 480 294920 16546
rect 293654 354 293766 480
rect 293236 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 295628 354 295656 16546
rect 297284 480 297312 16546
rect 298468 4004 298520 4010
rect 298468 3946 298520 3952
rect 298480 480 298508 3946
rect 299492 3482 299520 60114
rect 299572 31340 299624 31346
rect 299572 31282 299624 31288
rect 299584 4010 299612 31282
rect 300858 17232 300914 17241
rect 300858 17167 300914 17176
rect 300872 16574 300900 17167
rect 302252 16574 302280 78639
rect 324320 76696 324372 76702
rect 324320 76638 324372 76644
rect 305000 75336 305052 75342
rect 305000 75278 305052 75284
rect 303620 29912 303672 29918
rect 303620 29854 303672 29860
rect 303632 16574 303660 29854
rect 305012 16574 305040 75278
rect 322940 73840 322992 73846
rect 322940 73782 322992 73788
rect 318800 72752 318852 72758
rect 318800 72694 318852 72700
rect 317420 67040 317472 67046
rect 317420 66982 317472 66988
rect 306378 64288 306434 64297
rect 306378 64223 306434 64232
rect 300872 16546 301544 16574
rect 302252 16546 303200 16574
rect 303632 16546 303936 16574
rect 305012 16546 305592 16574
rect 299572 4004 299624 4010
rect 299572 3946 299624 3952
rect 300768 4004 300820 4010
rect 300768 3946 300820 3952
rect 299492 3454 299704 3482
rect 299676 480 299704 3454
rect 300780 480 300808 3946
rect 296046 354 296158 480
rect 295628 326 296158 354
rect 296046 -960 296158 326
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 354 301544 16546
rect 303172 480 303200 16546
rect 301934 354 302046 480
rect 301516 326 302046 354
rect 301934 -960 302046 326
rect 303130 -960 303242 480
rect 303908 354 303936 16546
rect 305564 480 305592 16546
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306392 354 306420 64223
rect 313280 61600 313332 61606
rect 313280 61542 313332 61548
rect 309140 40996 309192 41002
rect 309140 40938 309192 40944
rect 307022 36680 307078 36689
rect 307022 36615 307078 36624
rect 307036 3398 307064 36615
rect 309152 16574 309180 40938
rect 311162 35184 311218 35193
rect 311162 35119 311218 35128
rect 310520 22976 310572 22982
rect 310520 22918 310572 22924
rect 310532 16574 310560 22918
rect 309152 16546 309824 16574
rect 310532 16546 311112 16574
rect 307944 13320 307996 13326
rect 307944 13262 307996 13268
rect 307024 3392 307076 3398
rect 307024 3334 307076 3340
rect 307956 480 307984 13262
rect 309048 3392 309100 3398
rect 309048 3334 309100 3340
rect 309060 480 309088 3334
rect 306718 354 306830 480
rect 306392 326 306830 354
rect 306718 -960 306830 326
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 354 309824 16546
rect 311084 3482 311112 16546
rect 311176 4010 311204 35119
rect 313292 16574 313320 61542
rect 315304 54596 315356 54602
rect 315304 54538 315356 54544
rect 313292 16546 313872 16574
rect 311164 4004 311216 4010
rect 311164 3946 311216 3952
rect 312636 4004 312688 4010
rect 312636 3946 312688 3952
rect 311084 3454 311480 3482
rect 311452 480 311480 3454
rect 312648 480 312676 3946
rect 313844 480 313872 16546
rect 314660 14680 314712 14686
rect 314660 14622 314712 14628
rect 310214 354 310326 480
rect 309796 326 310326 354
rect 310214 -960 310326 326
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314672 354 314700 14622
rect 315316 4146 315344 54538
rect 317432 16574 317460 66982
rect 318812 16574 318840 72694
rect 320178 51912 320234 51921
rect 320178 51847 320234 51856
rect 320192 16574 320220 51847
rect 321560 35420 321612 35426
rect 321560 35362 321612 35368
rect 321572 16574 321600 35362
rect 317432 16546 318104 16574
rect 318812 16546 319760 16574
rect 320192 16546 320496 16574
rect 321572 16546 322152 16574
rect 316224 9104 316276 9110
rect 316224 9046 316276 9052
rect 315304 4140 315356 4146
rect 315304 4082 315356 4088
rect 316236 480 316264 9046
rect 317328 4140 317380 4146
rect 317328 4082 317380 4088
rect 317340 480 317368 4082
rect 314998 354 315110 480
rect 314672 326 315110 354
rect 314998 -960 315110 326
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 16546
rect 319732 480 319760 16546
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320468 354 320496 16546
rect 322124 480 322152 16546
rect 320886 354 320998 480
rect 320468 326 320998 354
rect 320886 -960 320998 326
rect 322082 -960 322194 480
rect 322952 354 322980 73782
rect 323584 72684 323636 72690
rect 323584 72626 323636 72632
rect 323596 4146 323624 72626
rect 323584 4140 323636 4146
rect 323584 4082 323636 4088
rect 324332 3210 324360 76638
rect 327736 73166 327764 139402
rect 464356 86970 464384 141199
rect 467116 100706 467144 142287
rect 574742 141128 574798 141137
rect 574742 141063 574798 141072
rect 467104 100700 467156 100706
rect 467104 100642 467156 100648
rect 464344 86964 464396 86970
rect 464344 86906 464396 86912
rect 523130 80744 523186 80753
rect 523130 80679 523186 80688
rect 340880 79484 340932 79490
rect 340880 79426 340932 79432
rect 327724 73160 327776 73166
rect 327724 73102 327776 73108
rect 332600 72616 332652 72622
rect 332600 72558 332652 72564
rect 327080 58744 327132 58750
rect 327080 58686 327132 58692
rect 324412 39568 324464 39574
rect 324412 39510 324464 39516
rect 324424 3398 324452 39510
rect 327092 16574 327120 58686
rect 331218 56128 331274 56137
rect 331218 56063 331274 56072
rect 329840 18760 329892 18766
rect 329840 18702 329892 18708
rect 329852 16574 329880 18702
rect 327092 16546 328040 16574
rect 329852 16546 330432 16574
rect 326804 4140 326856 4146
rect 326804 4082 326856 4088
rect 324412 3392 324464 3398
rect 324412 3334 324464 3340
rect 325608 3392 325660 3398
rect 325608 3334 325660 3340
rect 324332 3182 324452 3210
rect 324424 480 324452 3182
rect 325620 480 325648 3334
rect 326816 480 326844 4082
rect 328012 480 328040 16546
rect 328736 11960 328788 11966
rect 328736 11902 328788 11908
rect 323278 354 323390 480
rect 322952 326 323390 354
rect 323278 -960 323390 326
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 328748 354 328776 11902
rect 330404 480 330432 16546
rect 329166 354 329278 480
rect 328748 326 329278 354
rect 329166 -960 329278 326
rect 330362 -960 330474 480
rect 331232 354 331260 56063
rect 332612 3398 332640 72558
rect 333978 53272 334034 53281
rect 333978 53207 334034 53216
rect 332692 40928 332744 40934
rect 332692 40870 332744 40876
rect 332600 3392 332652 3398
rect 332600 3334 332652 3340
rect 332704 480 332732 40870
rect 333992 16574 334020 53207
rect 338118 50688 338174 50697
rect 338118 50623 338174 50632
rect 336738 21584 336794 21593
rect 336738 21519 336794 21528
rect 336752 16574 336780 21519
rect 338132 16574 338160 50623
rect 339500 28484 339552 28490
rect 339500 28426 339552 28432
rect 333992 16546 334664 16574
rect 336752 16546 337056 16574
rect 338132 16546 338712 16574
rect 333888 3392 333940 3398
rect 333888 3334 333940 3340
rect 333900 480 333928 3334
rect 331558 354 331670 480
rect 331232 326 331670 354
rect 331558 -960 331670 326
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 354 334664 16546
rect 336280 10532 336332 10538
rect 336280 10474 336332 10480
rect 336292 480 336320 10474
rect 335054 354 335166 480
rect 334636 326 335166 354
rect 335054 -960 335166 326
rect 336250 -960 336362 480
rect 337028 354 337056 16546
rect 338684 480 338712 16546
rect 337446 354 337558 480
rect 337028 326 337558 354
rect 337446 -960 337558 326
rect 338642 -960 338754 480
rect 339512 354 339540 28426
rect 340892 3398 340920 79426
rect 376760 79416 376812 79422
rect 376760 79358 376812 79364
rect 353300 76628 353352 76634
rect 353300 76570 353352 76576
rect 347780 73908 347832 73914
rect 347780 73850 347832 73856
rect 342904 72820 342956 72826
rect 342904 72762 342956 72768
rect 340972 72548 341024 72554
rect 340972 72490 341024 72496
rect 340880 3392 340932 3398
rect 340880 3334 340932 3340
rect 340984 480 341012 72490
rect 342916 3398 342944 72762
rect 345020 64252 345072 64258
rect 345020 64194 345072 64200
rect 345032 16574 345060 64194
rect 346400 32564 346452 32570
rect 346400 32506 346452 32512
rect 346412 16574 346440 32506
rect 347792 16574 347820 73850
rect 351920 60104 351972 60110
rect 351920 60046 351972 60052
rect 349160 57248 349212 57254
rect 349160 57190 349212 57196
rect 349172 16574 349200 57190
rect 350538 21448 350594 21457
rect 350538 21383 350594 21392
rect 350552 16574 350580 21383
rect 351932 16574 351960 60046
rect 353312 16574 353340 76570
rect 367100 76560 367152 76566
rect 367100 76502 367152 76508
rect 362960 69828 363012 69834
rect 362960 69770 363012 69776
rect 358820 68332 358872 68338
rect 358820 68274 358872 68280
rect 356060 51196 356112 51202
rect 356060 51138 356112 51144
rect 354678 21312 354734 21321
rect 354678 21247 354734 21256
rect 354692 16574 354720 21247
rect 356072 16574 356100 51138
rect 357440 33992 357492 33998
rect 357440 33934 357492 33940
rect 345032 16546 345336 16574
rect 346412 16546 346992 16574
rect 347792 16546 348096 16574
rect 349172 16546 349292 16574
rect 350552 16546 351224 16574
rect 351932 16546 352880 16574
rect 353312 16546 353616 16574
rect 354692 16546 355272 16574
rect 356072 16546 356376 16574
rect 343364 7812 343416 7818
rect 343364 7754 343416 7760
rect 342168 3392 342220 3398
rect 342168 3334 342220 3340
rect 342904 3392 342956 3398
rect 342904 3334 342956 3340
rect 342180 480 342208 3334
rect 343376 480 343404 7754
rect 344560 3392 344612 3398
rect 344560 3334 344612 3340
rect 344572 480 344600 3334
rect 339838 354 339950 480
rect 339512 326 339950 354
rect 339838 -960 339950 326
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345308 354 345336 16546
rect 346964 480 346992 16546
rect 348068 480 348096 16546
rect 349264 480 349292 16546
rect 350448 6520 350500 6526
rect 350448 6462 350500 6468
rect 350460 480 350488 6462
rect 345726 354 345838 480
rect 345308 326 345838 354
rect 345726 -960 345838 326
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351196 354 351224 16546
rect 352852 480 352880 16546
rect 351614 354 351726 480
rect 351196 326 351726 354
rect 351614 -960 351726 326
rect 352810 -960 352922 480
rect 353588 354 353616 16546
rect 355244 480 355272 16546
rect 356348 480 356376 16546
rect 357452 3210 357480 33934
rect 357532 19984 357584 19990
rect 357532 19926 357584 19932
rect 357544 3398 357572 19926
rect 358832 16574 358860 68274
rect 360200 31272 360252 31278
rect 360200 31214 360252 31220
rect 360212 16574 360240 31214
rect 360844 28416 360896 28422
rect 360844 28358 360896 28364
rect 358832 16546 359504 16574
rect 360212 16546 360792 16574
rect 357532 3392 357584 3398
rect 357532 3334 357584 3340
rect 358728 3392 358780 3398
rect 358728 3334 358780 3340
rect 357452 3182 357572 3210
rect 357544 480 357572 3182
rect 358740 480 358768 3334
rect 354006 354 354118 480
rect 353588 326 354118 354
rect 354006 -960 354118 326
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359476 354 359504 16546
rect 360764 3482 360792 16546
rect 360856 4010 360884 28358
rect 362972 16574 363000 69770
rect 364982 53136 365038 53145
rect 364982 53071 365038 53080
rect 362972 16546 363552 16574
rect 360844 4004 360896 4010
rect 360844 3946 360896 3952
rect 362316 4004 362368 4010
rect 362316 3946 362368 3952
rect 360764 3454 361160 3482
rect 361132 480 361160 3454
rect 362328 480 362356 3946
rect 363524 480 363552 16546
rect 364616 16040 364668 16046
rect 364616 15982 364668 15988
rect 364628 480 364656 15982
rect 364996 3398 365024 53071
rect 367112 16574 367140 76502
rect 368480 72480 368532 72486
rect 368480 72422 368532 72428
rect 368492 16574 368520 72422
rect 372618 62928 372674 62937
rect 372618 62863 372674 62872
rect 369858 54632 369914 54641
rect 369858 54567 369914 54576
rect 369872 16574 369900 54567
rect 372632 16574 372660 62863
rect 373998 50552 374054 50561
rect 373998 50487 374054 50496
rect 367112 16546 367784 16574
rect 368492 16546 369440 16574
rect 369872 16546 370176 16574
rect 372632 16546 372936 16574
rect 365812 7744 365864 7750
rect 365812 7686 365864 7692
rect 364984 3392 365036 3398
rect 364984 3334 365036 3340
rect 365824 480 365852 7686
rect 367008 3392 367060 3398
rect 367008 3334 367060 3340
rect 367020 480 367048 3334
rect 359894 354 360006 480
rect 359476 326 360006 354
rect 359894 -960 360006 326
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 354 367784 16546
rect 369412 480 369440 16546
rect 368174 354 368286 480
rect 367756 326 368286 354
rect 368174 -960 368286 326
rect 369370 -960 369482 480
rect 370148 354 370176 16546
rect 371700 4956 371752 4962
rect 371700 4898 371752 4904
rect 371712 480 371740 4898
rect 372908 480 372936 16546
rect 374012 1170 374040 50487
rect 374092 27056 374144 27062
rect 374092 26998 374144 27004
rect 374104 3398 374132 26998
rect 376772 16574 376800 79358
rect 448520 79348 448572 79354
rect 448520 79290 448572 79296
rect 393320 78124 393372 78130
rect 393320 78066 393372 78072
rect 389178 76528 389234 76537
rect 389178 76463 389234 76472
rect 380900 58676 380952 58682
rect 380900 58618 380952 58624
rect 378784 33924 378836 33930
rect 378784 33866 378836 33872
rect 378140 25696 378192 25702
rect 378140 25638 378192 25644
rect 378152 16574 378180 25638
rect 376772 16546 377720 16574
rect 378152 16546 378456 16574
rect 376024 11892 376076 11898
rect 376024 11834 376076 11840
rect 374092 3392 374144 3398
rect 374092 3334 374144 3340
rect 375288 3392 375340 3398
rect 375288 3334 375340 3340
rect 374012 1142 374132 1170
rect 374104 480 374132 1142
rect 375300 480 375328 3334
rect 370566 354 370678 480
rect 370148 326 370678 354
rect 370566 -960 370678 326
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 354 376064 11834
rect 377692 480 377720 16546
rect 376454 354 376566 480
rect 376036 326 376566 354
rect 376454 -960 376566 326
rect 377650 -960 377762 480
rect 378428 354 378456 16546
rect 378796 3398 378824 33866
rect 380912 16574 380940 58618
rect 382922 55992 382978 56001
rect 382922 55927 382978 55936
rect 382280 54528 382332 54534
rect 382280 54470 382332 54476
rect 380912 16546 381216 16574
rect 378784 3392 378836 3398
rect 378784 3334 378836 3340
rect 379980 3392 380032 3398
rect 379980 3334 380032 3340
rect 379992 480 380020 3334
rect 381188 480 381216 16546
rect 382292 3398 382320 54470
rect 382372 13252 382424 13258
rect 382372 13194 382424 13200
rect 382280 3392 382332 3398
rect 382280 3334 382332 3340
rect 382384 480 382412 13194
rect 382936 3126 382964 55927
rect 387798 49056 387854 49065
rect 387798 48991 387854 49000
rect 385960 14612 386012 14618
rect 385960 14554 386012 14560
rect 383568 3392 383620 3398
rect 383568 3334 383620 3340
rect 382924 3120 382976 3126
rect 382924 3062 382976 3068
rect 383580 480 383608 3334
rect 384764 3120 384816 3126
rect 384764 3062 384816 3068
rect 384776 480 384804 3062
rect 385972 480 386000 14554
rect 386696 10464 386748 10470
rect 386696 10406 386748 10412
rect 378846 354 378958 480
rect 378428 326 378958 354
rect 378846 -960 378958 326
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 386708 354 386736 10406
rect 387126 354 387238 480
rect 386708 326 387238 354
rect 387812 354 387840 48991
rect 389192 16574 389220 76463
rect 391940 53236 391992 53242
rect 391940 53178 391992 53184
rect 390558 45248 390614 45257
rect 390558 45183 390614 45192
rect 389192 16546 389496 16574
rect 389468 480 389496 16546
rect 390572 1834 390600 45183
rect 391952 16574 391980 53178
rect 393332 16574 393360 78066
rect 415492 78056 415544 78062
rect 415492 77998 415544 78004
rect 397460 69760 397512 69766
rect 397460 69702 397512 69708
rect 394698 60072 394754 60081
rect 394698 60007 394754 60016
rect 394712 16574 394740 60007
rect 396080 24336 396132 24342
rect 396080 24278 396132 24284
rect 391952 16546 392624 16574
rect 393332 16546 394280 16574
rect 394712 16546 395384 16574
rect 390652 13184 390704 13190
rect 390652 13126 390704 13132
rect 390560 1828 390612 1834
rect 390560 1770 390612 1776
rect 390664 480 390692 13126
rect 391848 1828 391900 1834
rect 391848 1770 391900 1776
rect 391860 480 391888 1770
rect 388230 354 388342 480
rect 387812 326 388342 354
rect 387126 -960 387238 326
rect 388230 -960 388342 326
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 354 392624 16546
rect 394252 480 394280 16546
rect 395356 480 395384 16546
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 24278
rect 397472 16574 397500 69702
rect 412640 62824 412692 62830
rect 412640 62766 412692 62772
rect 398840 61464 398892 61470
rect 398840 61406 398892 61412
rect 397472 16546 397776 16574
rect 397748 480 397776 16546
rect 398852 3210 398880 61406
rect 402980 60036 403032 60042
rect 402980 59978 403032 59984
rect 400864 51740 400916 51746
rect 400864 51682 400916 51688
rect 398932 22908 398984 22914
rect 398932 22850 398984 22856
rect 398944 3398 398972 22850
rect 400876 3398 400904 51682
rect 402992 16574 403020 59978
rect 405738 47832 405794 47841
rect 405738 47767 405794 47776
rect 404360 32496 404412 32502
rect 404360 32438 404412 32444
rect 402992 16546 403664 16574
rect 401324 3936 401376 3942
rect 401324 3878 401376 3884
rect 398932 3392 398984 3398
rect 398932 3334 398984 3340
rect 400128 3392 400180 3398
rect 400128 3334 400180 3340
rect 400864 3392 400916 3398
rect 400864 3334 400916 3340
rect 398852 3182 398972 3210
rect 398944 480 398972 3182
rect 400140 480 400168 3334
rect 401336 480 401364 3878
rect 402520 3392 402572 3398
rect 402520 3334 402572 3340
rect 402532 480 402560 3334
rect 403636 480 403664 16546
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404372 354 404400 32438
rect 405752 16574 405780 47767
rect 408498 43752 408554 43761
rect 408498 43687 408554 43696
rect 407212 31204 407264 31210
rect 407212 31146 407264 31152
rect 405752 16546 406056 16574
rect 406028 480 406056 16546
rect 407224 480 407252 31146
rect 408512 16574 408540 43687
rect 409880 29844 409932 29850
rect 409880 29786 409932 29792
rect 409892 16574 409920 29786
rect 408512 16546 409184 16574
rect 409892 16546 410840 16574
rect 408408 3868 408460 3874
rect 408408 3810 408460 3816
rect 408420 480 408448 3810
rect 404790 354 404902 480
rect 404372 326 404902 354
rect 404790 -960 404902 326
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 354 409184 16546
rect 410812 480 410840 16546
rect 411904 14544 411956 14550
rect 411904 14486 411956 14492
rect 411916 480 411944 14486
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 354 412680 62766
rect 414662 57488 414718 57497
rect 414662 57423 414718 57432
rect 414296 9036 414348 9042
rect 414296 8978 414348 8984
rect 414308 480 414336 8978
rect 414676 3398 414704 57423
rect 414664 3392 414716 3398
rect 414664 3334 414716 3340
rect 415504 480 415532 77998
rect 422300 77988 422352 77994
rect 422300 77930 422352 77936
rect 418802 50416 418858 50425
rect 418802 50351 418858 50360
rect 418158 25528 418214 25537
rect 418158 25463 418214 25472
rect 418172 16574 418200 25463
rect 418172 16546 418568 16574
rect 417424 11824 417476 11830
rect 417424 11766 417476 11772
rect 416688 3392 416740 3398
rect 416688 3334 416740 3340
rect 416700 480 416728 3334
rect 413070 354 413182 480
rect 412652 326 413182 354
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 11766
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 418540 354 418568 16546
rect 418816 3398 418844 50351
rect 422312 16574 422340 77930
rect 442264 75268 442316 75274
rect 442264 75210 442316 75216
rect 430580 69692 430632 69698
rect 430580 69634 430632 69640
rect 422944 67788 422996 67794
rect 422944 67730 422996 67736
rect 422312 16546 422616 16574
rect 420920 15972 420972 15978
rect 420920 15914 420972 15920
rect 418804 3392 418856 3398
rect 418804 3334 418856 3340
rect 420184 3392 420236 3398
rect 420184 3334 420236 3340
rect 420196 480 420224 3334
rect 418958 354 419070 480
rect 418540 326 419070 354
rect 417854 -960 417966 326
rect 418958 -960 419070 326
rect 420154 -960 420266 480
rect 420932 354 420960 15914
rect 422588 480 422616 16546
rect 422956 3398 422984 67730
rect 423770 59936 423826 59945
rect 423770 59871 423826 59880
rect 422944 3392 422996 3398
rect 422944 3334 422996 3340
rect 423784 480 423812 59871
rect 427818 43616 427874 43625
rect 427818 43551 427874 43560
rect 426440 42220 426492 42226
rect 426440 42162 426492 42168
rect 425060 24268 425112 24274
rect 425060 24210 425112 24216
rect 425072 16574 425100 24210
rect 426452 16574 426480 42162
rect 427832 16574 427860 43551
rect 430592 16574 430620 69634
rect 432604 65544 432656 65550
rect 432604 65486 432656 65492
rect 431960 21412 432012 21418
rect 431960 21354 432012 21360
rect 425072 16546 425744 16574
rect 426452 16546 426848 16574
rect 427832 16546 428504 16574
rect 430592 16546 430896 16574
rect 424968 3392 425020 3398
rect 424968 3334 425020 3340
rect 424980 480 425008 3334
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 425716 354 425744 16546
rect 426134 354 426246 480
rect 425716 326 426246 354
rect 426820 354 426848 16546
rect 428476 480 428504 16546
rect 429660 3800 429712 3806
rect 429660 3742 429712 3748
rect 429672 480 429700 3742
rect 430868 480 430896 16546
rect 431972 3330 432000 21354
rect 432052 10396 432104 10402
rect 432052 10338 432104 10344
rect 431960 3324 432012 3330
rect 431960 3266 432012 3272
rect 432064 480 432092 10338
rect 432616 3398 432644 65486
rect 440238 54496 440294 54505
rect 440238 54431 440294 54440
rect 437480 53168 437532 53174
rect 437480 53110 437532 53116
rect 435548 7676 435600 7682
rect 435548 7618 435600 7624
rect 432604 3392 432656 3398
rect 432604 3334 432656 3340
rect 434444 3392 434496 3398
rect 434444 3334 434496 3340
rect 433248 3324 433300 3330
rect 433248 3266 433300 3272
rect 433260 480 433288 3266
rect 434456 480 434484 3334
rect 435560 480 435588 7618
rect 436744 3732 436796 3738
rect 436744 3674 436796 3680
rect 436756 480 436784 3674
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 426134 -960 426246 326
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437492 354 437520 53110
rect 438860 28348 438912 28354
rect 438860 28290 438912 28296
rect 438872 16574 438900 28290
rect 438872 16546 439176 16574
rect 439148 480 439176 16546
rect 440252 3398 440280 54431
rect 440332 35352 440384 35358
rect 440332 35294 440384 35300
rect 440240 3392 440292 3398
rect 440240 3334 440292 3340
rect 440344 480 440372 35294
rect 442172 15904 442224 15910
rect 442172 15846 442224 15852
rect 442184 3482 442212 15846
rect 442276 3738 442304 75210
rect 444378 45112 444434 45121
rect 444378 45047 444434 45056
rect 444392 16574 444420 45047
rect 445760 17400 445812 17406
rect 445760 17342 445812 17348
rect 444392 16546 445064 16574
rect 443828 6452 443880 6458
rect 443828 6394 443880 6400
rect 442264 3732 442316 3738
rect 442264 3674 442316 3680
rect 442184 3454 442672 3482
rect 441528 3392 441580 3398
rect 441528 3334 441580 3340
rect 441540 480 441568 3334
rect 442644 480 442672 3454
rect 443840 480 443868 6394
rect 445036 480 445064 16546
rect 437910 354 438022 480
rect 437492 326 438022 354
rect 437910 -960 438022 326
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 445772 354 445800 17342
rect 447416 3664 447468 3670
rect 447416 3606 447468 3612
rect 447428 480 447456 3606
rect 448532 3210 448560 79290
rect 480260 78804 480312 78810
rect 480260 78746 480312 78752
rect 465170 78432 465226 78441
rect 465170 78367 465226 78376
rect 456798 78296 456854 78305
rect 456798 78231 456854 78240
rect 450544 55888 450596 55894
rect 450544 55830 450596 55836
rect 448612 49088 448664 49094
rect 448612 49030 448664 49036
rect 448624 3398 448652 49030
rect 450556 4146 450584 55830
rect 454038 46336 454094 46345
rect 454038 46271 454094 46280
rect 450912 6384 450964 6390
rect 450912 6326 450964 6332
rect 450544 4140 450596 4146
rect 450544 4082 450596 4088
rect 448612 3392 448664 3398
rect 448612 3334 448664 3340
rect 449808 3392 449860 3398
rect 449808 3334 449860 3340
rect 448532 3182 448652 3210
rect 448624 480 448652 3182
rect 449820 480 449848 3334
rect 450924 480 450952 6326
rect 453304 6316 453356 6322
rect 453304 6258 453356 6264
rect 452108 4140 452160 4146
rect 452108 4082 452160 4088
rect 452120 480 452148 4082
rect 453316 480 453344 6258
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454052 354 454080 46271
rect 455418 46200 455474 46209
rect 455418 46135 455474 46144
rect 455432 16574 455460 46135
rect 455432 16546 455736 16574
rect 455708 480 455736 16546
rect 456812 3398 456840 78231
rect 460938 72448 460994 72457
rect 460938 72383 460994 72392
rect 459560 61396 459612 61402
rect 459560 61338 459612 61344
rect 458178 43480 458234 43489
rect 458178 43415 458234 43424
rect 458192 16574 458220 43415
rect 459572 16574 459600 61338
rect 460952 16574 460980 72383
rect 464344 51128 464396 51134
rect 464344 51070 464396 51076
rect 463700 39500 463752 39506
rect 463700 39442 463752 39448
rect 462320 39432 462372 39438
rect 462320 39374 462372 39380
rect 458192 16546 459232 16574
rect 459572 16546 459968 16574
rect 460952 16546 461624 16574
rect 456892 4888 456944 4894
rect 456892 4830 456944 4836
rect 456800 3392 456852 3398
rect 456800 3334 456852 3340
rect 456904 480 456932 4830
rect 458088 3392 458140 3398
rect 458088 3334 458140 3340
rect 458100 480 458128 3334
rect 459204 480 459232 16546
rect 454470 354 454582 480
rect 454052 326 454582 354
rect 454470 -960 454582 326
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 16546
rect 461596 480 461624 16546
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462332 354 462360 39374
rect 463712 16574 463740 39442
rect 463712 16546 464016 16574
rect 463988 480 464016 16546
rect 464356 3058 464384 51070
rect 464344 3052 464396 3058
rect 464344 2994 464396 3000
rect 465184 480 465212 78367
rect 471978 78160 472034 78169
rect 471978 78095 472034 78104
rect 466458 47696 466514 47705
rect 466458 47631 466514 47640
rect 466472 16574 466500 47631
rect 468484 47592 468536 47598
rect 468484 47534 468536 47540
rect 466472 16546 467512 16574
rect 466276 3052 466328 3058
rect 466276 2994 466328 3000
rect 466288 480 466316 2994
rect 467484 480 467512 16546
rect 468496 3602 468524 47534
rect 470600 38072 470652 38078
rect 470600 38014 470652 38020
rect 468300 3596 468352 3602
rect 468300 3538 468352 3544
rect 468484 3596 468536 3602
rect 468484 3538 468536 3544
rect 469864 3596 469916 3602
rect 469864 3538 469916 3544
rect 462750 354 462862 480
rect 462332 326 462862 354
rect 462750 -960 462862 326
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468312 354 468340 3538
rect 469876 480 469904 3538
rect 468638 354 468750 480
rect 468312 326 468750 354
rect 468638 -960 468750 326
rect 469834 -960 469946 480
rect 470612 354 470640 38014
rect 471992 16574 472020 78095
rect 478142 71496 478198 71505
rect 478142 71431 478198 71440
rect 472624 64184 472676 64190
rect 472624 64126 472676 64132
rect 471992 16546 472296 16574
rect 472268 480 472296 16546
rect 472636 3534 472664 64126
rect 473450 57352 473506 57361
rect 473450 57287 473506 57296
rect 473464 16574 473492 57287
rect 476120 38004 476172 38010
rect 476120 37946 476172 37952
rect 474740 29776 474792 29782
rect 474740 29718 474792 29724
rect 474752 16574 474780 29718
rect 476132 16574 476160 37946
rect 477500 17332 477552 17338
rect 477500 17274 477552 17280
rect 473464 16546 474136 16574
rect 474752 16546 475792 16574
rect 476132 16546 476528 16574
rect 472624 3528 472676 3534
rect 472624 3470 472676 3476
rect 473452 3528 473504 3534
rect 473452 3470 473504 3476
rect 473464 480 473492 3470
rect 471030 354 471142 480
rect 470612 326 471142 354
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474108 354 474136 16546
rect 475764 480 475792 16546
rect 474526 354 474638 480
rect 474108 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476500 354 476528 16546
rect 477512 6914 477540 17274
rect 478156 16574 478184 71431
rect 480272 16574 480300 78746
rect 483020 78736 483072 78742
rect 483020 78678 483072 78684
rect 482282 75440 482338 75449
rect 482282 75375 482338 75384
rect 481640 36644 481692 36650
rect 481640 36586 481692 36592
rect 481652 16574 481680 36586
rect 478156 16546 478276 16574
rect 480272 16546 480576 16574
rect 481652 16546 481772 16574
rect 477512 6886 478184 6914
rect 478156 480 478184 6886
rect 478248 3602 478276 16546
rect 478236 3596 478288 3602
rect 478236 3538 478288 3544
rect 479340 3528 479392 3534
rect 479340 3470 479392 3476
rect 479352 480 479380 3470
rect 480548 480 480576 16546
rect 481744 480 481772 16546
rect 482192 13116 482244 13122
rect 482192 13058 482244 13064
rect 482204 490 482232 13058
rect 482296 3534 482324 75375
rect 483032 16574 483060 78678
rect 500960 77308 501012 77314
rect 500960 77250 501012 77256
rect 498842 71360 498898 71369
rect 498842 71295 498898 71304
rect 494058 66872 494114 66881
rect 494058 66807 494114 66816
rect 486422 65512 486478 65521
rect 486422 65447 486478 65456
rect 484400 56636 484452 56642
rect 484400 56578 484452 56584
rect 484412 16574 484440 56578
rect 486436 16574 486464 65447
rect 490010 47560 490066 47569
rect 490010 47495 490066 47504
rect 488540 33856 488592 33862
rect 488540 33798 488592 33804
rect 488552 16574 488580 33798
rect 490024 16574 490052 47495
rect 491300 40860 491352 40866
rect 491300 40802 491352 40808
rect 491312 16574 491340 40802
rect 492680 32428 492732 32434
rect 492680 32370 492732 32376
rect 492692 16574 492720 32370
rect 494072 16574 494100 66807
rect 495440 42152 495492 42158
rect 495440 42094 495492 42100
rect 483032 16546 484072 16574
rect 484412 16546 484808 16574
rect 486436 16546 486556 16574
rect 488552 16546 488856 16574
rect 490024 16546 490696 16574
rect 491312 16546 492352 16574
rect 492692 16546 493088 16574
rect 494072 16546 494744 16574
rect 482284 3528 482336 3534
rect 482284 3470 482336 3476
rect 476918 354 477030 480
rect 476500 326 477030 354
rect 476918 -960 477030 326
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482204 462 482416 490
rect 484044 480 484072 16546
rect 482388 354 482416 462
rect 482806 354 482918 480
rect 482388 326 482918 354
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 484780 354 484808 16546
rect 486424 14476 486476 14482
rect 486424 14418 486476 14424
rect 486436 480 486464 14418
rect 486528 4146 486556 16546
rect 486516 4140 486568 4146
rect 486516 4082 486568 4088
rect 487620 3460 487672 3466
rect 487620 3402 487672 3408
rect 487632 480 487660 3402
rect 488828 480 488856 16546
rect 489920 4140 489972 4146
rect 489920 4082 489972 4088
rect 489932 480 489960 4082
rect 485198 354 485310 480
rect 484780 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490668 354 490696 16546
rect 492324 480 492352 16546
rect 491086 354 491198 480
rect 490668 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493060 354 493088 16546
rect 494716 480 494744 16546
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495452 354 495480 42094
rect 498292 40792 498344 40798
rect 498292 40734 498344 40740
rect 498304 16574 498332 40734
rect 498304 16546 498792 16574
rect 497096 3732 497148 3738
rect 497096 3674 497148 3680
rect 497108 480 497136 3674
rect 498200 3596 498252 3602
rect 498200 3538 498252 3544
rect 498212 480 498240 3538
rect 498764 490 498792 16546
rect 498856 3466 498884 71295
rect 499578 55856 499634 55865
rect 499578 55791 499634 55800
rect 499592 16574 499620 55791
rect 500972 16574 501000 77250
rect 509882 75304 509938 75313
rect 509882 75239 509938 75248
rect 507860 67720 507912 67726
rect 507860 67662 507912 67668
rect 502984 49020 503036 49026
rect 502984 48962 503036 48968
rect 502340 29708 502392 29714
rect 502340 29650 502392 29656
rect 499592 16546 500632 16574
rect 500972 16546 501368 16574
rect 498844 3460 498896 3466
rect 498844 3402 498896 3408
rect 495870 354 495982 480
rect 495452 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 498764 462 498976 490
rect 500604 480 500632 16546
rect 498948 354 498976 462
rect 499366 354 499478 480
rect 498948 326 499478 354
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 501340 354 501368 16546
rect 502352 6914 502380 29650
rect 502996 16574 503024 48962
rect 503720 42084 503772 42090
rect 503720 42026 503772 42032
rect 502996 16546 503116 16574
rect 502352 6886 503024 6914
rect 502996 480 503024 6886
rect 503088 3058 503116 16546
rect 503076 3052 503128 3058
rect 503076 2994 503128 3000
rect 501758 354 501870 480
rect 501340 326 501870 354
rect 501758 -960 501870 326
rect 502954 -960 503066 480
rect 503732 354 503760 42026
rect 506572 28280 506624 28286
rect 506572 28222 506624 28228
rect 506584 6914 506612 28222
rect 507872 16574 507900 67662
rect 509240 26988 509292 26994
rect 509240 26930 509292 26936
rect 509252 16574 509280 26930
rect 507872 16546 508912 16574
rect 509252 16546 509648 16574
rect 506492 6886 506612 6914
rect 505376 3052 505428 3058
rect 505376 2994 505428 3000
rect 505388 480 505416 2994
rect 506492 480 506520 6886
rect 507676 3528 507728 3534
rect 507676 3470 507728 3476
rect 507688 480 507716 3470
rect 508884 480 508912 16546
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 509620 354 509648 16546
rect 509896 2990 509924 75239
rect 521660 75200 521712 75206
rect 521660 75142 521712 75148
rect 512000 63572 512052 63578
rect 512000 63514 512052 63520
rect 510620 26920 510672 26926
rect 510620 26862 510672 26868
rect 510632 16574 510660 26862
rect 510632 16546 511304 16574
rect 509884 2984 509936 2990
rect 509884 2926 509936 2932
rect 511276 480 511304 16546
rect 510038 354 510150 480
rect 509620 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512012 354 512040 63514
rect 514022 58576 514078 58585
rect 514022 58511 514078 58520
rect 513380 25628 513432 25634
rect 513380 25570 513432 25576
rect 512430 354 512542 480
rect 512012 326 512542 354
rect 513392 354 513420 25570
rect 514036 3058 514064 58511
rect 516784 53100 516836 53106
rect 516784 53042 516836 53048
rect 516140 39364 516192 39370
rect 516140 39306 516192 39312
rect 516152 16574 516180 39306
rect 516152 16546 516732 16574
rect 516704 3482 516732 16546
rect 516796 3602 516824 53042
rect 520922 44976 520978 44985
rect 520922 44911 520978 44920
rect 520280 24200 520332 24206
rect 520280 24142 520332 24148
rect 518900 17264 518952 17270
rect 518900 17206 518952 17212
rect 518912 16574 518940 17206
rect 518912 16546 519584 16574
rect 516784 3596 516836 3602
rect 516784 3538 516836 3544
rect 518348 3596 518400 3602
rect 518348 3538 518400 3544
rect 516704 3454 517192 3482
rect 514024 3052 514076 3058
rect 514024 2994 514076 3000
rect 515956 3052 516008 3058
rect 515956 2994 516008 3000
rect 514760 2984 514812 2990
rect 514760 2926 514812 2932
rect 514772 480 514800 2926
rect 515968 480 515996 2994
rect 517164 480 517192 3454
rect 518360 480 518388 3538
rect 519556 480 519584 16546
rect 513534 354 513646 480
rect 513392 326 513646 354
rect 512430 -960 512542 326
rect 513534 -960 513646 326
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520292 354 520320 24142
rect 520936 3262 520964 44911
rect 520924 3256 520976 3262
rect 520924 3198 520976 3204
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 521672 354 521700 75142
rect 523144 6914 523172 80679
rect 525800 80096 525852 80102
rect 525800 80038 525852 80044
rect 524418 75168 524474 75177
rect 524418 75103 524474 75112
rect 524432 16574 524460 75103
rect 525812 16574 525840 80038
rect 553400 75948 553452 75954
rect 553400 75890 553452 75896
rect 531318 71224 531374 71233
rect 531318 71159 531374 71168
rect 529940 66972 529992 66978
rect 529940 66914 529992 66920
rect 526442 61432 526498 61441
rect 526442 61367 526498 61376
rect 524432 16546 525472 16574
rect 525812 16546 526208 16574
rect 523052 6886 523172 6914
rect 523052 480 523080 6886
rect 524236 3256 524288 3262
rect 524236 3198 524288 3204
rect 524248 480 524276 3198
rect 525444 480 525472 16546
rect 521814 354 521926 480
rect 521672 326 521926 354
rect 520710 -960 520822 326
rect 521814 -960 521926 326
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526180 354 526208 16546
rect 526456 3534 526484 61367
rect 527824 36576 527876 36582
rect 527824 36518 527876 36524
rect 527180 22840 527232 22846
rect 527180 22782 527232 22788
rect 527192 6914 527220 22782
rect 527836 16574 527864 36518
rect 527836 16546 527956 16574
rect 527192 6886 527864 6914
rect 526444 3528 526496 3534
rect 526444 3470 526496 3476
rect 527836 480 527864 6886
rect 527928 4146 527956 16546
rect 527916 4140 527968 4146
rect 527916 4082 527968 4088
rect 529020 4140 529072 4146
rect 529020 4082 529072 4088
rect 529032 480 529060 4082
rect 526598 354 526710 480
rect 526180 326 526710 354
rect 526598 -960 526710 326
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 529952 354 529980 66914
rect 531332 480 531360 71159
rect 548522 71088 548578 71097
rect 548522 71023 548578 71032
rect 536840 67652 536892 67658
rect 536840 67594 536892 67600
rect 535458 44840 535514 44849
rect 535458 44775 535514 44784
rect 534080 37936 534132 37942
rect 534080 37878 534132 37884
rect 531412 25560 531464 25566
rect 531412 25502 531464 25508
rect 531424 16574 531452 25502
rect 534092 16574 534120 37878
rect 535472 16574 535500 44775
rect 536852 16574 536880 67594
rect 545764 66904 545816 66910
rect 545764 66846 545816 66852
rect 543738 64152 543794 64161
rect 543738 64087 543794 64096
rect 540242 62792 540298 62801
rect 540242 62727 540298 62736
rect 538864 35284 538916 35290
rect 538864 35226 538916 35232
rect 531424 16546 532096 16574
rect 534092 16546 534488 16574
rect 535472 16546 536144 16574
rect 536852 16546 537248 16574
rect 530094 354 530206 480
rect 529952 326 530206 354
rect 530094 -960 530206 326
rect 531290 -960 531402 480
rect 532068 354 532096 16546
rect 533712 3528 533764 3534
rect 533712 3470 533764 3476
rect 533724 480 533752 3470
rect 532486 354 532598 480
rect 532068 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534460 354 534488 16546
rect 536116 480 536144 16546
rect 537220 480 537248 16546
rect 538404 7608 538456 7614
rect 538404 7550 538456 7556
rect 538416 480 538444 7550
rect 538876 3534 538904 35226
rect 540256 3534 540284 62727
rect 542358 51776 542414 51785
rect 542358 51711 542414 51720
rect 542372 16574 542400 51711
rect 543752 16574 543780 64087
rect 542372 16546 542768 16574
rect 543752 16546 544424 16574
rect 541992 4820 542044 4826
rect 541992 4762 542044 4768
rect 538864 3528 538916 3534
rect 538864 3470 538916 3476
rect 539600 3528 539652 3534
rect 539600 3470 539652 3476
rect 540244 3528 540296 3534
rect 540244 3470 540296 3476
rect 539612 480 539640 3470
rect 540796 3460 540848 3466
rect 540796 3402 540848 3408
rect 540808 480 540836 3402
rect 542004 480 542032 4762
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 542740 354 542768 16546
rect 544396 480 544424 16546
rect 545488 11756 545540 11762
rect 545488 11698 545540 11704
rect 545500 480 545528 11698
rect 545776 3466 545804 66846
rect 546500 24132 546552 24138
rect 546500 24074 546552 24080
rect 545764 3460 545816 3466
rect 545764 3402 545816 3408
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546512 354 546540 24074
rect 548432 10328 548484 10334
rect 548432 10270 548484 10276
rect 547880 3528 547932 3534
rect 547880 3470 547932 3476
rect 547892 480 547920 3470
rect 548444 490 548472 10270
rect 548536 3194 548564 71023
rect 549260 40724 549312 40730
rect 549260 40666 549312 40672
rect 549272 16574 549300 40666
rect 552018 36544 552074 36553
rect 552018 36479 552074 36488
rect 549272 16546 550312 16574
rect 548524 3188 548576 3194
rect 548524 3130 548576 3136
rect 546654 354 546766 480
rect 546512 326 546766 354
rect 546654 -960 546766 326
rect 547850 -960 547962 480
rect 548444 462 548656 490
rect 550284 480 550312 16546
rect 552032 6914 552060 36479
rect 552664 22772 552716 22778
rect 552664 22714 552716 22720
rect 552676 16574 552704 22714
rect 553412 16574 553440 75890
rect 557538 69592 557594 69601
rect 557538 69527 557594 69536
rect 556158 50280 556214 50289
rect 556158 50215 556214 50224
rect 556172 16574 556200 50215
rect 557552 16574 557580 69527
rect 570604 64932 570656 64938
rect 570604 64874 570656 64880
rect 563704 60784 563756 60790
rect 563704 60726 563756 60732
rect 560944 45620 560996 45626
rect 560944 45562 560996 45568
rect 558920 35216 558972 35222
rect 558920 35158 558972 35164
rect 558932 16574 558960 35158
rect 552676 16546 552796 16574
rect 553412 16546 553808 16574
rect 556172 16546 556936 16574
rect 557552 16546 558592 16574
rect 558932 16546 559328 16574
rect 552032 6886 552704 6914
rect 551468 3188 551520 3194
rect 551468 3130 551520 3136
rect 551480 480 551508 3130
rect 552676 480 552704 6886
rect 552768 3534 552796 16546
rect 552756 3528 552808 3534
rect 552756 3470 552808 3476
rect 553780 480 553808 16546
rect 556160 8968 556212 8974
rect 556160 8910 556212 8916
rect 554964 3460 555016 3466
rect 554964 3402 555016 3408
rect 554976 480 555004 3402
rect 556172 480 556200 8910
rect 548628 354 548656 462
rect 549046 354 549158 480
rect 548628 326 549158 354
rect 549046 -960 549158 326
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 556908 354 556936 16546
rect 558564 480 558592 16546
rect 557326 354 557438 480
rect 556908 326 557438 354
rect 557326 -960 557438 326
rect 558522 -960 558634 480
rect 559300 354 559328 16546
rect 560852 3528 560904 3534
rect 560852 3470 560904 3476
rect 560864 480 560892 3470
rect 560956 3466 560984 45562
rect 561680 31136 561732 31142
rect 561680 31078 561732 31084
rect 561692 16574 561720 31078
rect 561692 16546 562088 16574
rect 560944 3460 560996 3466
rect 560944 3402 560996 3408
rect 562060 480 562088 16546
rect 563244 6248 563296 6254
rect 563244 6190 563296 6196
rect 563256 480 563284 6190
rect 563716 3534 563744 60726
rect 567842 57216 567898 57225
rect 567842 57151 567898 57160
rect 565818 48920 565874 48929
rect 565818 48855 565874 48864
rect 564532 31068 564584 31074
rect 564532 31010 564584 31016
rect 564544 6914 564572 31010
rect 565832 16574 565860 48855
rect 567200 18692 567252 18698
rect 567200 18634 567252 18640
rect 567212 16574 567240 18634
rect 565832 16546 566872 16574
rect 567212 16546 567608 16574
rect 564452 6886 564572 6914
rect 563704 3528 563756 3534
rect 563704 3470 563756 3476
rect 564452 480 564480 6886
rect 565636 3528 565688 3534
rect 565636 3470 565688 3476
rect 565648 480 565676 3470
rect 566844 480 566872 16546
rect 559718 354 559830 480
rect 559300 326 559830 354
rect 559718 -960 559830 326
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567580 354 567608 16546
rect 567856 3534 567884 57151
rect 569960 49768 570012 49774
rect 569960 49710 570012 49716
rect 569972 16574 570000 49710
rect 569972 16546 570368 16574
rect 567844 3528 567896 3534
rect 567844 3470 567896 3476
rect 569132 3528 569184 3534
rect 569132 3470 569184 3476
rect 569144 480 569172 3470
rect 570340 480 570368 16546
rect 570616 3126 570644 64874
rect 571984 53848 572036 53854
rect 571984 53790 572036 53796
rect 571340 18624 571392 18630
rect 571340 18566 571392 18572
rect 570604 3120 570656 3126
rect 570604 3062 570656 3068
rect 567998 354 568110 480
rect 567580 326 568110 354
rect 567998 -960 568110 326
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571352 354 571380 18566
rect 571996 3398 572024 53790
rect 574100 29640 574152 29646
rect 574100 29582 574152 29588
rect 574112 16574 574140 29582
rect 574756 20670 574784 141063
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 579988 86964 580040 86970
rect 579988 86906 580040 86912
rect 580000 86193 580028 86906
rect 579986 86184 580042 86193
rect 579986 86119 580042 86128
rect 579620 73160 579672 73166
rect 579620 73102 579672 73108
rect 579632 73001 579660 73102
rect 579618 72992 579674 73001
rect 579618 72927 579674 72936
rect 578240 43444 578292 43450
rect 578240 43386 578292 43392
rect 576860 33788 576912 33794
rect 576860 33730 576912 33736
rect 574744 20664 574796 20670
rect 574744 20606 574796 20612
rect 576872 16574 576900 33730
rect 578252 16574 578280 43386
rect 580172 20664 580224 20670
rect 580172 20606 580224 20612
rect 580184 19825 580212 20606
rect 580170 19816 580226 19825
rect 580170 19751 580226 19760
rect 574112 16546 575152 16574
rect 576872 16546 576992 16574
rect 578252 16546 578648 16574
rect 573916 3460 573968 3466
rect 573916 3402 573968 3408
rect 571984 3392 572036 3398
rect 571984 3334 572036 3340
rect 572720 3120 572772 3126
rect 572720 3062 572772 3068
rect 572732 480 572760 3062
rect 573928 480 573956 3402
rect 575124 480 575152 16546
rect 576308 3392 576360 3398
rect 576308 3334 576360 3340
rect 576320 480 576348 3334
rect 571494 354 571606 480
rect 571352 326 571606 354
rect 571494 -960 571606 326
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 576964 354 576992 16546
rect 578620 480 578648 16546
rect 580276 6633 580304 149058
rect 580354 142216 580410 142225
rect 580354 142151 580410 142160
rect 580368 33153 580396 142151
rect 580460 46345 580488 150418
rect 580540 143608 580592 143614
rect 580540 143550 580592 143556
rect 580552 59673 580580 143550
rect 580814 140992 580870 141001
rect 580814 140927 580870 140936
rect 580630 140856 580686 140865
rect 580630 140791 580686 140800
rect 580644 112849 580672 140791
rect 580828 126041 580856 140927
rect 580814 126032 580870 126041
rect 580814 125967 580870 125976
rect 580630 112840 580686 112849
rect 580630 112775 580686 112784
rect 580998 78024 581054 78033
rect 580998 77959 581054 77968
rect 580538 59664 580594 59673
rect 580538 59599 580594 59608
rect 580446 46336 580502 46345
rect 580446 46271 580502 46280
rect 580354 33144 580410 33153
rect 580354 33079 580410 33088
rect 580262 6624 580318 6633
rect 580262 6559 580318 6568
rect 581012 480 581040 77959
rect 581090 77888 581146 77897
rect 581090 77823 581146 77832
rect 581104 16574 581132 77823
rect 581104 16546 581776 16574
rect 577382 354 577494 480
rect 576964 326 577494 354
rect 577382 -960 577494 326
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 581748 354 581776 16546
rect 583392 6180 583444 6186
rect 583392 6122 583444 6128
rect 583404 480 583432 6122
rect 582166 354 582278 480
rect 581748 326 582278 354
rect 582166 -960 582278 326
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 3146 619112 3202 619168
rect 3238 606056 3294 606112
rect 3330 579944 3386 580000
rect 3422 566888 3478 566944
rect 3422 553832 3478 553888
rect 3422 527856 3478 527912
rect 3422 514820 3478 514856
rect 3422 514800 3424 514820
rect 3424 514800 3476 514820
rect 3476 514800 3478 514820
rect 3054 501744 3110 501800
rect 3422 475632 3478 475688
rect 3146 449520 3202 449576
rect 2870 410488 2926 410544
rect 2778 371340 2834 371376
rect 2778 371320 2780 371340
rect 2780 371320 2832 371340
rect 2832 371320 2834 371340
rect 3146 358400 3202 358456
rect 3330 319232 3386 319288
rect 3054 267144 3110 267200
rect 3514 462576 3570 462632
rect 3514 423544 3570 423600
rect 3514 397468 3516 397488
rect 3516 397468 3568 397488
rect 3568 397468 3570 397488
rect 3514 397432 3570 397468
rect 3514 345344 3570 345400
rect 3514 306176 3570 306232
rect 3514 293120 3570 293176
rect 2778 241032 2834 241088
rect 112534 262248 112590 262304
rect 3514 254088 3570 254144
rect 3514 214920 3570 214976
rect 3422 201864 3478 201920
rect 3422 188808 3478 188864
rect 3514 162832 3570 162888
rect 3146 149776 3202 149832
rect 8942 139440 8998 139496
rect 3238 136720 3294 136776
rect 3054 110608 3110 110664
rect 2778 77832 2834 77888
rect 2870 62736 2926 62792
rect 3514 84632 3570 84688
rect 6918 77968 6974 78024
rect 3514 71576 3570 71632
rect 3514 58520 3570 58576
rect 3514 32408 3570 32464
rect 3422 19352 3478 19408
rect 7562 75112 7618 75168
rect 3422 10240 3478 10296
rect 3422 6432 3478 6488
rect 20718 78104 20774 78160
rect 17222 71032 17278 71088
rect 12438 55800 12494 55856
rect 18602 68176 18658 68232
rect 17958 51720 18014 51776
rect 34518 76472 34574 76528
rect 22742 73752 22798 73808
rect 26238 68312 26294 68368
rect 25502 57160 25558 57216
rect 32402 61376 32458 61432
rect 27710 50224 27766 50280
rect 30378 48864 30434 48920
rect 40038 66816 40094 66872
rect 38658 64096 38714 64152
rect 39302 47504 39358 47560
rect 44270 46144 44326 46200
rect 49698 58520 49754 58576
rect 54482 73888 54538 73944
rect 57242 64232 57298 64288
rect 56598 53080 56654 53136
rect 67638 76608 67694 76664
rect 63498 43424 63554 43480
rect 75182 62872 75238 62928
rect 84198 66952 84254 67008
rect 77298 57296 77354 57352
rect 78678 50360 78734 50416
rect 81438 63008 81494 63064
rect 88338 55936 88394 55992
rect 93122 65456 93178 65512
rect 92478 54440 92534 54496
rect 93950 61512 94006 61568
rect 100298 195336 100354 195392
rect 97998 59880 98054 59936
rect 100206 78920 100262 78976
rect 101678 193976 101734 194032
rect 100390 74160 100446 74216
rect 100390 73752 100446 73808
rect 100666 191256 100722 191312
rect 99470 52400 99526 52456
rect 100574 52400 100630 52456
rect 99470 51720 99526 51776
rect 100758 77016 100814 77072
rect 100758 76472 100814 76528
rect 101402 149640 101458 149696
rect 101494 77016 101550 77072
rect 101862 191664 101918 191720
rect 101770 191528 101826 191584
rect 101402 64640 101458 64696
rect 101402 64096 101458 64152
rect 100758 57704 100814 57760
rect 101770 57704 101826 57760
rect 100758 57160 100814 57216
rect 102046 191392 102102 191448
rect 101954 190984 102010 191040
rect 101862 50224 101918 50280
rect 99470 49544 99526 49600
rect 100666 49544 100722 49600
rect 99470 48864 99526 48920
rect 100758 48184 100814 48240
rect 101954 48184 102010 48240
rect 100758 47504 100814 47560
rect 102782 151000 102838 151056
rect 102138 68312 102194 68368
rect 102230 68176 102286 68232
rect 102690 62056 102746 62112
rect 102138 61376 102194 61432
rect 102138 54576 102194 54632
rect 100758 46824 100814 46880
rect 102046 46824 102102 46880
rect 100758 46144 100814 46200
rect 103242 194248 103298 194304
rect 103150 78512 103206 78568
rect 102230 44104 102286 44160
rect 102782 44104 102838 44160
rect 102230 43424 102286 43480
rect 103058 68856 103114 68912
rect 103978 81912 104034 81968
rect 104530 66816 104586 66872
rect 104714 189624 104770 189680
rect 104254 64640 104310 64696
rect 104254 64232 104310 64288
rect 104162 59220 104218 59256
rect 104162 59200 104164 59220
rect 104164 59200 104216 59220
rect 104216 59200 104218 59220
rect 104162 58520 104218 58576
rect 103794 57840 103850 57896
rect 104714 57840 104770 57896
rect 103794 57296 103850 57352
rect 107198 199144 107254 199200
rect 105450 151272 105506 151328
rect 105358 151136 105414 151192
rect 105358 63416 105414 63472
rect 105910 198192 105966 198248
rect 105634 77968 105690 78024
rect 106922 196832 106978 196888
rect 106002 194112 106058 194168
rect 106094 191120 106150 191176
rect 106094 62056 106150 62112
rect 105450 53760 105506 53816
rect 105450 53080 105506 53136
rect 104806 50904 104862 50960
rect 108210 195472 108266 195528
rect 107474 190032 107530 190088
rect 107198 74024 107254 74080
rect 107382 71052 107438 71088
rect 107382 71032 107384 71052
rect 107384 71032 107436 71052
rect 107436 71032 107438 71052
rect 106922 66136 106978 66192
rect 107566 186904 107622 186960
rect 107474 63144 107530 63200
rect 108118 137808 108174 137864
rect 107566 55120 107622 55176
rect 107566 54576 107622 54632
rect 108302 66952 108358 67008
rect 108946 66136 109002 66192
rect 109590 76880 109646 76936
rect 110142 67496 110198 67552
rect 110970 146920 111026 146976
rect 110878 139032 110934 139088
rect 111430 73072 111486 73128
rect 110326 64640 110382 64696
rect 111706 76608 111762 76664
rect 112534 138624 112590 138680
rect 112442 75248 112498 75304
rect 111614 64504 111670 64560
rect 112258 60580 112314 60616
rect 112258 60560 112260 60580
rect 112260 60560 112312 60580
rect 112312 60560 112314 60580
rect 111798 59880 111854 59936
rect 115110 262384 115166 262440
rect 114006 138896 114062 138952
rect 113546 55936 113602 55992
rect 114098 138352 114154 138408
rect 115294 259664 115350 259720
rect 115018 142024 115074 142080
rect 115018 78648 115074 78704
rect 114098 68448 114154 68504
rect 115294 144064 115350 144120
rect 115754 75384 115810 75440
rect 115846 72936 115902 72992
rect 116858 143928 116914 143984
rect 116490 142160 116546 142216
rect 116490 139848 116546 139904
rect 116398 80824 116454 80880
rect 116490 78784 116546 78840
rect 116674 138080 116730 138136
rect 116674 72800 116730 72856
rect 116950 75248 117006 75304
rect 117778 92384 117834 92440
rect 117870 81096 117926 81152
rect 118422 76744 118478 76800
rect 118790 140664 118846 140720
rect 119434 259800 119490 259856
rect 120814 262656 120870 262712
rect 119434 140528 119490 140584
rect 119342 136584 119398 136640
rect 119526 140120 119582 140176
rect 119526 71304 119582 71360
rect 117686 69672 117742 69728
rect 119986 195744 120042 195800
rect 120446 147600 120502 147656
rect 119894 72664 119950 72720
rect 120078 52536 120134 52592
rect 120814 144472 120870 144528
rect 125598 261160 125654 261216
rect 133970 261024 134026 261080
rect 135902 265240 135958 265296
rect 137466 260888 137522 260944
rect 138662 262792 138718 262848
rect 140778 260072 140834 260128
rect 141422 259936 141478 259992
rect 142618 263880 142674 263936
rect 142250 262520 142306 262576
rect 142894 262520 142950 262576
rect 145010 263064 145066 263120
rect 145010 262248 145066 262304
rect 146206 263744 146262 263800
rect 145654 263064 145710 263120
rect 147034 264968 147090 265024
rect 146942 262384 146998 262440
rect 147678 260208 147734 260264
rect 148506 265104 148562 265160
rect 148368 260208 148424 260264
rect 147678 259800 147734 259856
rect 148138 259664 148194 259720
rect 151818 274624 151874 274680
rect 151082 263608 151138 263664
rect 150530 262656 150586 262712
rect 153658 262384 153714 262440
rect 158810 262656 158866 262712
rect 159914 262656 159970 262712
rect 160098 259936 160154 259992
rect 162030 262520 162086 262576
rect 161478 260752 161534 260808
rect 160926 259936 160982 259992
rect 163502 264968 163558 265024
rect 162674 260752 162730 260808
rect 162582 259800 162638 259856
rect 169022 265240 169078 265296
rect 167550 265104 167606 265160
rect 161202 259664 161258 259720
rect 149242 259528 149298 259584
rect 155222 259528 155278 259584
rect 187698 262928 187754 262984
rect 187698 262384 187754 262440
rect 187974 262384 188030 262440
rect 185674 259528 185730 259584
rect 120998 143112 121054 143168
rect 120630 74568 120686 74624
rect 120998 138488 121054 138544
rect 121182 196696 121238 196752
rect 121734 138080 121790 138136
rect 122010 148008 122066 148064
rect 121826 136584 121882 136640
rect 121734 132504 121790 132560
rect 121826 132368 121882 132424
rect 121826 122848 121882 122904
rect 121826 122712 121882 122768
rect 121826 113192 121882 113248
rect 121826 113056 121882 113112
rect 121826 103536 121882 103592
rect 121826 103400 121882 103456
rect 121826 93880 121882 93936
rect 120446 54984 120502 55040
rect 120446 54440 120502 54496
rect 122378 80960 122434 81016
rect 122562 147736 122618 147792
rect 122746 151544 122802 151600
rect 123574 194520 123630 194576
rect 122746 146648 122802 146704
rect 123574 142840 123630 142896
rect 123390 141888 123446 141944
rect 123390 139712 123446 139768
rect 123942 142160 123998 142216
rect 124586 141888 124642 141944
rect 124586 141072 124642 141128
rect 127714 200640 127770 200696
rect 125230 143248 125286 143304
rect 125598 142060 125600 142080
rect 125600 142060 125652 142080
rect 125652 142060 125654 142080
rect 125598 142024 125654 142060
rect 125138 141888 125194 141944
rect 124862 140256 124918 140312
rect 126518 141208 126574 141264
rect 126978 142296 127034 142352
rect 127070 140800 127126 140856
rect 124494 139576 124550 139632
rect 125506 139576 125562 139632
rect 127898 199008 127954 199064
rect 127806 142296 127862 142352
rect 127714 140528 127770 140584
rect 128082 198872 128138 198928
rect 127898 140664 127954 140720
rect 128358 193840 128414 193896
rect 131486 200504 131542 200560
rect 130106 199960 130162 200016
rect 128450 140936 128506 140992
rect 128082 140392 128138 140448
rect 131578 200096 131634 200152
rect 131762 199552 131818 199608
rect 131578 199416 131634 199472
rect 132130 200504 132186 200560
rect 131946 199824 132002 199880
rect 132222 199552 132278 199608
rect 131854 198736 131910 198792
rect 131762 196968 131818 197024
rect 130566 195200 130622 195256
rect 130106 194384 130162 194440
rect 129830 146240 129886 146296
rect 129094 140392 129150 140448
rect 127530 139576 127586 139632
rect 131026 192480 131082 192536
rect 130658 146784 130714 146840
rect 131854 147328 131910 147384
rect 131118 145424 131174 145480
rect 129462 139576 129518 139632
rect 132130 199416 132186 199472
rect 132314 199416 132370 199472
rect 132038 197920 132094 197976
rect 133004 199824 133060 199880
rect 132958 199724 132960 199744
rect 132960 199724 133012 199744
rect 133012 199724 133014 199744
rect 132958 199688 133014 199724
rect 132498 198328 132554 198384
rect 132406 198192 132462 198248
rect 132958 191528 133014 191584
rect 133234 198056 133290 198112
rect 133648 199858 133704 199914
rect 133510 198600 133566 198656
rect 133326 189896 133382 189952
rect 134752 199824 134808 199880
rect 133786 196288 133842 196344
rect 134338 193976 134394 194032
rect 134614 199436 134670 199472
rect 134614 199416 134616 199436
rect 134616 199416 134668 199436
rect 134668 199416 134670 199436
rect 134522 198600 134578 198656
rect 132222 147464 132278 147520
rect 134890 194248 134946 194304
rect 135580 199824 135636 199880
rect 135258 199416 135314 199472
rect 135258 199144 135314 199200
rect 135258 196152 135314 196208
rect 135350 195880 135406 195936
rect 135534 196016 135590 196072
rect 135442 195608 135498 195664
rect 136408 199858 136464 199914
rect 135902 199144 135958 199200
rect 136362 199144 136418 199200
rect 136868 199858 136924 199914
rect 137144 199858 137200 199914
rect 136546 196832 136602 196888
rect 136730 197104 136786 197160
rect 136822 196832 136878 196888
rect 137512 199858 137568 199914
rect 137190 198736 137246 198792
rect 137282 197240 137338 197296
rect 138340 199858 138396 199914
rect 138524 199858 138580 199914
rect 136178 148960 136234 149016
rect 135718 148824 135774 148880
rect 137466 196832 137522 196888
rect 138800 199858 138856 199914
rect 138110 198464 138166 198520
rect 138294 199144 138350 199200
rect 138662 196832 138718 196888
rect 137466 151408 137522 151464
rect 137098 147192 137154 147248
rect 135810 146104 135866 146160
rect 139260 199858 139316 199914
rect 139536 199858 139592 199914
rect 139904 199858 139960 199914
rect 140088 199858 140144 199914
rect 139398 199688 139454 199744
rect 138754 194112 138810 194168
rect 140042 199688 140098 199744
rect 139398 199144 139454 199200
rect 139766 197240 139822 197296
rect 138570 187176 138626 187232
rect 138478 151680 138534 151736
rect 140640 199824 140696 199880
rect 140916 199858 140972 199914
rect 141192 199858 141248 199914
rect 141560 199858 141616 199914
rect 140502 199688 140558 199744
rect 138662 144608 138718 144664
rect 139950 187040 140006 187096
rect 140962 199688 141018 199744
rect 141146 199416 141202 199472
rect 141238 198736 141294 198792
rect 140870 198192 140926 198248
rect 140962 198056 141018 198112
rect 140226 195744 140282 195800
rect 141422 198736 141478 198792
rect 141606 199416 141662 199472
rect 141790 199552 141846 199608
rect 141882 198736 141938 198792
rect 141882 195472 141938 195528
rect 142066 198736 142122 198792
rect 142664 199858 142720 199914
rect 142618 199416 142674 199472
rect 142434 195880 142490 195936
rect 142250 194248 142306 194304
rect 141054 151544 141110 151600
rect 140870 149776 140926 149832
rect 140042 141616 140098 141672
rect 139858 140256 139914 140312
rect 143124 199858 143180 199914
rect 143400 199858 143456 199914
rect 143032 199688 143088 199744
rect 144044 199858 144100 199914
rect 144228 199858 144284 199914
rect 145148 199858 145204 199914
rect 143354 199552 143410 199608
rect 143078 199416 143134 199472
rect 143078 198736 143134 198792
rect 143170 196832 143226 196888
rect 143814 199452 143816 199472
rect 143816 199452 143868 199472
rect 143868 199452 143870 199472
rect 143814 199416 143870 199452
rect 143998 199552 144054 199608
rect 143814 196424 143870 196480
rect 144182 199552 144238 199608
rect 144642 194384 144698 194440
rect 145102 199688 145158 199744
rect 145516 199858 145572 199914
rect 145470 199416 145526 199472
rect 145102 196832 145158 196888
rect 142526 144336 142582 144392
rect 143078 142976 143134 143032
rect 145838 199552 145894 199608
rect 146528 199858 146584 199914
rect 146712 199858 146768 199914
rect 146896 199858 146952 199914
rect 146850 199688 146906 199744
rect 147264 199858 147320 199914
rect 147448 199858 147504 199914
rect 147632 199858 147688 199914
rect 147034 199144 147090 199200
rect 147908 199858 147964 199914
rect 147402 196560 147458 196616
rect 147908 199722 147964 199778
rect 147678 199552 147734 199608
rect 147770 199416 147826 199472
rect 147862 198056 147918 198112
rect 148552 199858 148608 199914
rect 148736 199858 148792 199914
rect 148690 199688 148746 199744
rect 148506 199552 148562 199608
rect 147770 145560 147826 145616
rect 147678 144472 147734 144528
rect 149380 199858 149436 199914
rect 149564 199858 149620 199914
rect 149334 199552 149390 199608
rect 149518 199552 149574 199608
rect 150116 199858 150172 199914
rect 150392 199824 150448 199880
rect 150760 199858 150816 199914
rect 151496 199824 151552 199880
rect 149702 199416 149758 199472
rect 148874 194520 148930 194576
rect 149978 199552 150034 199608
rect 149702 195608 149758 195664
rect 149242 148552 149298 148608
rect 148598 148280 148654 148336
rect 149058 145832 149114 145888
rect 148598 144064 148654 144120
rect 150622 199688 150678 199744
rect 151956 199858 152012 199914
rect 151082 199280 151138 199336
rect 151174 196832 151230 196888
rect 151450 196560 151506 196616
rect 151726 148280 151782 148336
rect 153244 199858 153300 199914
rect 153520 199858 153576 199914
rect 153796 199858 153852 199914
rect 152646 199144 152702 199200
rect 152462 196968 152518 197024
rect 152738 192616 152794 192672
rect 153106 199552 153162 199608
rect 153198 196832 153254 196888
rect 153474 199552 153530 199608
rect 153658 198872 153714 198928
rect 153474 198056 153530 198112
rect 153566 197920 153622 197976
rect 152002 148416 152058 148472
rect 151910 148144 151966 148200
rect 151358 142704 151414 142760
rect 153750 195880 153806 195936
rect 154118 199688 154174 199744
rect 154532 199858 154588 199914
rect 153934 199552 153990 199608
rect 154532 199640 154588 199642
rect 154532 199588 154534 199640
rect 154534 199588 154586 199640
rect 154586 199588 154588 199640
rect 154900 199858 154956 199914
rect 154532 199586 154588 199588
rect 154302 195608 154358 195664
rect 154210 195336 154266 195392
rect 153842 192480 153898 192536
rect 153658 151272 153714 151328
rect 153566 148688 153622 148744
rect 153474 145696 153530 145752
rect 153290 141480 153346 141536
rect 154578 199416 154634 199472
rect 155452 199858 155508 199914
rect 155406 199688 155462 199744
rect 155728 199824 155784 199880
rect 155912 199858 155968 199914
rect 156096 199858 156152 199914
rect 155958 199688 156014 199744
rect 155590 199588 155592 199608
rect 155592 199588 155644 199608
rect 155644 199588 155646 199608
rect 155590 199552 155646 199588
rect 154026 141344 154082 141400
rect 155774 199552 155830 199608
rect 156142 199688 156198 199744
rect 156648 199858 156704 199914
rect 155958 199008 156014 199064
rect 156464 199688 156520 199744
rect 156602 199688 156658 199744
rect 156832 199722 156888 199778
rect 157108 199858 157164 199914
rect 156418 199416 156474 199472
rect 156786 199552 156842 199608
rect 157200 199722 157256 199778
rect 157752 199858 157808 199914
rect 157154 198872 157210 198928
rect 157522 199552 157578 199608
rect 157154 196832 157210 196888
rect 156142 144200 156198 144256
rect 157338 196560 157394 196616
rect 158028 199688 158084 199744
rect 158442 199688 158498 199744
rect 157982 199552 158038 199608
rect 157798 199028 157854 199064
rect 157798 199008 157800 199028
rect 157800 199008 157852 199028
rect 157852 199008 157854 199028
rect 157890 196560 157946 196616
rect 159500 199858 159556 199914
rect 158994 199552 159050 199608
rect 158626 198192 158682 198248
rect 158534 196016 158590 196072
rect 158994 199416 159050 199472
rect 158810 195336 158866 195392
rect 157338 142024 157394 142080
rect 157154 141344 157210 141400
rect 157890 148552 157946 148608
rect 159868 199858 159924 199914
rect 159546 198484 159602 198520
rect 159546 198464 159548 198484
rect 159548 198464 159600 198484
rect 159600 198464 159602 198484
rect 160328 199858 160384 199914
rect 160512 199858 160568 199914
rect 160788 199858 160844 199914
rect 160282 199552 160338 199608
rect 160834 199688 160890 199744
rect 161340 199858 161396 199914
rect 161616 199858 161672 199914
rect 161478 199776 161534 199778
rect 160466 199552 160522 199608
rect 160650 197240 160706 197296
rect 161018 199552 161074 199608
rect 161202 199724 161204 199744
rect 161204 199724 161256 199744
rect 161256 199724 161258 199744
rect 161202 199688 161258 199724
rect 161478 199724 161480 199776
rect 161480 199724 161532 199776
rect 161532 199724 161534 199776
rect 161478 199722 161534 199724
rect 161110 196696 161166 196752
rect 161202 196424 161258 196480
rect 161570 199416 161626 199472
rect 162076 199858 162132 199914
rect 162260 199858 162316 199914
rect 161754 196016 161810 196072
rect 161570 195744 161626 195800
rect 161478 195336 161534 195392
rect 162214 199688 162270 199744
rect 162030 195608 162086 195664
rect 162214 196696 162270 196752
rect 162904 199858 162960 199914
rect 162398 199552 162454 199608
rect 162398 199144 162454 199200
rect 162490 197784 162546 197840
rect 162398 196832 162454 196888
rect 162950 199552 163006 199608
rect 162582 195472 162638 195528
rect 163456 199858 163512 199914
rect 163502 199688 163558 199744
rect 163640 199722 163696 199778
rect 164100 199858 164156 199914
rect 164376 199858 164432 199914
rect 163686 199416 163742 199472
rect 163686 199300 163742 199336
rect 163686 199280 163688 199300
rect 163688 199280 163740 199300
rect 163740 199280 163742 199300
rect 163594 199008 163650 199064
rect 163594 196832 163650 196888
rect 163318 196424 163374 196480
rect 162490 144336 162546 144392
rect 160834 144064 160890 144120
rect 159638 142840 159694 142896
rect 161938 142704 161994 142760
rect 163410 196288 163466 196344
rect 163962 199572 164018 199608
rect 163962 199552 163964 199572
rect 163964 199552 164016 199572
rect 164016 199552 164018 199572
rect 163962 199280 164018 199336
rect 164606 199688 164662 199744
rect 164330 199144 164386 199200
rect 164330 197512 164386 197568
rect 164238 197104 164294 197160
rect 164146 196832 164202 196888
rect 164514 199552 164570 199608
rect 165204 199858 165260 199914
rect 164882 199688 164938 199744
rect 165158 199688 165214 199744
rect 164606 199008 164662 199064
rect 163042 145560 163098 145616
rect 163594 142840 163650 142896
rect 162582 139848 162638 139904
rect 165572 199858 165628 199914
rect 165250 199416 165306 199472
rect 165158 197240 165214 197296
rect 164974 196424 165030 196480
rect 165756 199688 165812 199744
rect 166032 199858 166088 199914
rect 165894 199416 165950 199472
rect 166308 199858 166364 199914
rect 167136 199858 167192 199914
rect 166078 199280 166134 199336
rect 166262 198872 166318 198928
rect 166078 196288 166134 196344
rect 166262 195744 166318 195800
rect 166630 196968 166686 197024
rect 166952 199688 167008 199744
rect 167090 199416 167146 199472
rect 166906 198736 166962 198792
rect 164330 144608 164386 144664
rect 165250 142976 165306 143032
rect 164606 139712 164662 139768
rect 167872 199858 167928 199914
rect 168056 199858 168112 199914
rect 168332 199858 168388 199914
rect 167826 199552 167882 199608
rect 167642 196152 167698 196208
rect 168976 199858 169032 199914
rect 169160 199858 169216 199914
rect 168608 199688 168664 199744
rect 168746 199688 168802 199744
rect 169712 199858 169768 199914
rect 168010 199552 168066 199608
rect 167918 195744 167974 195800
rect 167734 194520 167790 194576
rect 168470 199552 168526 199608
rect 168378 198328 168434 198384
rect 168286 196424 168342 196480
rect 168010 193160 168066 193216
rect 168746 199552 168802 199608
rect 168654 199416 168710 199472
rect 168654 199280 168710 199336
rect 168378 192208 168434 192264
rect 167182 151408 167238 151464
rect 167090 149504 167146 149560
rect 166998 148416 167054 148472
rect 168010 144472 168066 144528
rect 168838 195200 168894 195256
rect 169114 199588 169116 199608
rect 169116 199588 169168 199608
rect 169168 199588 169170 199608
rect 169114 199552 169170 199588
rect 169206 199280 169262 199336
rect 169712 199688 169768 199744
rect 169114 196424 169170 196480
rect 169022 196288 169078 196344
rect 168746 193296 168802 193352
rect 169390 196016 169446 196072
rect 168562 191120 168618 191176
rect 169666 199552 169722 199608
rect 169896 199858 169952 199914
rect 170080 199858 170136 199914
rect 170264 199858 170320 199914
rect 169574 196424 169630 196480
rect 169758 199008 169814 199064
rect 169942 199452 169944 199472
rect 169944 199452 169996 199472
rect 169996 199452 169998 199472
rect 169942 199416 169998 199452
rect 169850 196288 169906 196344
rect 169758 196152 169814 196208
rect 169758 193024 169814 193080
rect 170126 199552 170182 199608
rect 170126 196152 170182 196208
rect 170034 192072 170090 192128
rect 169942 147328 169998 147384
rect 170126 147192 170182 147248
rect 169758 139984 169814 140040
rect 170632 199858 170688 199914
rect 170908 199790 170964 199846
rect 171276 199858 171332 199914
rect 171230 199688 171286 199744
rect 171920 199858 171976 199914
rect 170678 199552 170734 199608
rect 170586 198192 170642 198248
rect 170310 147600 170366 147656
rect 170954 199416 171010 199472
rect 170862 198636 170864 198656
rect 170864 198636 170916 198656
rect 170916 198636 170918 198656
rect 170862 198600 170918 198636
rect 171230 198328 171286 198384
rect 171046 198056 171102 198112
rect 171322 197512 171378 197568
rect 171322 196424 171378 196480
rect 171598 197784 171654 197840
rect 171598 196016 171654 196072
rect 171138 147464 171194 147520
rect 172058 199688 172114 199744
rect 172196 199688 172252 199744
rect 172656 199858 172712 199914
rect 172932 199824 172988 199880
rect 172610 199688 172666 199744
rect 171782 197376 171838 197432
rect 171322 147056 171378 147112
rect 172242 198736 172298 198792
rect 172150 197920 172206 197976
rect 172058 196424 172114 196480
rect 173208 199824 173264 199880
rect 172610 197920 172666 197976
rect 173668 199824 173724 199880
rect 173070 198872 173126 198928
rect 173254 198328 173310 198384
rect 172794 197376 172850 197432
rect 172518 196288 172574 196344
rect 171782 145696 171838 145752
rect 172702 196288 172758 196344
rect 173162 196152 173218 196208
rect 174404 199858 174460 199914
rect 174588 199858 174644 199914
rect 173438 194384 173494 194440
rect 173622 193976 173678 194032
rect 172518 145968 172574 146024
rect 174266 199280 174322 199336
rect 174174 199008 174230 199064
rect 174174 198872 174230 198928
rect 174542 199708 174598 199744
rect 174542 199688 174544 199708
rect 174544 199688 174596 199708
rect 174596 199688 174598 199708
rect 174634 199280 174690 199336
rect 174634 194384 174690 194440
rect 174542 194248 174598 194304
rect 175232 199858 175288 199914
rect 175876 199858 175932 199914
rect 174174 150320 174230 150376
rect 175370 198464 175426 198520
rect 175186 197648 175242 197704
rect 174542 192072 174598 192128
rect 174358 150048 174414 150104
rect 173898 145832 173954 145888
rect 175462 197376 175518 197432
rect 175922 199144 175978 199200
rect 176014 198736 176070 198792
rect 176428 199858 176484 199914
rect 175922 193024 175978 193080
rect 175922 192208 175978 192264
rect 175646 189760 175702 189816
rect 175462 149640 175518 149696
rect 177072 199824 177128 199880
rect 177946 199588 177948 199608
rect 177948 199588 178000 199608
rect 178000 199588 178002 199608
rect 177946 199552 178002 199588
rect 177670 195064 177726 195120
rect 177118 189896 177174 189952
rect 176658 149776 176714 149832
rect 178222 199824 178278 199880
rect 176474 146104 176530 146160
rect 174542 141480 174598 141536
rect 179050 199688 179106 199744
rect 179050 199008 179106 199064
rect 180154 200504 180210 200560
rect 179418 146784 179474 146840
rect 180338 200368 180394 200424
rect 180338 144744 180394 144800
rect 182270 193840 182326 193896
rect 182822 140528 182878 140584
rect 183006 140256 183062 140312
rect 183834 194792 183890 194848
rect 183190 140392 183246 140448
rect 181258 139440 181314 139496
rect 185398 143112 185454 143168
rect 185398 142432 185454 142488
rect 185858 150456 185914 150512
rect 185674 143384 185730 143440
rect 185674 142568 185730 142624
rect 186042 152360 186098 152416
rect 123114 139304 123170 139360
rect 123850 139304 123906 139360
rect 129186 139304 129242 139360
rect 131946 139304 132002 139360
rect 166722 139304 166778 139360
rect 173438 139304 173494 139360
rect 184110 139304 184166 139360
rect 184386 139304 184442 139360
rect 185490 139304 185546 139360
rect 186502 140120 186558 140176
rect 186226 139304 186282 139360
rect 124126 78240 124182 78296
rect 130014 80552 130070 80608
rect 129738 80144 129794 80200
rect 128542 79872 128598 79928
rect 129002 78512 129058 78568
rect 128542 78376 128598 78432
rect 126978 77832 127034 77888
rect 129646 77832 129702 77888
rect 129554 77560 129610 77616
rect 129002 75112 129058 75168
rect 178038 80552 178094 80608
rect 130014 77288 130070 77344
rect 130474 75248 130530 75304
rect 129922 75112 129978 75168
rect 130842 77968 130898 78024
rect 130842 77288 130898 77344
rect 130934 75248 130990 75304
rect 132038 75792 132094 75848
rect 132636 79872 132692 79928
rect 133188 79906 133244 79962
rect 133556 79906 133612 79962
rect 132866 79756 132922 79792
rect 132866 79736 132868 79756
rect 132868 79736 132920 79756
rect 132920 79736 132922 79756
rect 133234 79736 133290 79792
rect 133418 79736 133474 79792
rect 134200 79906 134256 79962
rect 134752 79838 134808 79894
rect 132498 78240 132554 78296
rect 133050 79600 133106 79656
rect 133234 79600 133290 79656
rect 133326 77696 133382 77752
rect 134154 78512 134210 78568
rect 134154 78376 134210 78432
rect 134062 77288 134118 77344
rect 133970 76608 134026 76664
rect 134430 78920 134486 78976
rect 134338 78240 134394 78296
rect 134522 77852 134578 77888
rect 134522 77832 134524 77852
rect 134524 77832 134576 77852
rect 134576 77832 134578 77852
rect 134936 79906 134992 79962
rect 134706 77016 134762 77072
rect 135304 79872 135360 79928
rect 135672 79906 135728 79962
rect 135948 79906 136004 79962
rect 134982 79600 135038 79656
rect 135350 77288 135406 77344
rect 135534 79464 135590 79520
rect 135994 79736 136050 79792
rect 135810 77560 135866 77616
rect 136500 79906 136556 79962
rect 136454 79600 136510 79656
rect 136270 79464 136326 79520
rect 137052 79872 137108 79928
rect 137328 79906 137384 79962
rect 137006 79736 137062 79792
rect 136914 79600 136970 79656
rect 136730 78240 136786 78296
rect 136914 65728 136970 65784
rect 137282 79600 137338 79656
rect 137696 79736 137752 79792
rect 137880 79838 137936 79894
rect 137558 79464 137614 79520
rect 137926 78512 137982 78568
rect 138340 79736 138396 79792
rect 138524 79872 138580 79928
rect 138570 79772 138572 79792
rect 138572 79772 138624 79792
rect 138624 79772 138626 79792
rect 138570 79736 138626 79772
rect 138984 79906 139040 79962
rect 139168 79838 139224 79894
rect 139444 79872 139500 79928
rect 139720 79906 139776 79962
rect 140272 79906 140328 79962
rect 138110 66000 138166 66056
rect 138938 77968 138994 78024
rect 139214 79600 139270 79656
rect 139490 79328 139546 79384
rect 139674 79600 139730 79656
rect 139582 78512 139638 78568
rect 138478 66000 138534 66056
rect 139582 65592 139638 65648
rect 140226 79600 140282 79656
rect 140502 77832 140558 77888
rect 140824 79906 140880 79962
rect 141376 79872 141432 79928
rect 140962 76880 141018 76936
rect 140226 65592 140282 65648
rect 141422 78240 141478 78296
rect 141422 77832 141478 77888
rect 142296 79838 142352 79894
rect 142664 79872 142720 79928
rect 141698 78104 141754 78160
rect 142250 79328 142306 79384
rect 142158 77832 142214 77888
rect 142342 77424 142398 77480
rect 143216 79838 143272 79894
rect 143584 79872 143640 79928
rect 142710 68720 142766 68776
rect 142710 68040 142766 68096
rect 143446 79600 143502 79656
rect 143768 79770 143824 79826
rect 143952 79736 144008 79792
rect 143538 78920 143594 78976
rect 144274 79600 144330 79656
rect 144366 79328 144422 79384
rect 144826 79736 144882 79792
rect 145056 79906 145112 79962
rect 145240 79906 145296 79962
rect 144550 79636 144552 79656
rect 144552 79636 144604 79656
rect 144604 79636 144606 79656
rect 144550 79600 144606 79636
rect 144550 79464 144606 79520
rect 144458 77968 144514 78024
rect 144734 79464 144790 79520
rect 144182 74976 144238 75032
rect 144642 77832 144698 77888
rect 145102 79464 145158 79520
rect 145976 79906 146032 79962
rect 146160 79906 146216 79962
rect 146712 79906 146768 79962
rect 145930 79736 145986 79792
rect 146114 79464 146170 79520
rect 146206 76608 146262 76664
rect 146666 79600 146722 79656
rect 147264 79872 147320 79928
rect 147632 79772 147634 79792
rect 147634 79772 147686 79792
rect 147686 79772 147688 79792
rect 147632 79736 147688 79772
rect 147816 79906 147872 79962
rect 148184 79906 148240 79962
rect 147218 79620 147274 79656
rect 147218 79600 147220 79620
rect 147220 79600 147272 79620
rect 147272 79600 147274 79620
rect 147034 77424 147090 77480
rect 147126 67632 147182 67688
rect 147678 79600 147734 79656
rect 147862 79464 147918 79520
rect 147862 79328 147918 79384
rect 147586 77288 147642 77344
rect 148138 79328 148194 79384
rect 148552 79872 148608 79928
rect 148736 79906 148792 79962
rect 148414 79600 148470 79656
rect 149196 79872 149252 79928
rect 148690 79464 148746 79520
rect 148598 77424 148654 77480
rect 148506 69400 148562 69456
rect 149058 78512 149114 78568
rect 150576 79906 150632 79962
rect 150760 79838 150816 79894
rect 149334 78648 149390 78704
rect 148966 77560 149022 77616
rect 148874 77288 148930 77344
rect 148874 70080 148930 70136
rect 148874 69400 148930 69456
rect 149150 74024 149206 74080
rect 150070 79600 150126 79656
rect 149610 77288 149666 77344
rect 149518 71168 149574 71224
rect 150070 77288 150126 77344
rect 150254 79600 150310 79656
rect 150438 78512 150494 78568
rect 150346 77424 150402 77480
rect 149702 67496 149758 67552
rect 150346 71576 150402 71632
rect 150806 79464 150862 79520
rect 150714 77424 150770 77480
rect 151082 78104 151138 78160
rect 151266 79600 151322 79656
rect 151266 78784 151322 78840
rect 151174 73888 151230 73944
rect 151174 71712 151230 71768
rect 151450 79600 151506 79656
rect 151358 71712 151414 71768
rect 151864 79736 151920 79792
rect 151542 76472 151598 76528
rect 152278 79736 152334 79792
rect 152002 76744 152058 76800
rect 151726 74432 151782 74488
rect 151174 68584 151230 68640
rect 152692 79872 152748 79928
rect 152600 79772 152602 79792
rect 152602 79772 152654 79792
rect 152654 79772 152656 79792
rect 152600 79736 152656 79772
rect 152002 68856 152058 68912
rect 152738 77424 152794 77480
rect 154072 79906 154128 79962
rect 153290 79736 153346 79792
rect 152830 69808 152886 69864
rect 152738 68856 152794 68912
rect 153014 70488 153070 70544
rect 153290 79192 153346 79248
rect 153474 79600 153530 79656
rect 153474 73480 153530 73536
rect 153658 79636 153660 79656
rect 153660 79636 153712 79656
rect 153712 79636 153714 79656
rect 153658 79600 153714 79636
rect 153842 79600 153898 79656
rect 153382 68040 153438 68096
rect 153934 79328 153990 79384
rect 154440 79906 154496 79962
rect 154302 79736 154358 79792
rect 154394 79600 154450 79656
rect 154210 79464 154266 79520
rect 154302 77152 154358 77208
rect 154118 75520 154174 75576
rect 153658 69944 153714 70000
rect 154026 69944 154082 70000
rect 153934 68040 153990 68096
rect 154992 79906 155048 79962
rect 155268 79906 155324 79962
rect 154808 79824 154864 79826
rect 154808 79772 154810 79824
rect 154810 79772 154862 79824
rect 154862 79772 154864 79824
rect 154808 79770 154864 79772
rect 154486 76336 154542 76392
rect 155544 79872 155600 79928
rect 155912 79906 155968 79962
rect 154394 74296 154450 74352
rect 154854 78104 154910 78160
rect 154854 66136 154910 66192
rect 156096 79906 156152 79962
rect 156280 79906 156336 79962
rect 156740 79906 156796 79962
rect 155682 79600 155738 79656
rect 156050 79192 156106 79248
rect 155958 77968 156014 78024
rect 155498 71440 155554 71496
rect 156418 79600 156474 79656
rect 156326 79464 156382 79520
rect 156234 78240 156290 78296
rect 156694 79600 156750 79656
rect 156878 79600 156934 79656
rect 156602 75248 156658 75304
rect 156786 75656 156842 75712
rect 157292 79872 157348 79928
rect 157476 79906 157532 79962
rect 158120 79872 158176 79928
rect 156050 35128 156106 35184
rect 158580 79906 158636 79962
rect 157798 79192 157854 79248
rect 158442 79600 158498 79656
rect 158902 79736 158958 79792
rect 159316 79906 159372 79962
rect 159500 79872 159556 79928
rect 159960 79872 160016 79928
rect 158810 79464 158866 79520
rect 158902 78648 158958 78704
rect 159270 79600 159326 79656
rect 159776 79736 159832 79792
rect 159914 79736 159970 79792
rect 159454 78784 159510 78840
rect 159546 78648 159602 78704
rect 159546 75248 159602 75304
rect 159730 79192 159786 79248
rect 160328 79872 160384 79928
rect 160098 68856 160154 68912
rect 160466 79736 160522 79792
rect 160880 79872 160936 79928
rect 161800 79906 161856 79962
rect 161432 79736 161488 79792
rect 160374 79600 160430 79656
rect 161294 76880 161350 76936
rect 161202 76744 161258 76800
rect 161294 71304 161350 71360
rect 158902 6160 158958 6216
rect 161018 68856 161074 68912
rect 160190 8880 160246 8936
rect 161846 79600 161902 79656
rect 162122 79364 162124 79384
rect 162124 79364 162176 79384
rect 162176 79364 162178 79384
rect 162122 79328 162178 79364
rect 162122 79092 162124 79112
rect 162124 79092 162176 79112
rect 162176 79092 162178 79112
rect 162122 79056 162178 79092
rect 162536 79736 162592 79792
rect 162812 79872 162868 79928
rect 163088 79872 163144 79928
rect 162904 79736 162960 79792
rect 162306 76744 162362 76800
rect 162950 79600 163006 79656
rect 162582 77152 162638 77208
rect 163916 79872 163972 79928
rect 164192 79838 164248 79894
rect 164560 79872 164616 79928
rect 164744 79872 164800 79928
rect 163134 64504 163190 64560
rect 163134 63552 163190 63608
rect 163778 63552 163834 63608
rect 165020 79872 165076 79928
rect 164974 76744 165030 76800
rect 165664 79906 165720 79962
rect 165480 79838 165536 79894
rect 166032 79906 166088 79962
rect 165434 79600 165490 79656
rect 165342 77288 165398 77344
rect 165342 76916 165344 76936
rect 165344 76916 165396 76936
rect 165396 76916 165398 76936
rect 165342 76880 165398 76916
rect 165802 76744 165858 76800
rect 166952 79872 167008 79928
rect 166998 79736 167054 79792
rect 167320 79872 167376 79928
rect 166630 79600 166686 79656
rect 167688 79736 167744 79792
rect 167872 79872 167928 79928
rect 168056 79736 168112 79792
rect 168240 79906 168296 79962
rect 168608 79872 168664 79928
rect 167918 78240 167974 78296
rect 167826 76744 167882 76800
rect 168378 79736 168434 79792
rect 168700 79736 168756 79792
rect 168976 79872 169032 79928
rect 168286 76880 168342 76936
rect 168470 79464 168526 79520
rect 168470 79192 168526 79248
rect 168562 78376 168618 78432
rect 168746 79464 168802 79520
rect 169206 79192 169262 79248
rect 169620 79872 169676 79928
rect 169482 79600 169538 79656
rect 169298 76744 169354 76800
rect 169022 76336 169078 76392
rect 168930 75248 168986 75304
rect 169804 79906 169860 79962
rect 170356 79872 170412 79928
rect 170540 79872 170596 79928
rect 169850 79464 169906 79520
rect 169666 77424 169722 77480
rect 169482 73072 169538 73128
rect 170126 79600 170182 79656
rect 170724 79906 170780 79962
rect 171276 79872 171332 79928
rect 170494 78512 170550 78568
rect 170678 79464 170734 79520
rect 170770 79328 170826 79384
rect 170862 76744 170918 76800
rect 171138 78784 171194 78840
rect 171046 78512 171102 78568
rect 170954 75928 171010 75984
rect 171414 79056 171470 79112
rect 170954 72936 171010 72992
rect 171966 79620 172022 79656
rect 171966 79600 171968 79620
rect 171968 79600 172020 79620
rect 172020 79600 172022 79620
rect 171874 78104 171930 78160
rect 172472 79872 172528 79928
rect 172518 79772 172520 79792
rect 172520 79772 172572 79792
rect 172572 79772 172574 79792
rect 171690 75520 171746 75576
rect 172150 75112 172206 75168
rect 172518 79736 172574 79772
rect 172334 73888 172390 73944
rect 171506 69944 171562 70000
rect 171690 69808 171746 69864
rect 172150 69944 172206 70000
rect 172242 69808 172298 69864
rect 172794 76880 172850 76936
rect 173070 79736 173126 79792
rect 173852 79906 173908 79962
rect 173254 75792 173310 75848
rect 174220 79892 174276 79928
rect 174220 79872 174222 79892
rect 174222 79872 174274 79892
rect 174274 79872 174276 79892
rect 173990 79600 174046 79656
rect 173898 78920 173954 78976
rect 173806 76880 173862 76936
rect 173438 75384 173494 75440
rect 173714 75384 173770 75440
rect 173346 71576 173402 71632
rect 173530 73616 173586 73672
rect 171874 22616 171930 22672
rect 174864 79906 174920 79962
rect 175324 79872 175380 79928
rect 174726 79736 174782 79792
rect 174910 79736 174966 79792
rect 174634 76200 174690 76256
rect 174542 75384 174598 75440
rect 174818 77152 174874 77208
rect 174910 75384 174966 75440
rect 174726 71712 174782 71768
rect 174450 71440 174506 71496
rect 175094 78784 175150 78840
rect 175002 72800 175058 72856
rect 175186 72800 175242 72856
rect 175554 79600 175610 79656
rect 176060 79736 176116 79792
rect 176612 79838 176668 79894
rect 175738 77696 175794 77752
rect 175830 77560 175886 77616
rect 176290 78784 176346 78840
rect 176014 77560 176070 77616
rect 176796 79906 176852 79962
rect 176474 78512 176530 78568
rect 176198 72528 176254 72584
rect 176382 72528 176438 72584
rect 175922 69944 175978 70000
rect 177486 77968 177542 78024
rect 177854 79872 177910 79928
rect 177670 79736 177726 79792
rect 177670 79464 177726 79520
rect 177578 77832 177634 77888
rect 178038 79600 178094 79656
rect 178314 80280 178370 80336
rect 178222 79464 178278 79520
rect 178038 78512 178094 78568
rect 178038 76608 178094 76664
rect 178498 76608 178554 76664
rect 183466 80280 183522 80336
rect 179234 76608 179290 76664
rect 180982 79736 181038 79792
rect 183466 78512 183522 78568
rect 180062 75656 180118 75712
rect 180706 74976 180762 75032
rect 183466 77424 183522 77480
rect 184294 77424 184350 77480
rect 181534 73752 181590 73808
rect 182822 68312 182878 68368
rect 186226 79464 186282 79520
rect 186226 78512 186282 78568
rect 186226 74432 186282 74488
rect 187054 138080 187110 138136
rect 187054 137944 187110 138000
rect 187514 140528 187570 140584
rect 187514 139440 187570 139496
rect 187422 137808 187478 137864
rect 187330 137128 187386 137184
rect 187238 99456 187294 99512
rect 187238 98640 187294 98696
rect 187606 78512 187662 78568
rect 187698 77696 187754 77752
rect 187698 76200 187754 76256
rect 187606 71032 187662 71088
rect 187146 64504 187202 64560
rect 187974 73752 188030 73808
rect 187974 73480 188030 73536
rect 189262 262248 189318 262304
rect 188250 148552 188306 148608
rect 188434 148960 188490 149016
rect 188342 100816 188398 100872
rect 188618 99456 188674 99512
rect 188342 98776 188398 98832
rect 188250 98640 188306 98696
rect 188526 93744 188582 93800
rect 189078 100816 189134 100872
rect 188986 98776 189042 98832
rect 188434 68856 188490 68912
rect 189078 68856 189134 68912
rect 187882 60424 187938 60480
rect 187790 56208 187846 56264
rect 190090 259800 190146 259856
rect 189906 146920 189962 146976
rect 189630 142976 189686 143032
rect 190182 259664 190238 259720
rect 190090 142704 190146 142760
rect 190182 142024 190238 142080
rect 190826 259936 190882 259992
rect 191930 195608 191986 195664
rect 190826 142840 190882 142896
rect 190734 141344 190790 141400
rect 191286 138896 191342 138952
rect 192758 196560 192814 196616
rect 191930 57160 191986 57216
rect 190826 54576 190882 54632
rect 190734 53624 190790 53680
rect 190642 52264 190698 52320
rect 191746 52264 191802 52320
rect 191746 51856 191802 51912
rect 192482 138760 192538 138816
rect 193126 76472 193182 76528
rect 192758 56480 192814 56536
rect 193034 56480 193090 56536
rect 193034 56072 193090 56128
rect 192022 50632 192078 50688
rect 189998 34448 190054 34504
rect 190366 34448 190422 34504
rect 189998 33768 190054 33824
rect 193770 139304 193826 139360
rect 193678 139168 193734 139224
rect 194046 139032 194102 139088
rect 193954 81640 194010 81696
rect 193310 53080 193366 53136
rect 193218 52420 193274 52456
rect 193218 52400 193220 52420
rect 193220 52400 193272 52420
rect 193272 52400 193274 52420
rect 195242 139848 195298 139904
rect 195426 90344 195482 90400
rect 195334 81776 195390 81832
rect 196254 196696 196310 196752
rect 196070 195744 196126 195800
rect 195978 68176 196034 68232
rect 195426 36624 195482 36680
rect 196162 195472 196218 195528
rect 196438 147464 196494 147520
rect 196898 145560 196954 145616
rect 196806 82048 196862 82104
rect 196254 57296 196310 57352
rect 196254 56344 196310 56400
rect 197082 143112 197138 143168
rect 197450 197104 197506 197160
rect 196254 55936 196310 55992
rect 196162 49544 196218 49600
rect 196714 49544 196770 49600
rect 196714 49000 196770 49056
rect 198830 197240 198886 197296
rect 197450 48048 197506 48104
rect 196070 45192 196126 45248
rect 198738 146784 198794 146840
rect 198462 48048 198518 48104
rect 198462 47776 198518 47832
rect 201590 200232 201646 200288
rect 201130 200096 201186 200152
rect 199474 145696 199530 145752
rect 199566 137128 199622 137184
rect 199106 61920 199162 61976
rect 200210 196968 200266 197024
rect 199750 146240 199806 146296
rect 199750 137264 199806 137320
rect 199658 57432 199714 57488
rect 198830 50360 198886 50416
rect 200486 148280 200542 148336
rect 200210 55120 200266 55176
rect 200946 151136 201002 151192
rect 200854 138624 200910 138680
rect 200762 68856 200818 68912
rect 201222 81368 201278 81424
rect 202878 192752 202934 192808
rect 201406 55120 201462 55176
rect 201406 54440 201462 54496
rect 200486 43968 200542 44024
rect 201406 43968 201462 44024
rect 201406 43560 201462 43616
rect 202050 148416 202106 148472
rect 201958 136040 202014 136096
rect 203246 155624 203302 155680
rect 203154 155488 203210 155544
rect 203062 81912 203118 81968
rect 202970 78376 203026 78432
rect 201958 52400 202014 52456
rect 203338 155216 203394 155272
rect 203614 149096 203670 149152
rect 204258 187040 204314 187096
rect 203706 136584 203762 136640
rect 203706 135904 203762 135960
rect 203706 78104 203762 78160
rect 203430 73072 203486 73128
rect 203246 57568 203302 57624
rect 203338 54712 203394 54768
rect 203154 47912 203210 47968
rect 202050 46280 202106 46336
rect 203614 66000 203670 66056
rect 204166 57568 204222 57624
rect 204166 57296 204222 57352
rect 203982 54712 204038 54768
rect 204166 47912 204222 47968
rect 204166 47640 204222 47696
rect 364338 275168 364394 275224
rect 347778 262928 347834 262984
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 579802 590960 579858 591016
rect 580170 577632 580226 577688
rect 579802 564304 579858 564360
rect 580170 537784 580226 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 579986 471416 580042 471472
rect 580170 458088 580226 458144
rect 580170 431568 580226 431624
rect 580170 418240 580226 418296
rect 580170 404912 580226 404968
rect 580170 378392 580226 378448
rect 580262 365064 580318 365120
rect 580170 351908 580172 351928
rect 580172 351908 580224 351928
rect 580224 351908 580226 351928
rect 580170 351872 580226 351908
rect 580170 325216 580226 325272
rect 579986 312024 580042 312080
rect 580170 298696 580226 298752
rect 580170 272176 580226 272232
rect 477498 262792 477554 262848
rect 580170 258848 580226 258904
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 580446 232328 580502 232384
rect 580354 219000 580410 219056
rect 579802 205672 579858 205728
rect 208674 200368 208730 200424
rect 204626 199280 204682 199336
rect 204442 150184 204498 150240
rect 204350 66136 204406 66192
rect 208582 194384 208638 194440
rect 208490 194248 208546 194304
rect 207202 194112 207258 194168
rect 205638 190984 205694 191040
rect 204534 72936 204590 72992
rect 205086 71576 205142 71632
rect 205086 71168 205142 71224
rect 204718 66136 204774 66192
rect 204718 65456 204774 65512
rect 204442 49408 204498 49464
rect 204718 49408 204774 49464
rect 204718 48864 204774 48920
rect 204258 35808 204314 35864
rect 204258 35128 204314 35184
rect 205914 70216 205970 70272
rect 206190 190032 206246 190088
rect 206190 75384 206246 75440
rect 206650 80008 206706 80064
rect 206466 78784 206522 78840
rect 206558 75656 206614 75712
rect 206926 75656 206982 75712
rect 206926 75248 206982 75304
rect 206282 72800 206338 72856
rect 206006 70080 206062 70136
rect 205730 55800 205786 55856
rect 205638 26152 205694 26208
rect 205638 25472 205694 25528
rect 207018 21800 207074 21856
rect 207754 150356 207756 150376
rect 207756 150356 207808 150376
rect 207808 150356 207810 150376
rect 207754 150320 207810 150356
rect 207662 75792 207718 75848
rect 208214 75792 208270 75848
rect 208214 75112 208270 75168
rect 207202 50904 207258 50960
rect 207202 46688 207258 46744
rect 207110 21256 207166 21312
rect 207938 45620 207994 45656
rect 207938 45600 207940 45620
rect 207940 45600 207992 45620
rect 207992 45600 207994 45620
rect 208674 69944 208730 70000
rect 209870 198192 209926 198248
rect 209318 192480 209374 192536
rect 209226 77288 209282 77344
rect 209134 76472 209190 76528
rect 208582 52128 208638 52184
rect 208766 52128 208822 52184
rect 208766 51720 208822 51776
rect 208490 45464 208546 45520
rect 208490 44784 208546 44840
rect 209318 44104 209374 44160
rect 210238 189760 210294 189816
rect 210514 77152 210570 77208
rect 209870 48184 209926 48240
rect 209870 45328 209926 45384
rect 209778 17856 209834 17912
rect 211066 48184 211122 48240
rect 211066 47504 211122 47560
rect 211250 189896 211306 189952
rect 211526 80688 211582 80744
rect 212538 189624 212594 189680
rect 211986 77968 212042 78024
rect 211894 77832 211950 77888
rect 211618 74160 211674 74216
rect 211158 38528 211214 38584
rect 211066 17856 211122 17912
rect 211066 17176 211122 17232
rect 212446 38528 212502 38584
rect 212446 37848 212502 37904
rect 212814 198056 212870 198112
rect 212998 197920 213054 197976
rect 212998 71712 213054 71768
rect 212814 66816 212870 66872
rect 213918 64232 213974 64288
rect 213918 62736 213974 62792
rect 212722 62056 212778 62112
rect 213826 62056 213882 62112
rect 213826 61376 213882 61432
rect 212630 59200 212686 59256
rect 213826 59200 213882 59256
rect 213826 58520 213882 58576
rect 212630 30912 212686 30968
rect 212538 21528 212594 21584
rect 214654 151000 214710 151056
rect 214746 77016 214802 77072
rect 214102 57840 214158 57896
rect 215390 195200 215446 195256
rect 215574 68448 215630 68504
rect 215758 67496 215814 67552
rect 215482 63280 215538 63336
rect 215482 62736 215538 62792
rect 215390 60560 215446 60616
rect 215390 60016 215446 60072
rect 215298 57704 215354 57760
rect 215298 57160 215354 57216
rect 214010 51992 214066 52048
rect 216862 155352 216918 155408
rect 216770 63416 216826 63472
rect 218058 186904 218114 186960
rect 217138 76608 217194 76664
rect 217414 76608 217470 76664
rect 217138 76064 217194 76120
rect 580170 192480 580226 192536
rect 218242 74024 218298 74080
rect 218426 74296 218482 74352
rect 580170 179152 580226 179208
rect 580170 165824 580226 165880
rect 579986 152632 580042 152688
rect 467102 142296 467158 142352
rect 464342 141208 464398 141264
rect 218518 74024 218574 74080
rect 218426 73888 218482 73944
rect 218242 73344 218298 73400
rect 220818 68448 220874 68504
rect 218058 46824 218114 46880
rect 216862 37168 216918 37224
rect 217230 37168 217286 37224
rect 217230 36488 217286 36544
rect 227718 67496 227774 67552
rect 231858 60152 231914 60208
rect 237378 74024 237434 74080
rect 234710 33768 234766 33824
rect 251178 46416 251234 46472
rect 260102 76608 260158 76664
rect 259458 51992 259514 52048
rect 269118 73752 269174 73808
rect 263598 57568 263654 57624
rect 284298 73888 284354 73944
rect 276110 43832 276166 43888
rect 284390 56208 284446 56264
rect 302238 78648 302294 78704
rect 293958 37848 294014 37904
rect 300858 17176 300914 17232
rect 306378 64232 306434 64288
rect 307022 36624 307078 36680
rect 311162 35128 311218 35184
rect 320178 51856 320234 51912
rect 574742 141072 574798 141128
rect 523130 80688 523186 80744
rect 331218 56072 331274 56128
rect 333978 53216 334034 53272
rect 338118 50632 338174 50688
rect 336738 21528 336794 21584
rect 350538 21392 350594 21448
rect 354678 21256 354734 21312
rect 364982 53080 365038 53136
rect 372618 62872 372674 62928
rect 369858 54576 369914 54632
rect 373998 50496 374054 50552
rect 389178 76472 389234 76528
rect 382922 55936 382978 55992
rect 387798 49000 387854 49056
rect 390558 45192 390614 45248
rect 394698 60016 394754 60072
rect 405738 47776 405794 47832
rect 408498 43696 408554 43752
rect 414662 57432 414718 57488
rect 418802 50360 418858 50416
rect 418158 25472 418214 25528
rect 423770 59880 423826 59936
rect 427818 43560 427874 43616
rect 440238 54440 440294 54496
rect 444378 45056 444434 45112
rect 465170 78376 465226 78432
rect 456798 78240 456854 78296
rect 454038 46280 454094 46336
rect 455418 46144 455474 46200
rect 460938 72392 460994 72448
rect 458178 43424 458234 43480
rect 471978 78104 472034 78160
rect 466458 47640 466514 47696
rect 478142 71440 478198 71496
rect 473450 57296 473506 57352
rect 482282 75384 482338 75440
rect 498842 71304 498898 71360
rect 494058 66816 494114 66872
rect 486422 65456 486478 65512
rect 490010 47504 490066 47560
rect 499578 55800 499634 55856
rect 509882 75248 509938 75304
rect 514022 58520 514078 58576
rect 520922 44920 520978 44976
rect 524418 75112 524474 75168
rect 531318 71168 531374 71224
rect 526442 61376 526498 61432
rect 548522 71032 548578 71088
rect 535458 44784 535514 44840
rect 543738 64096 543794 64152
rect 540242 62736 540298 62792
rect 542358 51720 542414 51776
rect 552018 36488 552074 36544
rect 557538 69536 557594 69592
rect 556158 50224 556214 50280
rect 567842 57160 567898 57216
rect 565818 48864 565874 48920
rect 580170 99456 580226 99512
rect 579986 86128 580042 86184
rect 579618 72936 579674 72992
rect 580170 19760 580226 19816
rect 580354 142160 580410 142216
rect 580814 140936 580870 140992
rect 580630 140800 580686 140856
rect 580814 125976 580870 126032
rect 580630 112784 580686 112840
rect 580998 77968 581054 78024
rect 580538 59608 580594 59664
rect 580446 46280 580502 46336
rect 580354 33088 580410 33144
rect 580262 6568 580318 6624
rect 581090 77832 581146 77888
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3141 619170 3207 619173
rect -960 619168 3207 619170
rect -960 619112 3146 619168
rect 3202 619112 3207 619168
rect -960 619110 3207 619112
rect -960 619020 480 619110
rect 3141 619107 3207 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3233 606114 3299 606117
rect -960 606112 3299 606114
rect -960 606056 3238 606112
rect 3294 606056 3299 606112
rect -960 606054 3299 606056
rect -960 605964 480 606054
rect 3233 606051 3299 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 579797 564362 579863 564365
rect 583520 564362 584960 564452
rect 579797 564360 584960 564362
rect 579797 564304 579802 564360
rect 579858 564304 584960 564360
rect 579797 564302 584960 564304
rect 579797 564299 579863 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3417 553890 3483 553893
rect -960 553888 3483 553890
rect -960 553832 3422 553888
rect 3478 553832 3483 553888
rect -960 553830 3483 553832
rect -960 553740 480 553830
rect 3417 553827 3483 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3417 527914 3483 527917
rect -960 527912 3483 527914
rect -960 527856 3422 527912
rect 3478 527856 3483 527912
rect -960 527854 3483 527856
rect -960 527764 480 527854
rect 3417 527851 3483 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3417 514858 3483 514861
rect -960 514856 3483 514858
rect -960 514800 3422 514856
rect 3478 514800 3483 514856
rect -960 514798 3483 514800
rect -960 514708 480 514798
rect 3417 514795 3483 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3049 501802 3115 501805
rect -960 501800 3115 501802
rect -960 501744 3054 501800
rect 3110 501744 3115 501800
rect -960 501742 3115 501744
rect -960 501652 480 501742
rect 3049 501739 3115 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3417 475690 3483 475693
rect -960 475688 3483 475690
rect -960 475632 3422 475688
rect 3478 475632 3483 475688
rect -960 475630 3483 475632
rect -960 475540 480 475630
rect 3417 475627 3483 475630
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3509 462634 3575 462637
rect -960 462632 3575 462634
rect -960 462576 3514 462632
rect 3570 462576 3575 462632
rect -960 462574 3575 462576
rect -960 462484 480 462574
rect 3509 462571 3575 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3509 423602 3575 423605
rect -960 423600 3575 423602
rect -960 423544 3514 423600
rect 3570 423544 3575 423600
rect -960 423542 3575 423544
rect -960 423452 480 423542
rect 3509 423539 3575 423542
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 2865 410546 2931 410549
rect -960 410544 2931 410546
rect -960 410488 2870 410544
rect 2926 410488 2931 410544
rect -960 410486 2931 410488
rect -960 410396 480 410486
rect 2865 410483 2931 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3509 397490 3575 397493
rect -960 397488 3575 397490
rect -960 397432 3514 397488
rect 3570 397432 3575 397488
rect -960 397430 3575 397432
rect -960 397340 480 397430
rect 3509 397427 3575 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 2773 371378 2839 371381
rect -960 371376 2839 371378
rect -960 371320 2778 371376
rect 2834 371320 2839 371376
rect -960 371318 2839 371320
rect -960 371228 480 371318
rect 2773 371315 2839 371318
rect 580257 365122 580323 365125
rect 583520 365122 584960 365212
rect 580257 365120 584960 365122
rect 580257 365064 580262 365120
rect 580318 365064 584960 365120
rect 580257 365062 584960 365064
rect 580257 365059 580323 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3141 358458 3207 358461
rect -960 358456 3207 358458
rect -960 358400 3146 358456
rect 3202 358400 3207 358456
rect -960 358398 3207 358400
rect -960 358308 480 358398
rect 3141 358395 3207 358398
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3509 345402 3575 345405
rect -960 345400 3575 345402
rect -960 345344 3514 345400
rect 3570 345344 3575 345400
rect -960 345342 3575 345344
rect -960 345252 480 345342
rect 3509 345339 3575 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3325 319290 3391 319293
rect -960 319288 3391 319290
rect -960 319232 3330 319288
rect 3386 319232 3391 319288
rect -960 319230 3391 319232
rect -960 319140 480 319230
rect 3325 319227 3391 319230
rect 579981 312082 580047 312085
rect 583520 312082 584960 312172
rect 579981 312080 584960 312082
rect 579981 312024 579986 312080
rect 580042 312024 584960 312080
rect 579981 312022 584960 312024
rect 579981 312019 580047 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3509 306234 3575 306237
rect -960 306232 3575 306234
rect -960 306176 3514 306232
rect 3570 306176 3575 306232
rect -960 306174 3575 306176
rect -960 306084 480 306174
rect 3509 306171 3575 306174
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3509 293178 3575 293181
rect -960 293176 3575 293178
rect -960 293120 3514 293176
rect 3570 293120 3575 293176
rect -960 293118 3575 293120
rect -960 293028 480 293118
rect 3509 293115 3575 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 364333 275226 364399 275229
rect 190410 275224 364399 275226
rect 190410 275168 364338 275224
rect 364394 275168 364399 275224
rect 190410 275166 364399 275168
rect 151813 274682 151879 274685
rect 187734 274682 187740 274684
rect 151813 274680 187740 274682
rect 151813 274624 151818 274680
rect 151874 274624 187740 274680
rect 151813 274622 187740 274624
rect 151813 274619 151879 274622
rect 187734 274620 187740 274622
rect 187804 274682 187810 274684
rect 190410 274682 190470 275166
rect 364333 275163 364399 275166
rect 187804 274622 190470 274682
rect 187804 274620 187810 274622
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3049 267202 3115 267205
rect -960 267200 3115 267202
rect -960 267144 3054 267200
rect 3110 267144 3115 267200
rect -960 267142 3115 267144
rect -960 267052 480 267142
rect 3049 267139 3115 267142
rect 109534 265236 109540 265300
rect 109604 265298 109610 265300
rect 135897 265298 135963 265301
rect 109604 265296 135963 265298
rect 109604 265240 135902 265296
rect 135958 265240 135963 265296
rect 109604 265238 135963 265240
rect 109604 265236 109610 265238
rect 135897 265235 135963 265238
rect 169017 265298 169083 265301
rect 197670 265298 197676 265300
rect 169017 265296 197676 265298
rect 169017 265240 169022 265296
rect 169078 265240 197676 265296
rect 169017 265238 197676 265240
rect 169017 265235 169083 265238
rect 197670 265236 197676 265238
rect 197740 265236 197746 265300
rect 115790 265100 115796 265164
rect 115860 265162 115866 265164
rect 148501 265162 148567 265165
rect 115860 265160 148567 265162
rect 115860 265104 148506 265160
rect 148562 265104 148567 265160
rect 115860 265102 148567 265104
rect 115860 265100 115866 265102
rect 148501 265099 148567 265102
rect 167545 265162 167611 265165
rect 198958 265162 198964 265164
rect 167545 265160 198964 265162
rect 167545 265104 167550 265160
rect 167606 265104 198964 265160
rect 167545 265102 198964 265104
rect 167545 265099 167611 265102
rect 198958 265100 198964 265102
rect 199028 265100 199034 265164
rect 112846 264964 112852 265028
rect 112916 265026 112922 265028
rect 147029 265026 147095 265029
rect 112916 265024 147095 265026
rect 112916 264968 147034 265024
rect 147090 264968 147095 265024
rect 112916 264966 147095 264968
rect 112916 264964 112922 264966
rect 147029 264963 147095 264966
rect 163497 265026 163563 265029
rect 197486 265026 197492 265028
rect 163497 265024 197492 265026
rect 163497 264968 163502 265024
rect 163558 264968 197492 265024
rect 163497 264966 197492 264968
rect 163497 264963 163563 264966
rect 197486 264964 197492 264966
rect 197556 264964 197562 265028
rect 121126 263876 121132 263940
rect 121196 263938 121202 263940
rect 142613 263938 142679 263941
rect 121196 263936 142679 263938
rect 121196 263880 142618 263936
rect 142674 263880 142679 263936
rect 121196 263878 142679 263880
rect 121196 263876 121202 263878
rect 142613 263875 142679 263878
rect 121310 263740 121316 263804
rect 121380 263802 121386 263804
rect 146201 263802 146267 263805
rect 121380 263800 146267 263802
rect 121380 263744 146206 263800
rect 146262 263744 146267 263800
rect 121380 263742 146267 263744
rect 121380 263740 121386 263742
rect 146201 263739 146267 263742
rect 118366 263604 118372 263668
rect 118436 263666 118442 263668
rect 151077 263666 151143 263669
rect 118436 263664 151143 263666
rect 118436 263608 151082 263664
rect 151138 263608 151143 263664
rect 118436 263606 151143 263608
rect 118436 263604 118442 263606
rect 151077 263603 151143 263606
rect 145005 263122 145071 263125
rect 145649 263122 145715 263125
rect 145005 263120 145715 263122
rect 145005 263064 145010 263120
rect 145066 263064 145654 263120
rect 145710 263064 145715 263120
rect 145005 263062 145715 263064
rect 145005 263059 145071 263062
rect 145649 263059 145715 263062
rect 187693 262986 187759 262989
rect 347773 262986 347839 262989
rect 187693 262984 347839 262986
rect 187693 262928 187698 262984
rect 187754 262928 347778 262984
rect 347834 262928 347839 262984
rect 187693 262926 347839 262928
rect 187693 262923 187759 262926
rect 347773 262923 347839 262926
rect 114134 262788 114140 262852
rect 114204 262850 114210 262852
rect 138657 262850 138723 262853
rect 477493 262850 477559 262853
rect 114204 262848 138723 262850
rect 114204 262792 138662 262848
rect 138718 262792 138723 262848
rect 114204 262790 138723 262792
rect 114204 262788 114210 262790
rect 138657 262787 138723 262790
rect 151770 262848 477559 262850
rect 151770 262792 477498 262848
rect 477554 262792 477559 262848
rect 151770 262790 477559 262792
rect 120809 262714 120875 262717
rect 150525 262714 150591 262717
rect 151770 262714 151830 262790
rect 477493 262787 477559 262790
rect 120809 262712 151830 262714
rect 120809 262656 120814 262712
rect 120870 262656 150530 262712
rect 150586 262656 151830 262712
rect 120809 262654 151830 262656
rect 158805 262714 158871 262717
rect 159909 262714 159975 262717
rect 193622 262714 193628 262716
rect 158805 262712 193628 262714
rect 158805 262656 158810 262712
rect 158866 262656 159914 262712
rect 159970 262656 193628 262712
rect 158805 262654 193628 262656
rect 120809 262651 120875 262654
rect 150525 262651 150591 262654
rect 158805 262651 158871 262654
rect 159909 262651 159975 262654
rect 193622 262652 193628 262654
rect 193692 262652 193698 262716
rect 111558 262516 111564 262580
rect 111628 262578 111634 262580
rect 142245 262578 142311 262581
rect 142889 262578 142955 262581
rect 111628 262576 142955 262578
rect 111628 262520 142250 262576
rect 142306 262520 142894 262576
rect 142950 262520 142955 262576
rect 111628 262518 142955 262520
rect 111628 262516 111634 262518
rect 142245 262515 142311 262518
rect 142889 262515 142955 262518
rect 162025 262578 162091 262581
rect 193438 262578 193444 262580
rect 162025 262576 193444 262578
rect 162025 262520 162030 262576
rect 162086 262520 193444 262576
rect 162025 262518 193444 262520
rect 162025 262515 162091 262518
rect 193438 262516 193444 262518
rect 193508 262516 193514 262580
rect 115105 262442 115171 262445
rect 146937 262442 147003 262445
rect 115105 262440 147003 262442
rect 115105 262384 115110 262440
rect 115166 262384 146942 262440
rect 146998 262384 147003 262440
rect 115105 262382 147003 262384
rect 115105 262379 115171 262382
rect 146937 262379 147003 262382
rect 153653 262442 153719 262445
rect 187693 262442 187759 262445
rect 187969 262442 188035 262445
rect 153653 262440 188035 262442
rect 153653 262384 153658 262440
rect 153714 262384 187698 262440
rect 187754 262384 187974 262440
rect 188030 262384 188035 262440
rect 153653 262382 188035 262384
rect 153653 262379 153719 262382
rect 187693 262379 187759 262382
rect 187969 262379 188035 262382
rect 112529 262306 112595 262309
rect 145005 262306 145071 262309
rect 189257 262308 189323 262309
rect 189206 262306 189212 262308
rect 112529 262304 145071 262306
rect 112529 262248 112534 262304
rect 112590 262248 145010 262304
rect 145066 262248 145071 262304
rect 112529 262246 145071 262248
rect 189166 262246 189212 262306
rect 189276 262304 189323 262308
rect 189318 262248 189323 262304
rect 112529 262243 112595 262246
rect 145005 262243 145071 262246
rect 189206 262244 189212 262246
rect 189276 262244 189323 262248
rect 189257 262243 189323 262244
rect 111374 261156 111380 261220
rect 111444 261218 111450 261220
rect 125593 261218 125659 261221
rect 111444 261216 125659 261218
rect 111444 261160 125598 261216
rect 125654 261160 125659 261216
rect 111444 261158 125659 261160
rect 111444 261156 111450 261158
rect 125593 261155 125659 261158
rect 109350 261020 109356 261084
rect 109420 261082 109426 261084
rect 133965 261082 134031 261085
rect 109420 261080 134031 261082
rect 109420 261024 133970 261080
rect 134026 261024 134031 261080
rect 109420 261022 134031 261024
rect 109420 261020 109426 261022
rect 133965 261019 134031 261022
rect 111190 260884 111196 260948
rect 111260 260946 111266 260948
rect 137461 260946 137527 260949
rect 111260 260944 137527 260946
rect 111260 260888 137466 260944
rect 137522 260888 137527 260944
rect 111260 260886 137527 260888
rect 111260 260884 111266 260886
rect 137461 260883 137527 260886
rect 161473 260810 161539 260813
rect 162669 260810 162735 260813
rect 161473 260808 162735 260810
rect 161473 260752 161478 260808
rect 161534 260752 162674 260808
rect 162730 260752 162735 260808
rect 161473 260750 162735 260752
rect 161473 260747 161539 260750
rect 162669 260747 162735 260750
rect 147673 260266 147739 260269
rect 148363 260266 148429 260269
rect 147673 260264 148429 260266
rect 147673 260208 147678 260264
rect 147734 260208 148368 260264
rect 148424 260208 148429 260264
rect 147673 260206 148429 260208
rect 147673 260203 147739 260206
rect 148363 260203 148429 260206
rect 140773 260130 140839 260133
rect 140773 260128 140882 260130
rect 140773 260072 140778 260128
rect 140834 260072 140882 260128
rect 140773 260067 140882 260072
rect 116894 259932 116900 259996
rect 116964 259994 116970 259996
rect 140822 259994 140882 260067
rect 141417 259994 141483 259997
rect 116964 259992 141483 259994
rect 116964 259936 141422 259992
rect 141478 259936 141483 259992
rect 116964 259934 141483 259936
rect 116964 259932 116970 259934
rect 141417 259931 141483 259934
rect 160093 259994 160159 259997
rect 160921 259994 160987 259997
rect 190821 259994 190887 259997
rect 160093 259992 160987 259994
rect 160093 259936 160098 259992
rect 160154 259936 160926 259992
rect 160982 259936 160987 259992
rect 160093 259934 160987 259936
rect 160093 259931 160159 259934
rect 160921 259931 160987 259934
rect 180750 259992 190887 259994
rect 180750 259936 190826 259992
rect 190882 259936 190887 259992
rect 180750 259934 190887 259936
rect 119429 259858 119495 259861
rect 147673 259858 147739 259861
rect 119429 259856 147739 259858
rect 119429 259800 119434 259856
rect 119490 259800 147678 259856
rect 147734 259800 147739 259856
rect 119429 259798 147739 259800
rect 119429 259795 119495 259798
rect 147673 259795 147739 259798
rect 162577 259858 162643 259861
rect 180750 259858 180810 259934
rect 190821 259931 190887 259934
rect 190085 259858 190151 259861
rect 162577 259856 180810 259858
rect 162577 259800 162582 259856
rect 162638 259800 180810 259856
rect 162577 259798 180810 259800
rect 185350 259856 190151 259858
rect 185350 259800 190090 259856
rect 190146 259800 190151 259856
rect 185350 259798 190151 259800
rect 162577 259795 162643 259798
rect 115289 259722 115355 259725
rect 148133 259722 148199 259725
rect 115289 259720 148199 259722
rect 115289 259664 115294 259720
rect 115350 259664 148138 259720
rect 148194 259664 148199 259720
rect 115289 259662 148199 259664
rect 115289 259659 115355 259662
rect 148133 259659 148199 259662
rect 161197 259722 161263 259725
rect 185350 259722 185410 259798
rect 190085 259795 190151 259798
rect 190177 259722 190243 259725
rect 161197 259720 185410 259722
rect 161197 259664 161202 259720
rect 161258 259664 185410 259720
rect 161197 259662 185410 259664
rect 185534 259720 190243 259722
rect 185534 259664 190182 259720
rect 190238 259664 190243 259720
rect 185534 259662 190243 259664
rect 161197 259659 161263 259662
rect 116710 259524 116716 259588
rect 116780 259586 116786 259588
rect 149237 259586 149303 259589
rect 116780 259584 149303 259586
rect 116780 259528 149242 259584
rect 149298 259528 149303 259584
rect 116780 259526 149303 259528
rect 116780 259524 116786 259526
rect 149237 259523 149303 259526
rect 155217 259586 155283 259589
rect 185534 259586 185594 259662
rect 190177 259659 190243 259662
rect 155217 259584 185594 259586
rect 155217 259528 155222 259584
rect 155278 259528 185594 259584
rect 155217 259526 185594 259528
rect 185669 259586 185735 259589
rect 186078 259586 186084 259588
rect 185669 259584 186084 259586
rect 185669 259528 185674 259584
rect 185730 259528 186084 259584
rect 185669 259526 186084 259528
rect 155217 259523 155283 259526
rect 185669 259523 185735 259526
rect 186078 259524 186084 259526
rect 186148 259524 186154 259588
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3509 254146 3575 254149
rect -960 254144 3575 254146
rect -960 254088 3514 254144
rect 3570 254088 3575 254144
rect -960 254086 3575 254088
rect -960 253996 480 254086
rect 3509 254083 3575 254086
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 2773 241090 2839 241093
rect -960 241088 2839 241090
rect -960 241032 2778 241088
rect 2834 241032 2839 241088
rect -960 241030 2839 241032
rect -960 240940 480 241030
rect 2773 241027 2839 241030
rect 580441 232386 580507 232389
rect 583520 232386 584960 232476
rect 580441 232384 584960 232386
rect 580441 232328 580446 232384
rect 580502 232328 584960 232384
rect 580441 232326 584960 232328
rect 580441 232323 580507 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 580349 219058 580415 219061
rect 583520 219058 584960 219148
rect 580349 219056 584960 219058
rect 580349 219000 580354 219056
rect 580410 219000 584960 219056
rect 580349 218998 584960 219000
rect 580349 218995 580415 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3509 214978 3575 214981
rect -960 214976 3575 214978
rect -960 214920 3514 214976
rect 3570 214920 3575 214976
rect -960 214918 3575 214920
rect -960 214828 480 214918
rect 3509 214915 3575 214918
rect 186078 212468 186084 212532
rect 186148 212530 186154 212532
rect 187182 212530 187188 212532
rect 186148 212470 187188 212530
rect 186148 212468 186154 212470
rect 187182 212468 187188 212470
rect 187252 212468 187258 212532
rect 579797 205730 579863 205733
rect 583520 205730 584960 205820
rect 579797 205728 584960 205730
rect 579797 205672 579802 205728
rect 579858 205672 584960 205728
rect 579797 205670 584960 205672
rect 579797 205667 579863 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3417 201922 3483 201925
rect -960 201920 3483 201922
rect -960 201864 3422 201920
rect 3478 201864 3483 201920
rect -960 201862 3483 201864
rect -960 201772 480 201862
rect 3417 201859 3483 201862
rect 132166 201180 132172 201244
rect 132236 201242 132242 201244
rect 139894 201242 139900 201244
rect 132236 201182 139900 201242
rect 132236 201180 132242 201182
rect 139894 201180 139900 201182
rect 139964 201180 139970 201244
rect 131614 201044 131620 201108
rect 131684 201106 131690 201108
rect 138790 201106 138796 201108
rect 131684 201046 138796 201106
rect 131684 201044 131690 201046
rect 138790 201044 138796 201046
rect 138860 201044 138866 201108
rect 151486 200970 151492 200972
rect 131070 200910 151492 200970
rect 117078 200772 117084 200836
rect 117148 200834 117154 200836
rect 131070 200834 131130 200910
rect 151486 200908 151492 200910
rect 151556 200908 151562 200972
rect 117148 200774 131130 200834
rect 117148 200772 117154 200774
rect 131798 200772 131804 200836
rect 131868 200834 131874 200836
rect 136582 200834 136588 200836
rect 131868 200774 136588 200834
rect 131868 200772 131874 200774
rect 136582 200772 136588 200774
rect 136652 200772 136658 200836
rect 127709 200698 127775 200701
rect 153326 200698 153332 200700
rect 127709 200696 153332 200698
rect 127709 200640 127714 200696
rect 127770 200640 153332 200696
rect 127709 200638 153332 200640
rect 127709 200635 127775 200638
rect 153326 200636 153332 200638
rect 153396 200636 153402 200700
rect 106774 200500 106780 200564
rect 106844 200562 106850 200564
rect 131481 200562 131547 200565
rect 106844 200560 131547 200562
rect 106844 200504 131486 200560
rect 131542 200504 131547 200560
rect 106844 200502 131547 200504
rect 106844 200500 106850 200502
rect 131481 200499 131547 200502
rect 132125 200562 132191 200565
rect 140078 200562 140084 200564
rect 132125 200560 140084 200562
rect 132125 200504 132130 200560
rect 132186 200504 140084 200560
rect 132125 200502 140084 200504
rect 132125 200499 132191 200502
rect 140078 200500 140084 200502
rect 140148 200500 140154 200564
rect 180149 200562 180215 200565
rect 207054 200562 207060 200564
rect 180149 200560 207060 200562
rect 180149 200504 180154 200560
rect 180210 200504 207060 200560
rect 180149 200502 207060 200504
rect 180149 200499 180215 200502
rect 207054 200500 207060 200502
rect 207124 200500 207130 200564
rect 122414 200364 122420 200428
rect 122484 200426 122490 200428
rect 151670 200426 151676 200428
rect 122484 200366 151676 200426
rect 122484 200364 122490 200366
rect 151670 200364 151676 200366
rect 151740 200364 151746 200428
rect 180333 200426 180399 200429
rect 208669 200426 208735 200429
rect 152782 200366 156522 200426
rect 122598 200228 122604 200292
rect 122668 200290 122674 200292
rect 152782 200290 152842 200366
rect 122668 200230 152842 200290
rect 122668 200228 122674 200230
rect 131573 200154 131639 200157
rect 131573 200152 138582 200154
rect 131573 200096 131578 200152
rect 131634 200096 138582 200152
rect 131573 200094 138582 200096
rect 131573 200091 131639 200094
rect 130101 200018 130167 200021
rect 133454 200018 133460 200020
rect 130101 200016 133460 200018
rect 130101 199960 130106 200016
rect 130162 199960 133460 200016
rect 130101 199958 133460 199960
rect 130101 199955 130167 199958
rect 133454 199956 133460 199958
rect 133524 199956 133530 200020
rect 138522 199919 138582 200094
rect 140078 200092 140084 200156
rect 140148 200154 140154 200156
rect 154798 200154 154804 200156
rect 140148 200094 151048 200154
rect 140148 200092 140154 200094
rect 133643 199914 133709 199919
rect 131941 199882 132007 199885
rect 132999 199882 133065 199885
rect 133643 199884 133648 199914
rect 133704 199884 133709 199914
rect 136403 199914 136469 199919
rect 136863 199916 136929 199919
rect 131941 199880 133065 199882
rect 131941 199824 131946 199880
rect 132002 199824 133004 199880
rect 133060 199824 133065 199880
rect 131941 199822 133065 199824
rect 131941 199819 132007 199822
rect 132999 199819 133065 199822
rect 133638 199820 133644 199884
rect 133708 199882 133714 199884
rect 133708 199822 133766 199882
rect 133708 199820 133714 199822
rect 134190 199820 134196 199884
rect 134260 199882 134266 199884
rect 134747 199882 134813 199885
rect 134260 199880 134813 199882
rect 134260 199824 134752 199880
rect 134808 199824 134813 199880
rect 134260 199822 134813 199824
rect 134260 199820 134266 199822
rect 134747 199819 134813 199822
rect 135294 199820 135300 199884
rect 135364 199882 135370 199884
rect 135575 199882 135641 199885
rect 136403 199884 136408 199914
rect 136464 199884 136469 199914
rect 136590 199914 136929 199916
rect 135364 199880 135641 199882
rect 135364 199824 135580 199880
rect 135636 199824 135641 199880
rect 135364 199822 135641 199824
rect 135364 199820 135370 199822
rect 135575 199819 135641 199822
rect 136398 199820 136404 199884
rect 136468 199882 136474 199884
rect 136468 199822 136526 199882
rect 136590 199858 136868 199914
rect 136924 199858 136929 199914
rect 137139 199914 137205 199919
rect 137139 199884 137144 199914
rect 137200 199884 137205 199914
rect 137507 199914 137573 199919
rect 137507 199884 137512 199914
rect 137568 199884 137573 199914
rect 138335 199914 138401 199919
rect 136590 199856 136929 199858
rect 136468 199820 136474 199822
rect 132953 199746 133019 199749
rect 136590 199746 136650 199856
rect 136863 199853 136929 199856
rect 137134 199820 137140 199884
rect 137204 199882 137210 199884
rect 137204 199822 137262 199882
rect 137204 199820 137210 199822
rect 137502 199820 137508 199884
rect 137572 199882 137578 199884
rect 137572 199822 137630 199882
rect 137572 199820 137578 199822
rect 138054 199820 138060 199884
rect 138124 199882 138130 199884
rect 138335 199882 138340 199914
rect 138124 199858 138340 199882
rect 138396 199858 138401 199914
rect 138124 199853 138401 199858
rect 138519 199914 138585 199919
rect 138519 199858 138524 199914
rect 138580 199858 138585 199914
rect 138795 199914 138861 199919
rect 138795 199884 138800 199914
rect 138856 199884 138861 199914
rect 139255 199916 139321 199919
rect 139255 199914 139456 199916
rect 138519 199853 138585 199858
rect 138124 199822 138398 199853
rect 138124 199820 138130 199822
rect 138790 199820 138796 199884
rect 138860 199882 138866 199884
rect 138860 199822 138918 199882
rect 139255 199858 139260 199914
rect 139316 199858 139456 199914
rect 139531 199914 139597 199919
rect 139531 199884 139536 199914
rect 139592 199884 139597 199914
rect 139899 199914 139965 199919
rect 139899 199884 139904 199914
rect 139960 199884 139965 199914
rect 140083 199914 140149 199919
rect 139255 199856 139456 199858
rect 139255 199853 139321 199856
rect 138860 199820 138866 199822
rect 139396 199749 139456 199856
rect 139526 199820 139532 199884
rect 139596 199882 139602 199884
rect 139596 199822 139654 199882
rect 139596 199820 139602 199822
rect 139894 199820 139900 199884
rect 139964 199882 139970 199884
rect 139964 199822 140022 199882
rect 140083 199858 140088 199914
rect 140144 199858 140149 199914
rect 140911 199916 140977 199919
rect 140911 199914 141020 199916
rect 140083 199853 140149 199858
rect 140635 199880 140701 199885
rect 139964 199820 139970 199822
rect 140086 199749 140146 199853
rect 140635 199824 140640 199880
rect 140696 199824 140701 199880
rect 140911 199858 140916 199914
rect 140972 199884 141020 199914
rect 141187 199914 141253 199919
rect 140972 199858 141004 199884
rect 140911 199853 141004 199858
rect 140635 199819 140701 199824
rect 140960 199822 141004 199853
rect 140998 199820 141004 199822
rect 141068 199820 141074 199884
rect 141187 199858 141192 199914
rect 141248 199858 141253 199914
rect 141187 199853 141253 199858
rect 141555 199916 141621 199919
rect 141555 199914 141986 199916
rect 141555 199858 141560 199914
rect 141616 199882 141986 199914
rect 142659 199914 142725 199919
rect 143119 199916 143185 199919
rect 142286 199882 142292 199884
rect 141616 199858 142292 199882
rect 141555 199856 142292 199858
rect 141555 199853 141621 199856
rect 132953 199744 136650 199746
rect 132953 199688 132958 199744
rect 133014 199688 136650 199744
rect 132953 199686 136650 199688
rect 139393 199744 139459 199749
rect 139393 199688 139398 199744
rect 139454 199688 139459 199744
rect 132953 199683 133019 199686
rect 139393 199683 139459 199688
rect 140037 199744 140146 199749
rect 140037 199688 140042 199744
rect 140098 199688 140146 199744
rect 140037 199686 140146 199688
rect 140497 199746 140563 199749
rect 140638 199746 140698 199819
rect 140497 199744 140698 199746
rect 140497 199688 140502 199744
rect 140558 199688 140698 199744
rect 140497 199686 140698 199688
rect 140957 199746 141023 199749
rect 141190 199746 141250 199853
rect 141926 199822 142292 199856
rect 142286 199820 142292 199822
rect 142356 199820 142362 199884
rect 142659 199882 142664 199914
rect 142478 199858 142664 199882
rect 142720 199858 142725 199914
rect 143076 199914 143185 199916
rect 143076 199884 143124 199914
rect 142478 199853 142725 199858
rect 142478 199822 142722 199853
rect 140957 199744 141250 199746
rect 140957 199688 140962 199744
rect 141018 199688 141250 199744
rect 140957 199686 141250 199688
rect 140037 199683 140103 199686
rect 140497 199683 140563 199686
rect 140957 199683 141023 199686
rect 141550 199684 141556 199748
rect 141620 199746 141626 199748
rect 142478 199746 142538 199822
rect 143022 199820 143028 199884
rect 143092 199858 143124 199884
rect 143180 199858 143185 199914
rect 143092 199853 143185 199858
rect 143395 199914 143461 199919
rect 143395 199858 143400 199914
rect 143456 199858 143461 199914
rect 143395 199853 143461 199858
rect 144039 199916 144105 199919
rect 144223 199916 144289 199919
rect 144039 199914 144148 199916
rect 144039 199858 144044 199914
rect 144100 199858 144148 199914
rect 144039 199853 144148 199858
rect 144223 199914 144424 199916
rect 144223 199858 144228 199914
rect 144284 199858 144424 199914
rect 144223 199856 144424 199858
rect 144223 199853 144289 199856
rect 143092 199822 143136 199853
rect 143092 199820 143098 199822
rect 143027 199746 143093 199749
rect 141620 199686 142538 199746
rect 142662 199744 143093 199746
rect 142662 199688 143032 199744
rect 143088 199688 143093 199744
rect 142662 199686 143093 199688
rect 141620 199684 141626 199686
rect 131757 199612 131823 199613
rect 131757 199610 131804 199612
rect 131712 199608 131804 199610
rect 131712 199552 131762 199608
rect 131712 199550 131804 199552
rect 131757 199548 131804 199550
rect 131868 199548 131874 199612
rect 132217 199610 132283 199613
rect 141182 199610 141188 199612
rect 132217 199608 141188 199610
rect 132217 199552 132222 199608
rect 132278 199552 141188 199608
rect 132217 199550 141188 199552
rect 131757 199547 131823 199548
rect 132217 199547 132283 199550
rect 141182 199548 141188 199550
rect 141252 199548 141258 199612
rect 141785 199610 141851 199613
rect 141918 199610 141924 199612
rect 141785 199608 141924 199610
rect 141785 199552 141790 199608
rect 141846 199552 141924 199608
rect 141785 199550 141924 199552
rect 141785 199547 141851 199550
rect 141918 199548 141924 199550
rect 141988 199548 141994 199612
rect 142662 199477 142722 199686
rect 143027 199683 143093 199686
rect 143398 199613 143458 199853
rect 144088 199746 144148 199853
rect 142838 199548 142844 199612
rect 142908 199610 142914 199612
rect 142908 199550 143274 199610
rect 142908 199548 142914 199550
rect 131573 199476 131639 199477
rect 132125 199476 132191 199477
rect 131573 199474 131620 199476
rect 131528 199472 131620 199474
rect 131528 199416 131578 199472
rect 131528 199414 131620 199416
rect 131573 199412 131620 199414
rect 131684 199412 131690 199476
rect 132125 199474 132172 199476
rect 132080 199472 132172 199474
rect 132080 199416 132130 199472
rect 132080 199414 132172 199416
rect 132125 199412 132172 199414
rect 132236 199412 132242 199476
rect 132309 199474 132375 199477
rect 134609 199474 134675 199477
rect 132309 199472 134675 199474
rect 132309 199416 132314 199472
rect 132370 199416 134614 199472
rect 134670 199416 134675 199472
rect 132309 199414 134675 199416
rect 131573 199411 131639 199412
rect 132125 199411 132191 199412
rect 132309 199411 132375 199414
rect 134609 199411 134675 199414
rect 135253 199474 135319 199477
rect 137134 199474 137140 199476
rect 135253 199472 137140 199474
rect 135253 199416 135258 199472
rect 135314 199416 137140 199472
rect 135253 199414 137140 199416
rect 135253 199411 135319 199414
rect 137134 199412 137140 199414
rect 137204 199412 137210 199476
rect 141141 199474 141207 199477
rect 141601 199474 141667 199477
rect 141141 199472 141667 199474
rect 141141 199416 141146 199472
rect 141202 199416 141606 199472
rect 141662 199416 141667 199472
rect 141141 199414 141667 199416
rect 141141 199411 141207 199414
rect 141601 199411 141667 199414
rect 142613 199472 142722 199477
rect 142613 199416 142618 199472
rect 142674 199416 142722 199472
rect 142613 199414 142722 199416
rect 142613 199411 142679 199414
rect 142838 199412 142844 199476
rect 142908 199474 142914 199476
rect 143073 199474 143139 199477
rect 142908 199472 143139 199474
rect 142908 199416 143078 199472
rect 143134 199416 143139 199472
rect 142908 199414 143139 199416
rect 143214 199474 143274 199550
rect 143349 199608 143458 199613
rect 143349 199552 143354 199608
rect 143410 199552 143458 199608
rect 143349 199550 143458 199552
rect 143950 199686 144148 199746
rect 143950 199613 144010 199686
rect 143950 199608 144059 199613
rect 143950 199552 143998 199608
rect 144054 199552 144059 199608
rect 143950 199550 144059 199552
rect 143349 199547 143415 199550
rect 143993 199547 144059 199550
rect 144177 199610 144243 199613
rect 144364 199610 144424 199856
rect 145143 199914 145209 199919
rect 145511 199916 145577 199919
rect 145143 199858 145148 199914
rect 145204 199858 145209 199914
rect 145143 199853 145209 199858
rect 145330 199914 145577 199916
rect 145330 199858 145516 199914
rect 145572 199858 145577 199914
rect 146523 199914 146589 199919
rect 146523 199882 146528 199914
rect 145330 199856 145577 199858
rect 145146 199749 145206 199853
rect 145097 199744 145206 199749
rect 145097 199688 145102 199744
rect 145158 199688 145206 199744
rect 145097 199686 145206 199688
rect 145097 199683 145163 199686
rect 144177 199608 144424 199610
rect 144177 199552 144182 199608
rect 144238 199552 144424 199608
rect 144177 199550 144424 199552
rect 144177 199547 144243 199550
rect 143809 199474 143875 199477
rect 143214 199472 143875 199474
rect 143214 199416 143814 199472
rect 143870 199416 143875 199472
rect 143214 199414 143875 199416
rect 145330 199474 145390 199856
rect 145511 199853 145577 199856
rect 145836 199858 146528 199882
rect 146584 199858 146589 199914
rect 146707 199914 146773 199919
rect 146707 199884 146712 199914
rect 146768 199884 146773 199914
rect 146891 199914 146957 199919
rect 145836 199853 146589 199858
rect 145836 199822 146586 199853
rect 145836 199613 145896 199822
rect 146702 199820 146708 199884
rect 146772 199882 146778 199884
rect 146772 199822 146830 199882
rect 146891 199858 146896 199914
rect 146952 199858 146957 199914
rect 147259 199914 147325 199919
rect 147259 199884 147264 199914
rect 147320 199884 147325 199914
rect 147443 199914 147509 199919
rect 146891 199853 146957 199858
rect 146772 199820 146778 199822
rect 146894 199749 146954 199853
rect 147254 199820 147260 199884
rect 147324 199882 147330 199884
rect 147324 199822 147382 199882
rect 147443 199858 147448 199914
rect 147504 199858 147509 199914
rect 147443 199853 147509 199858
rect 147627 199914 147693 199919
rect 147627 199858 147632 199914
rect 147688 199858 147693 199914
rect 147627 199853 147693 199858
rect 147903 199916 147969 199919
rect 147903 199914 148196 199916
rect 147903 199858 147908 199914
rect 147964 199884 148196 199914
rect 148547 199914 148613 199919
rect 147964 199858 148180 199884
rect 147903 199856 148180 199858
rect 147903 199853 147969 199856
rect 147324 199820 147330 199822
rect 146845 199744 146954 199749
rect 146845 199688 146850 199744
rect 146906 199688 146954 199744
rect 146845 199686 146954 199688
rect 146845 199683 146911 199686
rect 145833 199608 145899 199613
rect 145833 199552 145838 199608
rect 145894 199552 145899 199608
rect 145833 199547 145899 199552
rect 146518 199548 146524 199612
rect 146588 199610 146594 199612
rect 147446 199610 147506 199853
rect 146588 199550 147506 199610
rect 147630 199613 147690 199853
rect 148136 199822 148180 199856
rect 148174 199820 148180 199822
rect 148244 199820 148250 199884
rect 148547 199858 148552 199914
rect 148608 199858 148613 199914
rect 148547 199853 148613 199858
rect 148731 199914 148797 199919
rect 148731 199858 148736 199914
rect 148792 199858 148797 199914
rect 149375 199916 149441 199919
rect 149559 199916 149625 199919
rect 150111 199916 150177 199919
rect 149375 199914 149484 199916
rect 149375 199882 149380 199914
rect 148731 199853 148797 199858
rect 149286 199858 149380 199882
rect 149436 199858 149484 199914
rect 147903 199780 147969 199783
rect 147903 199778 148012 199780
rect 147903 199722 147908 199778
rect 147964 199746 148012 199778
rect 147964 199722 148242 199746
rect 147903 199717 148242 199722
rect 147952 199686 148242 199717
rect 147630 199608 147739 199613
rect 147630 199552 147678 199608
rect 147734 199552 147739 199608
rect 147630 199550 147739 199552
rect 146588 199548 146594 199550
rect 147673 199547 147739 199550
rect 145465 199474 145531 199477
rect 145330 199472 145531 199474
rect 145330 199416 145470 199472
rect 145526 199416 145531 199472
rect 145330 199414 145531 199416
rect 142908 199412 142914 199414
rect 143073 199411 143139 199414
rect 143809 199411 143875 199414
rect 145465 199411 145531 199414
rect 147765 199474 147831 199477
rect 148182 199474 148242 199686
rect 148550 199613 148610 199853
rect 148734 199749 148794 199853
rect 148685 199744 148794 199749
rect 148685 199688 148690 199744
rect 148746 199688 148794 199744
rect 148685 199686 148794 199688
rect 149286 199822 149484 199858
rect 149559 199914 149760 199916
rect 149559 199858 149564 199914
rect 149620 199858 149760 199914
rect 149559 199856 149760 199858
rect 149559 199853 149625 199856
rect 148685 199683 148751 199686
rect 148501 199608 148610 199613
rect 148501 199552 148506 199608
rect 148562 199552 148610 199608
rect 148501 199550 148610 199552
rect 149286 199613 149346 199822
rect 149286 199608 149395 199613
rect 149286 199552 149334 199608
rect 149390 199552 149395 199608
rect 149286 199550 149395 199552
rect 148501 199547 148567 199550
rect 149329 199547 149395 199550
rect 149513 199610 149579 199613
rect 149700 199610 149760 199856
rect 149976 199914 150177 199916
rect 149976 199858 150116 199914
rect 150172 199858 150177 199914
rect 150755 199914 150821 199919
rect 149976 199856 150177 199858
rect 149976 199613 150036 199856
rect 150111 199853 150177 199856
rect 150387 199880 150453 199885
rect 150387 199824 150392 199880
rect 150448 199824 150453 199880
rect 150755 199858 150760 199914
rect 150816 199858 150821 199914
rect 150755 199853 150821 199858
rect 150387 199819 150453 199824
rect 150390 199746 150450 199819
rect 150617 199746 150683 199749
rect 150390 199744 150683 199746
rect 150390 199688 150622 199744
rect 150678 199688 150683 199744
rect 150390 199686 150683 199688
rect 150617 199683 150683 199686
rect 149513 199608 149760 199610
rect 149513 199552 149518 199608
rect 149574 199552 149760 199608
rect 149513 199550 149760 199552
rect 149973 199608 150039 199613
rect 149973 199552 149978 199608
rect 150034 199552 150039 199608
rect 149513 199547 149579 199550
rect 149973 199547 150039 199552
rect 147765 199472 148242 199474
rect 147765 199416 147770 199472
rect 147826 199416 148242 199472
rect 147765 199414 148242 199416
rect 149697 199474 149763 199477
rect 150758 199474 150818 199853
rect 150988 199610 151048 200094
rect 154530 200094 154804 200154
rect 154530 199919 154590 200094
rect 154798 200092 154804 200094
rect 154868 200092 154874 200156
rect 151951 199916 152017 199919
rect 153239 199916 153305 199919
rect 151951 199914 152060 199916
rect 151491 199884 151557 199885
rect 151486 199882 151492 199884
rect 151400 199822 151492 199882
rect 151486 199820 151492 199822
rect 151556 199820 151562 199884
rect 151951 199858 151956 199914
rect 152012 199882 152060 199914
rect 153196 199914 153305 199916
rect 153196 199884 153244 199914
rect 152958 199882 152964 199884
rect 152012 199858 152964 199882
rect 151951 199853 152964 199858
rect 152000 199822 152964 199853
rect 152958 199820 152964 199822
rect 153028 199820 153034 199884
rect 153142 199820 153148 199884
rect 153212 199858 153244 199884
rect 153300 199858 153305 199914
rect 153515 199914 153581 199919
rect 153515 199884 153520 199914
rect 153576 199884 153581 199914
rect 153791 199916 153857 199919
rect 153791 199914 153900 199916
rect 153212 199853 153305 199858
rect 153212 199822 153256 199853
rect 153212 199820 153218 199822
rect 153510 199820 153516 199884
rect 153580 199882 153586 199884
rect 153580 199822 153638 199882
rect 153791 199858 153796 199914
rect 153852 199884 153900 199914
rect 154527 199914 154593 199919
rect 154895 199916 154961 199919
rect 153852 199858 153884 199884
rect 153791 199853 153884 199858
rect 153840 199822 153884 199853
rect 153580 199820 153586 199822
rect 153878 199820 153884 199822
rect 153948 199820 153954 199884
rect 154527 199858 154532 199914
rect 154588 199858 154593 199914
rect 154527 199853 154593 199858
rect 154852 199914 154961 199916
rect 154852 199858 154900 199914
rect 154956 199882 154961 199914
rect 155447 199916 155513 199919
rect 155447 199914 155648 199916
rect 155166 199882 155172 199884
rect 154956 199858 155172 199882
rect 154852 199822 155172 199858
rect 155166 199820 155172 199822
rect 155236 199820 155242 199884
rect 155447 199858 155452 199914
rect 155508 199858 155648 199914
rect 155907 199914 155973 199919
rect 155447 199856 155648 199858
rect 155447 199853 155513 199856
rect 151491 199819 151557 199820
rect 151670 199684 151676 199748
rect 151740 199746 151746 199748
rect 154113 199746 154179 199749
rect 151740 199744 154179 199746
rect 151740 199688 154118 199744
rect 154174 199688 154179 199744
rect 151740 199686 154179 199688
rect 151740 199684 151746 199686
rect 154113 199683 154179 199686
rect 155401 199746 155467 199749
rect 155588 199746 155648 199856
rect 155723 199880 155789 199885
rect 155723 199824 155728 199880
rect 155784 199824 155789 199880
rect 155907 199858 155912 199914
rect 155968 199858 155973 199914
rect 155907 199853 155973 199858
rect 156091 199914 156157 199919
rect 156091 199858 156096 199914
rect 156152 199858 156157 199914
rect 156091 199853 156157 199858
rect 155723 199819 155789 199824
rect 155401 199744 155648 199746
rect 155401 199688 155406 199744
rect 155462 199688 155648 199744
rect 155401 199686 155648 199688
rect 155401 199683 155467 199686
rect 154527 199642 154593 199647
rect 153101 199610 153167 199613
rect 150988 199608 153167 199610
rect 150988 199552 153106 199608
rect 153162 199552 153167 199608
rect 150988 199550 153167 199552
rect 153101 199547 153167 199550
rect 153326 199548 153332 199612
rect 153396 199610 153402 199612
rect 153469 199610 153535 199613
rect 153396 199608 153535 199610
rect 153396 199552 153474 199608
rect 153530 199552 153535 199608
rect 153396 199550 153535 199552
rect 153396 199548 153402 199550
rect 153469 199547 153535 199550
rect 153929 199610 153995 199613
rect 154527 199610 154532 199642
rect 153929 199608 154532 199610
rect 153929 199552 153934 199608
rect 153990 199586 154532 199608
rect 154588 199586 154593 199642
rect 155726 199613 155786 199819
rect 155910 199749 155970 199853
rect 156094 199749 156154 199853
rect 156462 199749 156522 200366
rect 180333 200424 208735 200426
rect 180333 200368 180338 200424
rect 180394 200368 208674 200424
rect 208730 200368 208735 200424
rect 180333 200366 208735 200368
rect 180333 200363 180399 200366
rect 208669 200363 208735 200366
rect 168414 200228 168420 200292
rect 168484 200290 168490 200292
rect 201585 200290 201651 200293
rect 168484 200288 201651 200290
rect 168484 200232 201590 200288
rect 201646 200232 201651 200288
rect 168484 200230 201651 200232
rect 168484 200228 168490 200230
rect 201585 200227 201651 200230
rect 166390 200092 166396 200156
rect 166460 200154 166466 200156
rect 201125 200154 201191 200157
rect 166460 200152 201191 200154
rect 166460 200096 201130 200152
rect 201186 200096 201191 200152
rect 166460 200094 201191 200096
rect 166460 200092 166466 200094
rect 201125 200091 201191 200094
rect 169518 200018 169524 200020
rect 169296 199958 169524 200018
rect 156643 199914 156709 199919
rect 157103 199916 157169 199919
rect 156643 199884 156648 199914
rect 156704 199884 156709 199914
rect 157060 199914 157169 199916
rect 156638 199820 156644 199884
rect 156708 199882 156714 199884
rect 156708 199822 156766 199882
rect 157060 199858 157108 199914
rect 157164 199858 157169 199914
rect 157747 199914 157813 199919
rect 157747 199884 157752 199914
rect 157808 199884 157813 199914
rect 159495 199916 159561 199919
rect 159863 199916 159929 199919
rect 159495 199914 159604 199916
rect 157060 199853 157169 199858
rect 156708 199820 156714 199822
rect 156827 199778 156893 199783
rect 155910 199744 156019 199749
rect 155910 199688 155958 199744
rect 156014 199688 156019 199744
rect 155910 199686 156019 199688
rect 156094 199744 156203 199749
rect 156094 199688 156142 199744
rect 156198 199688 156203 199744
rect 156094 199686 156203 199688
rect 155953 199683 156019 199686
rect 156137 199683 156203 199686
rect 156459 199744 156525 199749
rect 156459 199688 156464 199744
rect 156520 199688 156525 199744
rect 156459 199683 156525 199688
rect 156597 199746 156663 199749
rect 156827 199746 156832 199778
rect 156597 199744 156832 199746
rect 156597 199688 156602 199744
rect 156658 199722 156832 199744
rect 156888 199722 156893 199778
rect 156658 199717 156893 199722
rect 156658 199688 156890 199717
rect 156597 199686 156890 199688
rect 156597 199683 156663 199686
rect 153990 199581 154593 199586
rect 155585 199608 155651 199613
rect 153990 199552 154590 199581
rect 153929 199550 154590 199552
rect 155585 199552 155590 199608
rect 155646 199552 155651 199608
rect 153929 199547 153995 199550
rect 155585 199547 155651 199552
rect 155726 199608 155835 199613
rect 155726 199552 155774 199608
rect 155830 199552 155835 199608
rect 155726 199550 155835 199552
rect 155769 199547 155835 199550
rect 156781 199610 156847 199613
rect 157060 199610 157120 199853
rect 157742 199820 157748 199884
rect 157812 199882 157818 199884
rect 157812 199822 157870 199882
rect 159495 199858 159500 199914
rect 159556 199858 159604 199914
rect 159495 199853 159604 199858
rect 159863 199914 159972 199916
rect 159863 199858 159868 199914
rect 159924 199882 159972 199914
rect 160323 199914 160389 199919
rect 160134 199882 160140 199884
rect 159924 199858 160140 199882
rect 159863 199853 160140 199858
rect 157812 199820 157818 199822
rect 157195 199778 157261 199783
rect 157195 199748 157200 199778
rect 157256 199748 157261 199778
rect 157190 199684 157196 199748
rect 157260 199746 157266 199748
rect 157260 199686 157318 199746
rect 157260 199684 157266 199686
rect 157558 199684 157564 199748
rect 157628 199746 157634 199748
rect 158023 199746 158089 199749
rect 158437 199746 158503 199749
rect 157628 199744 158089 199746
rect 157628 199688 158028 199744
rect 158084 199688 158089 199744
rect 157628 199686 158089 199688
rect 157628 199684 157634 199686
rect 158023 199683 158089 199686
rect 158164 199744 158503 199746
rect 158164 199688 158442 199744
rect 158498 199688 158503 199744
rect 158164 199686 158503 199688
rect 156781 199608 157120 199610
rect 156781 199552 156786 199608
rect 156842 199552 157120 199608
rect 156781 199550 157120 199552
rect 157517 199610 157583 199613
rect 157977 199610 158043 199613
rect 157517 199608 158043 199610
rect 157517 199552 157522 199608
rect 157578 199552 157982 199608
rect 158038 199552 158043 199608
rect 157517 199550 158043 199552
rect 156781 199547 156847 199550
rect 157517 199547 157583 199550
rect 157977 199547 158043 199550
rect 149697 199472 150818 199474
rect 149697 199416 149702 199472
rect 149758 199416 150818 199472
rect 149697 199414 150818 199416
rect 154573 199476 154639 199477
rect 154573 199472 154620 199476
rect 154684 199474 154690 199476
rect 154573 199416 154578 199472
rect 147765 199411 147831 199414
rect 149697 199411 149763 199414
rect 154573 199412 154620 199416
rect 154684 199414 154730 199474
rect 154684 199412 154690 199414
rect 154573 199411 154639 199412
rect 118550 199276 118556 199340
rect 118620 199338 118626 199340
rect 151077 199338 151143 199341
rect 118620 199336 151143 199338
rect 118620 199280 151082 199336
rect 151138 199280 151143 199336
rect 118620 199278 151143 199280
rect 155588 199338 155648 199547
rect 156413 199474 156479 199477
rect 158164 199474 158224 199686
rect 158437 199683 158503 199686
rect 158989 199608 159055 199613
rect 158989 199552 158994 199608
rect 159050 199552 159055 199608
rect 158989 199547 159055 199552
rect 158992 199477 159052 199547
rect 156413 199472 158224 199474
rect 156413 199416 156418 199472
rect 156474 199416 158224 199472
rect 156413 199414 158224 199416
rect 158989 199472 159055 199477
rect 158989 199416 158994 199472
rect 159050 199416 159055 199472
rect 156413 199411 156479 199414
rect 158989 199411 159055 199416
rect 159544 199338 159604 199853
rect 159912 199822 160140 199853
rect 160134 199820 160140 199822
rect 160204 199820 160210 199884
rect 160323 199858 160328 199914
rect 160384 199858 160389 199914
rect 160323 199853 160389 199858
rect 160507 199914 160573 199919
rect 160507 199858 160512 199914
rect 160568 199858 160573 199914
rect 160507 199853 160573 199858
rect 160783 199914 160849 199919
rect 161335 199916 161401 199919
rect 160783 199858 160788 199914
rect 160844 199858 160849 199914
rect 161108 199914 161401 199916
rect 161108 199884 161340 199914
rect 160783 199853 160849 199858
rect 160326 199613 160386 199853
rect 160510 199613 160570 199853
rect 160786 199749 160846 199853
rect 161054 199820 161060 199884
rect 161124 199858 161340 199884
rect 161396 199858 161401 199914
rect 161124 199856 161401 199858
rect 161124 199822 161168 199856
rect 161335 199853 161401 199856
rect 161611 199914 161677 199919
rect 162071 199916 162137 199919
rect 161611 199858 161616 199914
rect 161672 199858 161677 199914
rect 161936 199914 162137 199916
rect 161611 199853 161677 199858
rect 161124 199820 161130 199822
rect 161473 199780 161539 199783
rect 161430 199778 161539 199780
rect 160786 199744 160895 199749
rect 161197 199748 161263 199749
rect 161430 199748 161478 199778
rect 161197 199746 161244 199748
rect 160786 199688 160834 199744
rect 160890 199688 160895 199744
rect 160786 199686 160895 199688
rect 161152 199744 161244 199746
rect 161152 199688 161202 199744
rect 161152 199686 161244 199688
rect 160829 199683 160895 199686
rect 161197 199684 161244 199686
rect 161308 199684 161314 199748
rect 161422 199746 161428 199748
rect 161416 199686 161428 199746
rect 161534 199722 161539 199778
rect 161422 199684 161428 199686
rect 161492 199717 161539 199722
rect 161492 199684 161498 199717
rect 161197 199683 161263 199684
rect 160277 199608 160386 199613
rect 160277 199552 160282 199608
rect 160338 199552 160386 199608
rect 160277 199550 160386 199552
rect 160461 199608 160570 199613
rect 160461 199552 160466 199608
rect 160522 199552 160570 199608
rect 160461 199550 160570 199552
rect 161013 199610 161079 199613
rect 161614 199610 161674 199853
rect 161790 199820 161796 199884
rect 161860 199882 161866 199884
rect 161936 199882 162076 199914
rect 161860 199858 162076 199882
rect 162132 199858 162137 199914
rect 161860 199856 162137 199858
rect 161860 199822 161996 199856
rect 162071 199853 162137 199856
rect 162255 199914 162321 199919
rect 162255 199858 162260 199914
rect 162316 199858 162321 199914
rect 162255 199853 162321 199858
rect 162899 199914 162965 199919
rect 162899 199858 162904 199914
rect 162960 199858 162965 199914
rect 163451 199914 163517 199919
rect 162899 199853 162965 199858
rect 161860 199820 161866 199822
rect 162258 199749 162318 199853
rect 162209 199744 162318 199749
rect 162209 199688 162214 199744
rect 162270 199688 162318 199744
rect 162209 199686 162318 199688
rect 162209 199683 162275 199686
rect 162902 199613 162962 199853
rect 163078 199820 163084 199884
rect 163148 199882 163154 199884
rect 163451 199882 163456 199914
rect 163148 199858 163456 199882
rect 163512 199858 163517 199914
rect 164095 199914 164161 199919
rect 163148 199853 163517 199858
rect 163148 199822 163514 199853
rect 163148 199820 163154 199822
rect 163814 199820 163820 199884
rect 163884 199882 163890 199884
rect 164095 199882 164100 199914
rect 163884 199858 164100 199882
rect 164156 199858 164161 199914
rect 163884 199853 164161 199858
rect 164371 199914 164437 199919
rect 165199 199916 165265 199919
rect 164371 199858 164376 199914
rect 164432 199858 164437 199914
rect 164972 199914 165265 199916
rect 164972 199884 165204 199914
rect 164371 199853 164437 199858
rect 163884 199822 164158 199853
rect 163884 199820 163890 199822
rect 163635 199778 163701 199783
rect 163497 199748 163563 199749
rect 163635 199748 163640 199778
rect 163696 199748 163701 199778
rect 163446 199746 163452 199748
rect 163406 199686 163452 199746
rect 163516 199744 163563 199748
rect 163558 199688 163563 199744
rect 163446 199684 163452 199686
rect 163516 199684 163563 199688
rect 163630 199684 163636 199748
rect 163700 199746 163706 199748
rect 163700 199686 163758 199746
rect 163700 199684 163706 199686
rect 163497 199683 163563 199684
rect 161013 199608 161674 199610
rect 161013 199552 161018 199608
rect 161074 199552 161674 199608
rect 161013 199550 161674 199552
rect 162393 199610 162459 199613
rect 162526 199610 162532 199612
rect 162393 199608 162532 199610
rect 162393 199552 162398 199608
rect 162454 199552 162532 199608
rect 162393 199550 162532 199552
rect 160277 199547 160343 199550
rect 160461 199547 160527 199550
rect 161013 199547 161079 199550
rect 162393 199547 162459 199550
rect 162526 199548 162532 199550
rect 162596 199548 162602 199612
rect 162902 199608 163011 199613
rect 162902 199552 162950 199608
rect 163006 199552 163011 199608
rect 162902 199550 163011 199552
rect 162945 199547 163011 199550
rect 163262 199548 163268 199612
rect 163332 199610 163338 199612
rect 163957 199610 164023 199613
rect 163332 199608 164023 199610
rect 163332 199552 163962 199608
rect 164018 199552 164023 199608
rect 163332 199550 164023 199552
rect 163332 199548 163338 199550
rect 163957 199547 164023 199550
rect 161238 199412 161244 199476
rect 161308 199474 161314 199476
rect 161565 199474 161631 199477
rect 163681 199476 163747 199477
rect 161308 199472 161631 199474
rect 161308 199416 161570 199472
rect 161626 199416 161631 199472
rect 161308 199414 161631 199416
rect 161308 199412 161314 199414
rect 161565 199411 161631 199414
rect 163630 199412 163636 199476
rect 163700 199474 163747 199476
rect 164374 199474 164434 199853
rect 164918 199820 164924 199884
rect 164988 199858 165204 199884
rect 165260 199858 165265 199914
rect 164988 199856 165265 199858
rect 164988 199822 165032 199856
rect 165199 199853 165265 199856
rect 165567 199916 165633 199919
rect 165567 199914 165860 199916
rect 165567 199858 165572 199914
rect 165628 199884 165860 199914
rect 166027 199914 166093 199919
rect 166027 199884 166032 199914
rect 166088 199884 166093 199914
rect 166303 199916 166369 199919
rect 166303 199914 166642 199916
rect 165628 199858 165844 199884
rect 165567 199856 165844 199858
rect 165567 199853 165633 199856
rect 165800 199822 165844 199856
rect 164988 199820 164994 199822
rect 165838 199820 165844 199822
rect 165908 199820 165914 199884
rect 166022 199820 166028 199884
rect 166092 199882 166098 199884
rect 166092 199822 166150 199882
rect 166303 199858 166308 199914
rect 166364 199884 166642 199914
rect 167131 199914 167197 199919
rect 166364 199858 166580 199884
rect 166303 199856 166580 199858
rect 166303 199853 166369 199856
rect 166092 199820 166098 199822
rect 166574 199820 166580 199856
rect 166644 199820 166650 199884
rect 167131 199858 167136 199914
rect 167192 199882 167197 199914
rect 167867 199914 167933 199919
rect 167494 199882 167500 199884
rect 167192 199858 167500 199882
rect 167131 199853 167500 199858
rect 167134 199822 167500 199853
rect 167494 199820 167500 199822
rect 167564 199820 167570 199884
rect 167678 199820 167684 199884
rect 167748 199882 167754 199884
rect 167867 199882 167872 199914
rect 167748 199858 167872 199882
rect 167928 199858 167933 199914
rect 167748 199853 167933 199858
rect 168051 199914 168117 199919
rect 168051 199858 168056 199914
rect 168112 199858 168117 199914
rect 168051 199853 168117 199858
rect 168327 199916 168393 199919
rect 168327 199914 168436 199916
rect 168327 199858 168332 199914
rect 168388 199882 168436 199914
rect 168971 199914 169037 199919
rect 168598 199882 168604 199884
rect 168388 199858 168604 199882
rect 168327 199853 168604 199858
rect 167748 199822 167930 199853
rect 167748 199820 167754 199822
rect 164601 199746 164667 199749
rect 164734 199746 164740 199748
rect 164601 199744 164740 199746
rect 164601 199688 164606 199744
rect 164662 199688 164740 199744
rect 164601 199686 164740 199688
rect 164601 199683 164667 199686
rect 164734 199684 164740 199686
rect 164804 199684 164810 199748
rect 164877 199746 164943 199749
rect 165153 199746 165219 199749
rect 164877 199744 165219 199746
rect 164877 199688 164882 199744
rect 164938 199688 165158 199744
rect 165214 199688 165219 199744
rect 164877 199686 165219 199688
rect 164877 199683 164943 199686
rect 165153 199683 165219 199686
rect 165286 199684 165292 199748
rect 165356 199746 165362 199748
rect 165751 199746 165817 199749
rect 165356 199744 165817 199746
rect 165356 199688 165756 199744
rect 165812 199688 165817 199744
rect 165356 199686 165817 199688
rect 165356 199684 165362 199686
rect 165751 199683 165817 199686
rect 166947 199744 167013 199749
rect 166947 199688 166952 199744
rect 167008 199688 167013 199744
rect 166947 199683 167013 199688
rect 164509 199610 164575 199613
rect 166950 199610 167010 199683
rect 168054 199613 168114 199853
rect 168376 199822 168604 199853
rect 168598 199820 168604 199822
rect 168668 199820 168674 199884
rect 168782 199820 168788 199884
rect 168852 199882 168858 199884
rect 168971 199882 168976 199914
rect 168852 199858 168976 199882
rect 169032 199858 169037 199914
rect 168852 199853 169037 199858
rect 169155 199914 169221 199919
rect 169155 199858 169160 199914
rect 169216 199882 169221 199914
rect 169296 199882 169356 199958
rect 169518 199956 169524 199958
rect 169588 199956 169594 200020
rect 170806 199956 170812 200020
rect 170876 200018 170882 200020
rect 170876 199958 171012 200018
rect 170876 199956 170882 199958
rect 169707 199914 169773 199919
rect 169707 199882 169712 199914
rect 169216 199858 169356 199882
rect 169155 199853 169356 199858
rect 168852 199822 169034 199853
rect 169158 199822 169356 199853
rect 169434 199858 169712 199882
rect 169768 199858 169773 199914
rect 169891 199914 169957 199919
rect 169891 199884 169896 199914
rect 169952 199884 169957 199914
rect 170075 199914 170141 199919
rect 169434 199853 169773 199858
rect 169434 199822 169770 199853
rect 168852 199820 168858 199822
rect 168603 199744 168669 199749
rect 168603 199688 168608 199744
rect 168664 199688 168669 199744
rect 168603 199683 168669 199688
rect 168741 199746 168807 199749
rect 168741 199744 169034 199746
rect 168741 199688 168746 199744
rect 168802 199688 169034 199744
rect 168741 199686 169034 199688
rect 168741 199683 168807 199686
rect 167821 199610 167887 199613
rect 164509 199608 166826 199610
rect 164509 199552 164514 199608
rect 164570 199552 166826 199608
rect 164509 199550 166826 199552
rect 166950 199608 167887 199610
rect 166950 199552 167826 199608
rect 167882 199552 167887 199608
rect 166950 199550 167887 199552
rect 164509 199547 164575 199550
rect 165245 199474 165311 199477
rect 163700 199472 163792 199474
rect 163742 199416 163792 199472
rect 163700 199414 163792 199416
rect 164374 199472 165311 199474
rect 164374 199416 165250 199472
rect 165306 199416 165311 199472
rect 164374 199414 165311 199416
rect 163700 199412 163747 199414
rect 163681 199411 163747 199412
rect 165245 199411 165311 199414
rect 165889 199474 165955 199477
rect 166390 199474 166396 199476
rect 165889 199472 166396 199474
rect 165889 199416 165894 199472
rect 165950 199416 166396 199472
rect 165889 199414 166396 199416
rect 165889 199411 165955 199414
rect 166390 199412 166396 199414
rect 166460 199412 166466 199476
rect 166766 199474 166826 199550
rect 167821 199547 167887 199550
rect 168005 199608 168114 199613
rect 168465 199612 168531 199613
rect 168414 199610 168420 199612
rect 168005 199552 168010 199608
rect 168066 199552 168114 199608
rect 168005 199550 168114 199552
rect 168374 199550 168420 199610
rect 168484 199608 168531 199612
rect 168526 199552 168531 199608
rect 168005 199547 168071 199550
rect 168414 199548 168420 199550
rect 168484 199548 168531 199552
rect 168606 199610 168666 199683
rect 168741 199610 168807 199613
rect 168606 199608 168807 199610
rect 168606 199552 168746 199608
rect 168802 199552 168807 199608
rect 168606 199550 168807 199552
rect 168465 199547 168531 199548
rect 168741 199547 168807 199550
rect 167085 199474 167151 199477
rect 166766 199472 167151 199474
rect 166766 199416 167090 199472
rect 167146 199416 167151 199472
rect 166766 199414 167151 199416
rect 167085 199411 167151 199414
rect 168649 199474 168715 199477
rect 168974 199474 169034 199686
rect 169109 199612 169175 199613
rect 169109 199608 169156 199612
rect 169220 199610 169226 199612
rect 169434 199610 169494 199822
rect 169886 199820 169892 199884
rect 169956 199882 169962 199884
rect 169956 199822 170014 199882
rect 170075 199858 170080 199914
rect 170136 199858 170141 199914
rect 170075 199853 170141 199858
rect 170259 199914 170325 199919
rect 170259 199858 170264 199914
rect 170320 199858 170325 199914
rect 170627 199914 170693 199919
rect 170627 199884 170632 199914
rect 170688 199884 170693 199914
rect 170259 199853 170325 199858
rect 169956 199820 169962 199822
rect 169707 199746 169773 199749
rect 170078 199748 170138 199853
rect 169707 199744 170000 199746
rect 169707 199688 169712 199744
rect 169768 199688 170000 199744
rect 169707 199686 170000 199688
rect 169707 199683 169773 199686
rect 169661 199610 169727 199613
rect 169109 199552 169114 199608
rect 169109 199548 169156 199552
rect 169220 199550 169266 199610
rect 169434 199608 169727 199610
rect 169434 199552 169666 199608
rect 169722 199552 169727 199608
rect 169434 199550 169727 199552
rect 169940 199610 170000 199686
rect 170070 199684 170076 199748
rect 170140 199684 170146 199748
rect 170121 199610 170187 199613
rect 169940 199608 170187 199610
rect 169940 199552 170126 199608
rect 170182 199552 170187 199608
rect 169940 199550 170187 199552
rect 169220 199548 169226 199550
rect 169109 199547 169175 199548
rect 169661 199547 169727 199550
rect 170121 199547 170187 199550
rect 169334 199474 169340 199476
rect 168649 199472 168850 199474
rect 168649 199416 168654 199472
rect 168710 199416 168850 199472
rect 168649 199414 168850 199416
rect 168974 199414 169340 199474
rect 168649 199411 168715 199414
rect 163681 199338 163747 199341
rect 163957 199338 164023 199341
rect 155588 199278 156522 199338
rect 159544 199336 163747 199338
rect 159544 199280 163686 199336
rect 163742 199280 163747 199336
rect 159544 199278 163747 199280
rect 118620 199276 118626 199278
rect 151077 199275 151143 199278
rect 107193 199202 107259 199205
rect 135253 199202 135319 199205
rect 107193 199200 135319 199202
rect 107193 199144 107198 199200
rect 107254 199144 135258 199200
rect 135314 199144 135319 199200
rect 107193 199142 135319 199144
rect 107193 199139 107259 199142
rect 135253 199139 135319 199142
rect 135478 199140 135484 199204
rect 135548 199202 135554 199204
rect 135897 199202 135963 199205
rect 136357 199204 136423 199205
rect 136357 199202 136404 199204
rect 135548 199200 135963 199202
rect 135548 199144 135902 199200
rect 135958 199144 135963 199200
rect 135548 199142 135963 199144
rect 136312 199200 136404 199202
rect 136312 199144 136362 199200
rect 136312 199142 136404 199144
rect 135548 199140 135554 199142
rect 135897 199139 135963 199142
rect 136357 199140 136404 199142
rect 136468 199140 136474 199204
rect 136582 199140 136588 199204
rect 136652 199202 136658 199204
rect 138289 199202 138355 199205
rect 136652 199200 138355 199202
rect 136652 199144 138294 199200
rect 138350 199144 138355 199200
rect 136652 199142 138355 199144
rect 136652 199140 136658 199142
rect 136357 199139 136423 199140
rect 138289 199139 138355 199142
rect 139393 199202 139459 199205
rect 147029 199202 147095 199205
rect 139393 199200 147095 199202
rect 139393 199144 139398 199200
rect 139454 199144 147034 199200
rect 147090 199144 147095 199200
rect 139393 199142 147095 199144
rect 139393 199139 139459 199142
rect 147029 199139 147095 199142
rect 152641 199202 152707 199205
rect 156462 199202 156522 199278
rect 163681 199275 163747 199278
rect 163822 199336 164023 199338
rect 163822 199280 163962 199336
rect 164018 199280 164023 199336
rect 163822 199278 164023 199280
rect 162393 199202 162459 199205
rect 152641 199200 156338 199202
rect 152641 199144 152646 199200
rect 152702 199144 156338 199200
rect 152641 199142 156338 199144
rect 156462 199200 162459 199202
rect 156462 199144 162398 199200
rect 162454 199144 162459 199200
rect 156462 199142 162459 199144
rect 152641 199139 152707 199142
rect 127893 199066 127959 199069
rect 155953 199066 156019 199069
rect 127893 199064 156019 199066
rect 127893 199008 127898 199064
rect 127954 199008 155958 199064
rect 156014 199008 156019 199064
rect 127893 199006 156019 199008
rect 127893 199003 127959 199006
rect 155953 199003 156019 199006
rect 128077 198930 128143 198933
rect 153653 198930 153719 198933
rect 128077 198928 153719 198930
rect 128077 198872 128082 198928
rect 128138 198872 153658 198928
rect 153714 198872 153719 198928
rect 128077 198870 153719 198872
rect 128077 198867 128143 198870
rect 153653 198867 153719 198870
rect 131849 198794 131915 198797
rect 137185 198794 137251 198797
rect 131849 198792 137251 198794
rect 131849 198736 131854 198792
rect 131910 198736 137190 198792
rect 137246 198736 137251 198792
rect 131849 198734 137251 198736
rect 131849 198731 131915 198734
rect 137185 198731 137251 198734
rect 141233 198794 141299 198797
rect 141417 198794 141483 198797
rect 141877 198796 141943 198797
rect 141877 198794 141924 198796
rect 141233 198792 141483 198794
rect 141233 198736 141238 198792
rect 141294 198736 141422 198792
rect 141478 198736 141483 198792
rect 141233 198734 141483 198736
rect 141832 198792 141924 198794
rect 141832 198736 141882 198792
rect 141832 198734 141924 198736
rect 141233 198731 141299 198734
rect 141417 198731 141483 198734
rect 141877 198732 141924 198734
rect 141988 198732 141994 198796
rect 142061 198794 142127 198797
rect 143073 198796 143139 198797
rect 142654 198794 142660 198796
rect 142061 198792 142660 198794
rect 142061 198736 142066 198792
rect 142122 198736 142660 198792
rect 142061 198734 142660 198736
rect 141877 198731 141943 198732
rect 142061 198731 142127 198734
rect 142654 198732 142660 198734
rect 142724 198732 142730 198796
rect 143022 198732 143028 198796
rect 143092 198794 143139 198796
rect 156278 198794 156338 199142
rect 162393 199139 162459 199142
rect 157793 199066 157859 199069
rect 163589 199066 163655 199069
rect 157793 199064 163655 199066
rect 157793 199008 157798 199064
rect 157854 199008 163594 199064
rect 163650 199008 163655 199064
rect 157793 199006 163655 199008
rect 157793 199003 157859 199006
rect 163589 199003 163655 199006
rect 157149 198930 157215 198933
rect 163822 198930 163882 199278
rect 163957 199275 164023 199278
rect 166073 199338 166139 199341
rect 168649 199338 168715 199341
rect 166073 199336 168715 199338
rect 166073 199280 166078 199336
rect 166134 199280 168654 199336
rect 168710 199280 168715 199336
rect 166073 199278 168715 199280
rect 168790 199338 168850 199414
rect 169334 199412 169340 199414
rect 169404 199412 169410 199476
rect 169702 199412 169708 199476
rect 169772 199474 169778 199476
rect 169937 199474 170003 199477
rect 169772 199472 170003 199474
rect 169772 199416 169942 199472
rect 169998 199416 170003 199472
rect 169772 199414 170003 199416
rect 170262 199474 170322 199853
rect 170622 199820 170628 199884
rect 170692 199882 170698 199884
rect 170692 199822 170750 199882
rect 170952 199851 171012 199958
rect 172830 199956 172836 200020
rect 172900 200018 172906 200020
rect 174118 200018 174124 200020
rect 172900 199958 174124 200018
rect 172900 199956 172906 199958
rect 174118 199956 174124 199958
rect 174188 199956 174194 200020
rect 171271 199916 171337 199919
rect 171915 199916 171981 199919
rect 171271 199914 171380 199916
rect 171271 199858 171276 199914
rect 171332 199884 171380 199914
rect 171872 199914 171981 199916
rect 171332 199858 171364 199884
rect 171271 199853 171364 199858
rect 170903 199846 171012 199851
rect 170692 199820 170698 199822
rect 170903 199790 170908 199846
rect 170964 199790 171012 199846
rect 171320 199822 171364 199853
rect 171358 199820 171364 199822
rect 171428 199820 171434 199884
rect 171542 199820 171548 199884
rect 171612 199882 171618 199884
rect 171872 199882 171920 199914
rect 171612 199858 171920 199882
rect 171976 199858 171981 199914
rect 172651 199914 172717 199919
rect 174399 199916 174465 199919
rect 172651 199884 172656 199914
rect 172712 199884 172717 199914
rect 174264 199914 174465 199916
rect 172462 199882 172468 199884
rect 171612 199853 171981 199858
rect 171612 199822 171932 199853
rect 172240 199822 172468 199882
rect 171612 199820 171618 199822
rect 170903 199788 171012 199790
rect 170903 199785 170969 199788
rect 172240 199749 172300 199822
rect 172462 199820 172468 199822
rect 172532 199820 172538 199884
rect 172646 199820 172652 199884
rect 172716 199882 172722 199884
rect 172927 199882 172993 199885
rect 172716 199822 172774 199882
rect 172927 199880 173036 199882
rect 172927 199824 172932 199880
rect 172988 199824 173036 199880
rect 172716 199820 172722 199822
rect 172927 199819 173036 199824
rect 173203 199880 173269 199885
rect 173203 199824 173208 199880
rect 173264 199824 173269 199880
rect 173203 199819 173269 199824
rect 173382 199820 173388 199884
rect 173452 199882 173458 199884
rect 173663 199882 173729 199885
rect 173452 199880 173729 199882
rect 173452 199824 173668 199880
rect 173724 199824 173729 199880
rect 173452 199822 173729 199824
rect 173452 199820 173458 199822
rect 173663 199819 173729 199822
rect 174264 199858 174404 199914
rect 174460 199858 174465 199914
rect 174264 199856 174465 199858
rect 171225 199746 171291 199749
rect 171726 199746 171732 199748
rect 171225 199744 171732 199746
rect 171225 199688 171230 199744
rect 171286 199688 171732 199744
rect 171225 199686 171732 199688
rect 171225 199683 171291 199686
rect 171726 199684 171732 199686
rect 171796 199684 171802 199748
rect 171910 199684 171916 199748
rect 171980 199746 171986 199748
rect 172053 199746 172119 199749
rect 171980 199744 172119 199746
rect 171980 199688 172058 199744
rect 172114 199688 172119 199744
rect 171980 199686 172119 199688
rect 171980 199684 171986 199686
rect 172053 199683 172119 199686
rect 172191 199744 172300 199749
rect 172191 199688 172196 199744
rect 172252 199688 172300 199744
rect 172191 199686 172300 199688
rect 172191 199683 172257 199686
rect 172462 199684 172468 199748
rect 172532 199746 172538 199748
rect 172605 199746 172671 199749
rect 172976 199748 173036 199819
rect 172532 199744 172671 199746
rect 172532 199688 172610 199744
rect 172666 199688 172671 199744
rect 172532 199686 172671 199688
rect 172532 199684 172538 199686
rect 172605 199683 172671 199686
rect 172968 199684 172974 199748
rect 173038 199684 173044 199748
rect 173206 199746 173266 199819
rect 174264 199748 174324 199856
rect 174399 199853 174465 199856
rect 174583 199916 174649 199919
rect 174583 199914 174922 199916
rect 174583 199858 174588 199914
rect 174644 199884 174922 199914
rect 175227 199914 175293 199919
rect 174644 199858 174860 199884
rect 174583 199856 174860 199858
rect 174583 199853 174649 199856
rect 174854 199820 174860 199856
rect 174924 199820 174930 199884
rect 175227 199858 175232 199914
rect 175288 199882 175293 199914
rect 175871 199916 175937 199919
rect 176423 199916 176489 199919
rect 175871 199914 175980 199916
rect 175406 199882 175412 199884
rect 175288 199858 175412 199882
rect 175227 199853 175412 199858
rect 175230 199822 175412 199853
rect 175406 199820 175412 199822
rect 175476 199820 175482 199884
rect 175871 199858 175876 199914
rect 175932 199884 175980 199914
rect 176423 199914 176532 199916
rect 175932 199858 175964 199884
rect 175871 199853 175964 199858
rect 175920 199822 175964 199853
rect 175958 199820 175964 199822
rect 176028 199820 176034 199884
rect 176423 199858 176428 199914
rect 176484 199884 176532 199914
rect 176484 199858 176516 199884
rect 176423 199853 176516 199858
rect 176472 199822 176516 199853
rect 176510 199820 176516 199822
rect 176580 199820 176586 199884
rect 177067 199882 177133 199885
rect 178217 199882 178283 199885
rect 177067 199880 178283 199882
rect 177067 199824 177072 199880
rect 177128 199824 178222 199880
rect 178278 199824 178283 199880
rect 177067 199822 178283 199824
rect 177067 199819 177133 199822
rect 178217 199819 178283 199822
rect 173566 199746 173572 199748
rect 173206 199686 173572 199746
rect 173566 199684 173572 199686
rect 173636 199684 173642 199748
rect 174264 199686 174308 199748
rect 174302 199684 174308 199686
rect 174372 199684 174378 199748
rect 174537 199746 174603 199749
rect 179045 199746 179111 199749
rect 174537 199744 179111 199746
rect 174537 199688 174542 199744
rect 174598 199688 179050 199744
rect 179106 199688 179111 199744
rect 174537 199686 179111 199688
rect 174537 199683 174603 199686
rect 179045 199683 179111 199686
rect 170673 199610 170739 199613
rect 177941 199610 178007 199613
rect 170673 199608 178007 199610
rect 170673 199552 170678 199608
rect 170734 199552 177946 199608
rect 178002 199552 178007 199608
rect 170673 199550 178007 199552
rect 170673 199547 170739 199550
rect 177941 199547 178007 199550
rect 170949 199474 171015 199477
rect 170262 199472 171015 199474
rect 170262 199416 170954 199472
rect 171010 199416 171015 199472
rect 170262 199414 171015 199416
rect 169772 199412 169778 199414
rect 169937 199411 170003 199414
rect 170949 199411 171015 199414
rect 171726 199412 171732 199476
rect 171796 199474 171802 199476
rect 171796 199414 179430 199474
rect 171796 199412 171802 199414
rect 168966 199338 168972 199340
rect 168790 199278 168972 199338
rect 166073 199275 166139 199278
rect 168649 199275 168715 199278
rect 168966 199276 168972 199278
rect 169036 199276 169042 199340
rect 169201 199338 169267 199341
rect 174261 199338 174327 199341
rect 169201 199336 174327 199338
rect 169201 199280 169206 199336
rect 169262 199280 174266 199336
rect 174322 199280 174327 199336
rect 169201 199278 174327 199280
rect 169201 199275 169267 199278
rect 174261 199275 174327 199278
rect 174629 199338 174695 199341
rect 174854 199338 174860 199340
rect 174629 199336 174860 199338
rect 174629 199280 174634 199336
rect 174690 199280 174860 199336
rect 174629 199278 174860 199280
rect 174629 199275 174695 199278
rect 174854 199276 174860 199278
rect 174924 199276 174930 199340
rect 179370 199338 179430 199414
rect 204621 199338 204687 199341
rect 179370 199336 204687 199338
rect 179370 199280 204626 199336
rect 204682 199280 204687 199336
rect 179370 199278 204687 199280
rect 204621 199275 204687 199278
rect 164325 199202 164391 199205
rect 175917 199202 175983 199205
rect 200798 199202 200804 199204
rect 164325 199200 175983 199202
rect 164325 199144 164330 199200
rect 164386 199144 175922 199200
rect 175978 199144 175983 199200
rect 164325 199142 175983 199144
rect 164325 199139 164391 199142
rect 175917 199139 175983 199142
rect 176702 199142 200804 199202
rect 164601 199066 164667 199069
rect 169753 199066 169819 199069
rect 164601 199064 169819 199066
rect 164601 199008 164606 199064
rect 164662 199008 169758 199064
rect 169814 199008 169819 199064
rect 164601 199006 169819 199008
rect 164601 199003 164667 199006
rect 169753 199003 169819 199006
rect 174169 199066 174235 199069
rect 176702 199066 176762 199142
rect 200798 199140 200804 199142
rect 200868 199140 200874 199204
rect 174169 199064 176762 199066
rect 174169 199008 174174 199064
rect 174230 199008 176762 199064
rect 174169 199006 176762 199008
rect 179045 199066 179111 199069
rect 200614 199066 200620 199068
rect 179045 199064 200620 199066
rect 179045 199008 179050 199064
rect 179106 199008 200620 199064
rect 179045 199006 200620 199008
rect 174169 199003 174235 199006
rect 179045 199003 179111 199006
rect 200614 199004 200620 199006
rect 200684 199004 200690 199068
rect 157149 198928 163882 198930
rect 157149 198872 157154 198928
rect 157210 198872 163882 198928
rect 157149 198870 163882 198872
rect 166257 198930 166323 198933
rect 173065 198930 173131 198933
rect 174169 198932 174235 198933
rect 166257 198928 173131 198930
rect 166257 198872 166262 198928
rect 166318 198872 173070 198928
rect 173126 198872 173131 198928
rect 166257 198870 173131 198872
rect 157149 198867 157215 198870
rect 166257 198867 166323 198870
rect 173065 198867 173131 198870
rect 174118 198868 174124 198932
rect 174188 198930 174235 198932
rect 174188 198928 174280 198930
rect 174230 198872 174280 198928
rect 174188 198870 174280 198872
rect 174188 198868 174235 198870
rect 174486 198868 174492 198932
rect 174556 198930 174562 198932
rect 200982 198930 200988 198932
rect 174556 198870 200988 198930
rect 174556 198868 174562 198870
rect 200982 198868 200988 198870
rect 201052 198868 201058 198932
rect 174169 198867 174235 198868
rect 163262 198794 163268 198796
rect 143092 198792 143184 198794
rect 143134 198736 143184 198792
rect 143092 198734 143184 198736
rect 156278 198734 163268 198794
rect 143092 198732 143139 198734
rect 163262 198732 163268 198734
rect 163332 198732 163338 198796
rect 166901 198794 166967 198797
rect 172237 198794 172303 198797
rect 166901 198792 172303 198794
rect 166901 198736 166906 198792
rect 166962 198736 172242 198792
rect 172298 198736 172303 198792
rect 166901 198734 172303 198736
rect 143073 198731 143139 198732
rect 166901 198731 166967 198734
rect 172237 198731 172303 198734
rect 176009 198794 176075 198797
rect 189022 198794 189028 198796
rect 176009 198792 189028 198794
rect 176009 198736 176014 198792
rect 176070 198736 189028 198792
rect 176009 198734 189028 198736
rect 176009 198731 176075 198734
rect 189022 198732 189028 198734
rect 189092 198732 189098 198796
rect 133505 198658 133571 198661
rect 133638 198658 133644 198660
rect 133505 198656 133644 198658
rect 133505 198600 133510 198656
rect 133566 198600 133644 198656
rect 133505 198598 133644 198600
rect 133505 198595 133571 198598
rect 133638 198596 133644 198598
rect 133708 198596 133714 198660
rect 134374 198596 134380 198660
rect 134444 198658 134450 198660
rect 134517 198658 134583 198661
rect 134444 198656 134583 198658
rect 134444 198600 134522 198656
rect 134578 198600 134583 198656
rect 134444 198598 134583 198600
rect 134444 198596 134450 198598
rect 134517 198595 134583 198598
rect 169150 198596 169156 198660
rect 169220 198658 169226 198660
rect 170857 198658 170923 198661
rect 169220 198656 170923 198658
rect 169220 198600 170862 198656
rect 170918 198600 170923 198656
rect 169220 198598 170923 198600
rect 169220 198596 169226 198598
rect 170857 198595 170923 198598
rect 171542 198596 171548 198660
rect 171612 198658 171618 198660
rect 187918 198658 187924 198660
rect 171612 198598 187924 198658
rect 171612 198596 171618 198598
rect 187918 198596 187924 198598
rect 187988 198596 187994 198660
rect 138105 198522 138171 198525
rect 138422 198522 138428 198524
rect 138105 198520 138428 198522
rect 138105 198464 138110 198520
rect 138166 198464 138428 198520
rect 138105 198462 138428 198464
rect 138105 198459 138171 198462
rect 138422 198460 138428 198462
rect 138492 198460 138498 198524
rect 155166 198460 155172 198524
rect 155236 198522 155242 198524
rect 159541 198522 159607 198525
rect 155236 198520 159607 198522
rect 155236 198464 159546 198520
rect 159602 198464 159607 198520
rect 155236 198462 159607 198464
rect 155236 198460 155242 198462
rect 159541 198459 159607 198462
rect 175365 198522 175431 198525
rect 175590 198522 175596 198524
rect 175365 198520 175596 198522
rect 175365 198464 175370 198520
rect 175426 198464 175596 198520
rect 175365 198462 175596 198464
rect 175365 198459 175431 198462
rect 175590 198460 175596 198462
rect 175660 198460 175666 198524
rect 107510 198324 107516 198388
rect 107580 198386 107586 198388
rect 132493 198386 132559 198389
rect 107580 198384 132559 198386
rect 107580 198328 132498 198384
rect 132554 198328 132559 198384
rect 107580 198326 132559 198328
rect 107580 198324 107586 198326
rect 132493 198323 132559 198326
rect 161238 198324 161244 198388
rect 161308 198386 161314 198388
rect 168373 198386 168439 198389
rect 161308 198384 168439 198386
rect 161308 198328 168378 198384
rect 168434 198328 168439 198384
rect 161308 198326 168439 198328
rect 161308 198324 161314 198326
rect 168373 198323 168439 198326
rect 168598 198324 168604 198388
rect 168668 198386 168674 198388
rect 171225 198386 171291 198389
rect 168668 198384 171291 198386
rect 168668 198328 171230 198384
rect 171286 198328 171291 198384
rect 168668 198326 171291 198328
rect 168668 198324 168674 198326
rect 171225 198323 171291 198326
rect 173249 198386 173315 198389
rect 201166 198386 201172 198388
rect 173249 198384 201172 198386
rect 173249 198328 173254 198384
rect 173310 198328 201172 198384
rect 173249 198326 201172 198328
rect 173249 198323 173315 198326
rect 201166 198324 201172 198326
rect 201236 198324 201242 198388
rect 105905 198250 105971 198253
rect 132401 198250 132467 198253
rect 105905 198248 132467 198250
rect 105905 198192 105910 198248
rect 105966 198192 132406 198248
rect 132462 198192 132467 198248
rect 105905 198190 132467 198192
rect 105905 198187 105971 198190
rect 132401 198187 132467 198190
rect 140865 198250 140931 198253
rect 143574 198250 143580 198252
rect 140865 198248 143580 198250
rect 140865 198192 140870 198248
rect 140926 198192 143580 198248
rect 140865 198190 143580 198192
rect 140865 198187 140931 198190
rect 143574 198188 143580 198190
rect 143644 198188 143650 198252
rect 148910 198188 148916 198252
rect 148980 198250 148986 198252
rect 158621 198250 158687 198253
rect 148980 198248 158687 198250
rect 148980 198192 158626 198248
rect 158682 198192 158687 198248
rect 148980 198190 158687 198192
rect 148980 198188 148986 198190
rect 158621 198187 158687 198190
rect 170581 198250 170647 198253
rect 209865 198250 209931 198253
rect 170581 198248 209931 198250
rect 170581 198192 170586 198248
rect 170642 198192 209870 198248
rect 209926 198192 209931 198248
rect 170581 198190 209931 198192
rect 170581 198187 170647 198190
rect 209865 198187 209931 198190
rect 106958 198052 106964 198116
rect 107028 198114 107034 198116
rect 133229 198114 133295 198117
rect 140957 198116 141023 198117
rect 140957 198114 141004 198116
rect 107028 198112 133295 198114
rect 107028 198056 133234 198112
rect 133290 198056 133295 198112
rect 107028 198054 133295 198056
rect 140912 198112 141004 198114
rect 140912 198056 140962 198112
rect 140912 198054 141004 198056
rect 107028 198052 107034 198054
rect 133229 198051 133295 198054
rect 140957 198052 141004 198054
rect 141068 198052 141074 198116
rect 147857 198114 147923 198117
rect 153469 198116 153535 198117
rect 148174 198114 148180 198116
rect 147857 198112 148180 198114
rect 147857 198056 147862 198112
rect 147918 198056 148180 198112
rect 147857 198054 148180 198056
rect 140957 198051 141023 198052
rect 147857 198051 147923 198054
rect 148174 198052 148180 198054
rect 148244 198052 148250 198116
rect 153469 198114 153516 198116
rect 153424 198112 153516 198114
rect 153424 198056 153474 198112
rect 153424 198054 153516 198056
rect 153469 198052 153516 198054
rect 153580 198052 153586 198116
rect 171041 198114 171107 198117
rect 212809 198114 212875 198117
rect 171041 198112 212875 198114
rect 171041 198056 171046 198112
rect 171102 198056 212814 198112
rect 212870 198056 212875 198112
rect 171041 198054 212875 198056
rect 153469 198051 153535 198052
rect 171041 198051 171107 198054
rect 212809 198051 212875 198054
rect 102910 197916 102916 197980
rect 102980 197978 102986 197980
rect 132033 197978 132099 197981
rect 102980 197976 132099 197978
rect 102980 197920 132038 197976
rect 132094 197920 132099 197976
rect 102980 197918 132099 197920
rect 102980 197916 102986 197918
rect 132033 197915 132099 197918
rect 153142 197916 153148 197980
rect 153212 197978 153218 197980
rect 153561 197978 153627 197981
rect 153212 197976 153627 197978
rect 153212 197920 153566 197976
rect 153622 197920 153627 197976
rect 153212 197918 153627 197920
rect 153212 197916 153218 197918
rect 153561 197915 153627 197918
rect 154430 197916 154436 197980
rect 154500 197978 154506 197980
rect 165286 197978 165292 197980
rect 154500 197918 165292 197978
rect 154500 197916 154506 197918
rect 165286 197916 165292 197918
rect 165356 197916 165362 197980
rect 172145 197978 172211 197981
rect 172278 197978 172284 197980
rect 172145 197976 172284 197978
rect 172145 197920 172150 197976
rect 172206 197920 172284 197976
rect 172145 197918 172284 197920
rect 172145 197915 172211 197918
rect 172278 197916 172284 197918
rect 172348 197916 172354 197980
rect 172605 197978 172671 197981
rect 212993 197978 213059 197981
rect 172605 197976 213059 197978
rect 172605 197920 172610 197976
rect 172666 197920 212998 197976
rect 213054 197920 213059 197976
rect 172605 197918 213059 197920
rect 172605 197915 172671 197918
rect 212993 197915 213059 197918
rect 157742 197780 157748 197844
rect 157812 197842 157818 197844
rect 162485 197842 162551 197845
rect 157812 197840 162551 197842
rect 157812 197784 162490 197840
rect 162546 197784 162551 197840
rect 157812 197782 162551 197784
rect 157812 197780 157818 197782
rect 162485 197779 162551 197782
rect 171593 197842 171659 197845
rect 186998 197842 187004 197844
rect 171593 197840 187004 197842
rect 171593 197784 171598 197840
rect 171654 197784 187004 197840
rect 171593 197782 187004 197784
rect 171593 197779 171659 197782
rect 186998 197780 187004 197782
rect 187068 197780 187074 197844
rect 175181 197706 175247 197709
rect 176326 197706 176332 197708
rect 175181 197704 176332 197706
rect 175181 197648 175186 197704
rect 175242 197648 176332 197704
rect 175181 197646 176332 197648
rect 175181 197643 175247 197646
rect 176326 197644 176332 197646
rect 176396 197644 176402 197708
rect 164325 197570 164391 197573
rect 164918 197570 164924 197572
rect 164325 197568 164924 197570
rect 164325 197512 164330 197568
rect 164386 197512 164924 197568
rect 164325 197510 164924 197512
rect 164325 197507 164391 197510
rect 164918 197508 164924 197510
rect 164988 197508 164994 197572
rect 171317 197570 171383 197573
rect 188102 197570 188108 197572
rect 171317 197568 188108 197570
rect 171317 197512 171322 197568
rect 171378 197512 188108 197568
rect 171317 197510 188108 197512
rect 171317 197507 171383 197510
rect 188102 197508 188108 197510
rect 188172 197508 188178 197572
rect 164734 197372 164740 197436
rect 164804 197434 164810 197436
rect 171777 197434 171843 197437
rect 164804 197432 171843 197434
rect 164804 197376 171782 197432
rect 171838 197376 171843 197432
rect 164804 197374 171843 197376
rect 164804 197372 164810 197374
rect 171777 197371 171843 197374
rect 172789 197434 172855 197437
rect 173750 197434 173756 197436
rect 172789 197432 173756 197434
rect 172789 197376 172794 197432
rect 172850 197376 173756 197432
rect 172789 197374 173756 197376
rect 172789 197371 172855 197374
rect 173750 197372 173756 197374
rect 173820 197372 173826 197436
rect 175457 197434 175523 197437
rect 175958 197434 175964 197436
rect 175457 197432 175964 197434
rect 175457 197376 175462 197432
rect 175518 197376 175964 197432
rect 175457 197374 175964 197376
rect 175457 197371 175523 197374
rect 175958 197372 175964 197374
rect 176028 197372 176034 197436
rect 136582 197236 136588 197300
rect 136652 197298 136658 197300
rect 137277 197298 137343 197301
rect 139761 197300 139827 197301
rect 139710 197298 139716 197300
rect 136652 197296 137343 197298
rect 136652 197240 137282 197296
rect 137338 197240 137343 197296
rect 136652 197238 137343 197240
rect 139670 197238 139716 197298
rect 139780 197296 139827 197300
rect 139822 197240 139827 197296
rect 136652 197236 136658 197238
rect 137277 197235 137343 197238
rect 139710 197236 139716 197238
rect 139780 197236 139827 197240
rect 139761 197235 139827 197236
rect 160645 197298 160711 197301
rect 162342 197298 162348 197300
rect 160645 197296 162348 197298
rect 160645 197240 160650 197296
rect 160706 197240 162348 197296
rect 160645 197238 162348 197240
rect 160645 197235 160711 197238
rect 162342 197236 162348 197238
rect 162412 197236 162418 197300
rect 165153 197298 165219 197301
rect 198825 197298 198891 197301
rect 165153 197296 198891 197298
rect 165153 197240 165158 197296
rect 165214 197240 198830 197296
rect 198886 197240 198891 197296
rect 165153 197238 198891 197240
rect 165153 197235 165219 197238
rect 198825 197235 198891 197238
rect 136725 197162 136791 197165
rect 136950 197162 136956 197164
rect 136725 197160 136956 197162
rect 136725 197104 136730 197160
rect 136786 197104 136956 197160
rect 136725 197102 136956 197104
rect 136725 197099 136791 197102
rect 136950 197100 136956 197102
rect 137020 197100 137026 197164
rect 164233 197162 164299 197165
rect 197445 197162 197511 197165
rect 164233 197160 197511 197162
rect 164233 197104 164238 197160
rect 164294 197104 197450 197160
rect 197506 197104 197511 197160
rect 164233 197102 197511 197104
rect 164233 197099 164299 197102
rect 197445 197099 197511 197102
rect 131757 197026 131823 197029
rect 152457 197026 152523 197029
rect 131757 197024 152523 197026
rect 131757 196968 131762 197024
rect 131818 196968 152462 197024
rect 152518 196968 152523 197024
rect 131757 196966 152523 196968
rect 131757 196963 131823 196966
rect 152457 196963 152523 196966
rect 166625 197026 166691 197029
rect 200205 197026 200271 197029
rect 166625 197024 200271 197026
rect 166625 196968 166630 197024
rect 166686 196968 200210 197024
rect 200266 196968 200271 197024
rect 166625 196966 200271 196968
rect 166625 196963 166691 196966
rect 200205 196963 200271 196966
rect 106917 196890 106983 196893
rect 136541 196890 136607 196893
rect 136817 196892 136883 196893
rect 136766 196890 136772 196892
rect 106917 196888 136607 196890
rect 106917 196832 106922 196888
rect 106978 196832 136546 196888
rect 136602 196832 136607 196888
rect 106917 196830 136607 196832
rect 136726 196830 136772 196890
rect 136836 196888 136883 196892
rect 137461 196892 137527 196893
rect 137461 196890 137508 196892
rect 136878 196832 136883 196888
rect 106917 196827 106983 196830
rect 136541 196827 136607 196830
rect 136766 196828 136772 196830
rect 136836 196828 136883 196832
rect 137416 196888 137508 196890
rect 137416 196832 137466 196888
rect 137416 196830 137508 196832
rect 136817 196827 136883 196828
rect 137461 196828 137508 196830
rect 137572 196828 137578 196892
rect 138054 196828 138060 196892
rect 138124 196890 138130 196892
rect 138657 196890 138723 196893
rect 138124 196888 138723 196890
rect 138124 196832 138662 196888
rect 138718 196832 138723 196888
rect 138124 196830 138723 196832
rect 138124 196828 138130 196830
rect 137461 196827 137527 196828
rect 138657 196827 138723 196830
rect 142470 196828 142476 196892
rect 142540 196890 142546 196892
rect 143165 196890 143231 196893
rect 142540 196888 143231 196890
rect 142540 196832 143170 196888
rect 143226 196832 143231 196888
rect 142540 196830 143231 196832
rect 142540 196828 142546 196830
rect 143165 196827 143231 196830
rect 145097 196890 145163 196893
rect 146702 196890 146708 196892
rect 145097 196888 146708 196890
rect 145097 196832 145102 196888
rect 145158 196832 146708 196888
rect 145097 196830 146708 196832
rect 145097 196827 145163 196830
rect 146702 196828 146708 196830
rect 146772 196828 146778 196892
rect 147070 196828 147076 196892
rect 147140 196890 147146 196892
rect 151169 196890 151235 196893
rect 153193 196890 153259 196893
rect 157149 196892 157215 196893
rect 157149 196890 157196 196892
rect 147140 196888 151235 196890
rect 147140 196832 151174 196888
rect 151230 196832 151235 196888
rect 147140 196830 151235 196832
rect 147140 196828 147146 196830
rect 151169 196827 151235 196830
rect 151494 196888 153259 196890
rect 151494 196832 153198 196888
rect 153254 196832 153259 196888
rect 151494 196830 153259 196832
rect 157104 196888 157196 196890
rect 157104 196832 157154 196888
rect 157104 196830 157196 196832
rect 121177 196754 121243 196757
rect 151494 196754 151554 196830
rect 153193 196827 153259 196830
rect 157149 196828 157196 196830
rect 157260 196828 157266 196892
rect 162393 196890 162459 196893
rect 162526 196890 162532 196892
rect 162393 196888 162532 196890
rect 162393 196832 162398 196888
rect 162454 196832 162532 196888
rect 162393 196830 162532 196832
rect 157149 196827 157215 196828
rect 162393 196827 162459 196830
rect 162526 196828 162532 196830
rect 162596 196828 162602 196892
rect 163446 196828 163452 196892
rect 163516 196890 163522 196892
rect 163589 196890 163655 196893
rect 163516 196888 163655 196890
rect 163516 196832 163594 196888
rect 163650 196832 163655 196888
rect 163516 196830 163655 196832
rect 163516 196828 163522 196830
rect 163589 196827 163655 196830
rect 164141 196890 164207 196893
rect 197302 196890 197308 196892
rect 164141 196888 197308 196890
rect 164141 196832 164146 196888
rect 164202 196832 197308 196888
rect 164141 196830 197308 196832
rect 164141 196827 164207 196830
rect 197302 196828 197308 196830
rect 197372 196828 197378 196892
rect 121177 196752 151554 196754
rect 121177 196696 121182 196752
rect 121238 196696 151554 196752
rect 121177 196694 151554 196696
rect 121177 196691 121243 196694
rect 157190 196692 157196 196756
rect 157260 196754 157266 196756
rect 161105 196754 161171 196757
rect 157260 196752 161171 196754
rect 157260 196696 161110 196752
rect 161166 196696 161171 196752
rect 157260 196694 161171 196696
rect 157260 196692 157266 196694
rect 161105 196691 161171 196694
rect 162209 196754 162275 196757
rect 196249 196754 196315 196757
rect 162209 196752 196315 196754
rect 162209 196696 162214 196752
rect 162270 196696 196254 196752
rect 196310 196696 196315 196752
rect 162209 196694 196315 196696
rect 162209 196691 162275 196694
rect 196249 196691 196315 196694
rect 113030 196556 113036 196620
rect 113100 196618 113106 196620
rect 147397 196618 147463 196621
rect 113100 196616 147463 196618
rect 113100 196560 147402 196616
rect 147458 196560 147463 196616
rect 113100 196558 147463 196560
rect 113100 196556 113106 196558
rect 147397 196555 147463 196558
rect 148174 196556 148180 196620
rect 148244 196618 148250 196620
rect 151445 196618 151511 196621
rect 148244 196616 151511 196618
rect 148244 196560 151450 196616
rect 151506 196560 151511 196616
rect 148244 196558 151511 196560
rect 148244 196556 148250 196558
rect 151445 196555 151511 196558
rect 157333 196618 157399 196621
rect 157558 196618 157564 196620
rect 157333 196616 157564 196618
rect 157333 196560 157338 196616
rect 157394 196560 157564 196616
rect 157333 196558 157564 196560
rect 157333 196555 157399 196558
rect 157558 196556 157564 196558
rect 157628 196556 157634 196620
rect 157885 196618 157951 196621
rect 192753 196618 192819 196621
rect 157885 196616 192819 196618
rect 157885 196560 157890 196616
rect 157946 196560 192758 196616
rect 192814 196560 192819 196616
rect 157885 196558 192819 196560
rect 157885 196555 157951 196558
rect 192753 196555 192819 196558
rect 142286 196420 142292 196484
rect 142356 196482 142362 196484
rect 143809 196482 143875 196485
rect 142356 196480 143875 196482
rect 142356 196424 143814 196480
rect 143870 196424 143875 196480
rect 142356 196422 143875 196424
rect 142356 196420 142362 196422
rect 143809 196419 143875 196422
rect 161054 196420 161060 196484
rect 161124 196482 161130 196484
rect 161197 196482 161263 196485
rect 161124 196480 161263 196482
rect 161124 196424 161202 196480
rect 161258 196424 161263 196480
rect 161124 196422 161263 196424
rect 161124 196420 161130 196422
rect 161197 196419 161263 196422
rect 163078 196420 163084 196484
rect 163148 196482 163154 196484
rect 163313 196482 163379 196485
rect 164969 196484 165035 196485
rect 164918 196482 164924 196484
rect 163148 196480 163379 196482
rect 163148 196424 163318 196480
rect 163374 196424 163379 196480
rect 163148 196422 163379 196424
rect 164878 196422 164924 196482
rect 164988 196480 165035 196484
rect 165030 196424 165035 196480
rect 163148 196420 163154 196422
rect 163313 196419 163379 196422
rect 164918 196420 164924 196422
rect 164988 196420 165035 196424
rect 167678 196420 167684 196484
rect 167748 196482 167754 196484
rect 168281 196482 168347 196485
rect 167748 196480 168347 196482
rect 167748 196424 168286 196480
rect 168342 196424 168347 196480
rect 167748 196422 168347 196424
rect 167748 196420 167754 196422
rect 164969 196419 165035 196420
rect 168281 196419 168347 196422
rect 169109 196484 169175 196485
rect 169109 196480 169156 196484
rect 169220 196482 169226 196484
rect 169569 196482 169635 196485
rect 171317 196484 171383 196485
rect 170806 196482 170812 196484
rect 169109 196424 169114 196480
rect 169109 196420 169156 196424
rect 169220 196422 169266 196482
rect 169569 196480 170812 196482
rect 169569 196424 169574 196480
rect 169630 196424 170812 196480
rect 169569 196422 170812 196424
rect 169220 196420 169226 196422
rect 169109 196419 169175 196420
rect 169569 196419 169635 196422
rect 170806 196420 170812 196422
rect 170876 196420 170882 196484
rect 171317 196482 171364 196484
rect 171272 196480 171364 196482
rect 171272 196424 171322 196480
rect 171272 196422 171364 196424
rect 171317 196420 171364 196422
rect 171428 196420 171434 196484
rect 172053 196482 172119 196485
rect 193254 196482 193260 196484
rect 172053 196480 193260 196482
rect 172053 196424 172058 196480
rect 172114 196424 193260 196480
rect 172053 196422 193260 196424
rect 171317 196419 171383 196420
rect 172053 196419 172119 196422
rect 193254 196420 193260 196422
rect 193324 196420 193330 196484
rect 133781 196346 133847 196349
rect 134006 196346 134012 196348
rect 133781 196344 134012 196346
rect 133781 196288 133786 196344
rect 133842 196288 134012 196344
rect 133781 196286 134012 196288
rect 133781 196283 133847 196286
rect 134006 196284 134012 196286
rect 134076 196284 134082 196348
rect 163405 196346 163471 196349
rect 166073 196348 166139 196349
rect 163814 196346 163820 196348
rect 163405 196344 163820 196346
rect 163405 196288 163410 196344
rect 163466 196288 163820 196344
rect 163405 196286 163820 196288
rect 163405 196283 163471 196286
rect 163814 196284 163820 196286
rect 163884 196284 163890 196348
rect 166022 196284 166028 196348
rect 166092 196346 166139 196348
rect 166092 196344 166184 196346
rect 166134 196288 166184 196344
rect 166092 196286 166184 196288
rect 166092 196284 166139 196286
rect 168782 196284 168788 196348
rect 168852 196346 168858 196348
rect 169017 196346 169083 196349
rect 168852 196344 169083 196346
rect 168852 196288 169022 196344
rect 169078 196288 169083 196344
rect 168852 196286 169083 196288
rect 168852 196284 168858 196286
rect 166073 196283 166139 196284
rect 169017 196283 169083 196286
rect 169845 196346 169911 196349
rect 172513 196348 172579 196349
rect 170070 196346 170076 196348
rect 169845 196344 170076 196346
rect 169845 196288 169850 196344
rect 169906 196288 170076 196344
rect 169845 196286 170076 196288
rect 169845 196283 169911 196286
rect 170070 196284 170076 196286
rect 170140 196284 170146 196348
rect 172462 196284 172468 196348
rect 172532 196346 172579 196348
rect 172697 196346 172763 196349
rect 173382 196346 173388 196348
rect 172532 196344 172624 196346
rect 172574 196288 172624 196344
rect 172532 196286 172624 196288
rect 172697 196344 173388 196346
rect 172697 196288 172702 196344
rect 172758 196288 173388 196344
rect 172697 196286 173388 196288
rect 172532 196284 172579 196286
rect 172513 196283 172579 196284
rect 172697 196283 172763 196286
rect 173382 196284 173388 196286
rect 173452 196284 173458 196348
rect 135253 196212 135319 196213
rect 135253 196210 135300 196212
rect 135208 196208 135300 196210
rect 135208 196152 135258 196208
rect 135208 196150 135300 196152
rect 135253 196148 135300 196150
rect 135364 196148 135370 196212
rect 167494 196148 167500 196212
rect 167564 196210 167570 196212
rect 167637 196210 167703 196213
rect 167564 196208 167703 196210
rect 167564 196152 167642 196208
rect 167698 196152 167703 196208
rect 167564 196150 167703 196152
rect 167564 196148 167570 196150
rect 135253 196147 135319 196148
rect 167637 196147 167703 196150
rect 169518 196148 169524 196212
rect 169588 196210 169594 196212
rect 169753 196210 169819 196213
rect 169588 196208 169819 196210
rect 169588 196152 169758 196208
rect 169814 196152 169819 196208
rect 169588 196150 169819 196152
rect 169588 196148 169594 196150
rect 169753 196147 169819 196150
rect 170121 196210 170187 196213
rect 170622 196210 170628 196212
rect 170121 196208 170628 196210
rect 170121 196152 170126 196208
rect 170182 196152 170628 196208
rect 170121 196150 170628 196152
rect 170121 196147 170187 196150
rect 170622 196148 170628 196150
rect 170692 196148 170698 196212
rect 171910 196148 171916 196212
rect 171980 196210 171986 196212
rect 173157 196210 173223 196213
rect 171980 196208 173223 196210
rect 171980 196152 173162 196208
rect 173218 196152 173223 196208
rect 171980 196150 173223 196152
rect 171980 196148 171986 196150
rect 173157 196147 173223 196150
rect 135294 196012 135300 196076
rect 135364 196074 135370 196076
rect 135529 196074 135595 196077
rect 135364 196072 135595 196074
rect 135364 196016 135534 196072
rect 135590 196016 135595 196072
rect 135364 196014 135595 196016
rect 135364 196012 135370 196014
rect 135529 196011 135595 196014
rect 158110 196012 158116 196076
rect 158180 196074 158186 196076
rect 158529 196074 158595 196077
rect 158180 196072 158595 196074
rect 158180 196016 158534 196072
rect 158590 196016 158595 196072
rect 158180 196014 158595 196016
rect 158180 196012 158186 196014
rect 158529 196011 158595 196014
rect 161422 196012 161428 196076
rect 161492 196074 161498 196076
rect 161749 196074 161815 196077
rect 161492 196072 161815 196074
rect 161492 196016 161754 196072
rect 161810 196016 161815 196072
rect 161492 196014 161815 196016
rect 161492 196012 161498 196014
rect 161749 196011 161815 196014
rect 165838 196012 165844 196076
rect 165908 196074 165914 196076
rect 169385 196074 169451 196077
rect 165908 196072 169451 196074
rect 165908 196016 169390 196072
rect 169446 196016 169451 196072
rect 165908 196014 169451 196016
rect 165908 196012 165914 196014
rect 169385 196011 169451 196014
rect 169886 196012 169892 196076
rect 169956 196074 169962 196076
rect 171593 196074 171659 196077
rect 169956 196072 171659 196074
rect 169956 196016 171598 196072
rect 171654 196016 171659 196072
rect 169956 196014 171659 196016
rect 169956 196012 169962 196014
rect 171593 196011 171659 196014
rect 135345 195938 135411 195941
rect 135662 195938 135668 195940
rect 135345 195936 135668 195938
rect 135345 195880 135350 195936
rect 135406 195880 135668 195936
rect 135345 195878 135668 195880
rect 135345 195875 135411 195878
rect 135662 195876 135668 195878
rect 135732 195876 135738 195940
rect 142429 195938 142495 195941
rect 142838 195938 142844 195940
rect 142429 195936 142844 195938
rect 142429 195880 142434 195936
rect 142490 195880 142844 195936
rect 142429 195878 142844 195880
rect 142429 195875 142495 195878
rect 142838 195876 142844 195878
rect 142908 195876 142914 195940
rect 153745 195938 153811 195941
rect 184054 195938 184060 195940
rect 153745 195936 184060 195938
rect 153745 195880 153750 195936
rect 153806 195880 184060 195936
rect 153745 195878 184060 195880
rect 153745 195875 153811 195878
rect 184054 195876 184060 195878
rect 184124 195876 184130 195940
rect 119981 195802 120047 195805
rect 130326 195802 130332 195804
rect 119981 195800 130332 195802
rect 119981 195744 119986 195800
rect 120042 195744 130332 195800
rect 119981 195742 130332 195744
rect 119981 195739 120047 195742
rect 130326 195740 130332 195742
rect 130396 195740 130402 195804
rect 139526 195740 139532 195804
rect 139596 195802 139602 195804
rect 140221 195802 140287 195805
rect 139596 195800 140287 195802
rect 139596 195744 140226 195800
rect 140282 195744 140287 195800
rect 139596 195742 140287 195744
rect 139596 195740 139602 195742
rect 140221 195739 140287 195742
rect 161565 195802 161631 195805
rect 161790 195802 161796 195804
rect 161565 195800 161796 195802
rect 161565 195744 161570 195800
rect 161626 195744 161796 195800
rect 161565 195742 161796 195744
rect 161565 195739 161631 195742
rect 161790 195740 161796 195742
rect 161860 195740 161866 195804
rect 166257 195802 166323 195805
rect 166574 195802 166580 195804
rect 166257 195800 166580 195802
rect 166257 195744 166262 195800
rect 166318 195744 166580 195800
rect 166257 195742 166580 195744
rect 166257 195739 166323 195742
rect 166574 195740 166580 195742
rect 166644 195740 166650 195804
rect 167913 195802 167979 195805
rect 196065 195802 196131 195805
rect 167913 195800 196131 195802
rect 167913 195744 167918 195800
rect 167974 195744 196070 195800
rect 196126 195744 196131 195800
rect 167913 195742 196131 195744
rect 167913 195739 167979 195742
rect 196065 195739 196131 195742
rect 104014 195604 104020 195668
rect 104084 195666 104090 195668
rect 135437 195666 135503 195669
rect 104084 195664 135503 195666
rect 104084 195608 135442 195664
rect 135498 195608 135503 195664
rect 104084 195606 135503 195608
rect 104084 195604 104090 195606
rect 135437 195603 135503 195606
rect 146886 195604 146892 195668
rect 146956 195666 146962 195668
rect 149697 195666 149763 195669
rect 146956 195664 149763 195666
rect 146956 195608 149702 195664
rect 149758 195608 149763 195664
rect 146956 195606 149763 195608
rect 146956 195604 146962 195606
rect 149697 195603 149763 195606
rect 153878 195604 153884 195668
rect 153948 195666 153954 195668
rect 154297 195666 154363 195669
rect 153948 195664 154363 195666
rect 153948 195608 154302 195664
rect 154358 195608 154363 195664
rect 153948 195606 154363 195608
rect 153948 195604 153954 195606
rect 154297 195603 154363 195606
rect 162025 195666 162091 195669
rect 191925 195666 191991 195669
rect 162025 195664 191991 195666
rect 162025 195608 162030 195664
rect 162086 195608 191930 195664
rect 191986 195608 191991 195664
rect 162025 195606 191991 195608
rect 162025 195603 162091 195606
rect 191925 195603 191991 195606
rect 108205 195530 108271 195533
rect 141877 195530 141943 195533
rect 108205 195528 141943 195530
rect 108205 195472 108210 195528
rect 108266 195472 141882 195528
rect 141938 195472 141943 195528
rect 108205 195470 141943 195472
rect 108205 195467 108271 195470
rect 141877 195467 141943 195470
rect 162577 195530 162643 195533
rect 196157 195530 196223 195533
rect 162577 195528 196223 195530
rect 162577 195472 162582 195528
rect 162638 195472 196162 195528
rect 196218 195472 196223 195528
rect 162577 195470 196223 195472
rect 162577 195467 162643 195470
rect 196157 195467 196223 195470
rect 100293 195394 100359 195397
rect 154205 195394 154271 195397
rect 100293 195392 154271 195394
rect 100293 195336 100298 195392
rect 100354 195336 154210 195392
rect 154266 195336 154271 195392
rect 100293 195334 154271 195336
rect 100293 195331 100359 195334
rect 154205 195331 154271 195334
rect 158805 195394 158871 195397
rect 160134 195394 160140 195396
rect 158805 195392 160140 195394
rect 158805 195336 158810 195392
rect 158866 195336 160140 195392
rect 158805 195334 160140 195336
rect 158805 195331 158871 195334
rect 160134 195332 160140 195334
rect 160204 195332 160210 195396
rect 161473 195394 161539 195397
rect 194542 195394 194548 195396
rect 161473 195392 194548 195394
rect 161473 195336 161478 195392
rect 161534 195336 194548 195392
rect 161473 195334 194548 195336
rect 161473 195331 161539 195334
rect 194542 195332 194548 195334
rect 194612 195332 194618 195396
rect 119838 195196 119844 195260
rect 119908 195258 119914 195260
rect 130561 195258 130627 195261
rect 119908 195256 130627 195258
rect 119908 195200 130566 195256
rect 130622 195200 130627 195256
rect 119908 195198 130627 195200
rect 119908 195196 119914 195198
rect 130561 195195 130627 195198
rect 168833 195258 168899 195261
rect 215385 195258 215451 195261
rect 168833 195256 215451 195258
rect 168833 195200 168838 195256
rect 168894 195200 215390 195256
rect 215446 195200 215451 195256
rect 168833 195198 215451 195200
rect 168833 195195 168899 195198
rect 215385 195195 215451 195198
rect 177665 195122 177731 195125
rect 199326 195122 199332 195124
rect 177665 195120 199332 195122
rect 177665 195064 177670 195120
rect 177726 195064 199332 195120
rect 177665 195062 199332 195064
rect 177665 195059 177731 195062
rect 199326 195060 199332 195062
rect 199396 195060 199402 195124
rect 175406 194788 175412 194852
rect 175476 194850 175482 194852
rect 183829 194850 183895 194853
rect 175476 194848 183895 194850
rect 175476 194792 183834 194848
rect 183890 194792 183895 194848
rect 175476 194790 183895 194792
rect 175476 194788 175482 194790
rect 183829 194787 183895 194790
rect 123569 194578 123635 194581
rect 148869 194578 148935 194581
rect 123569 194576 148935 194578
rect 123569 194520 123574 194576
rect 123630 194520 148874 194576
rect 148930 194520 148935 194576
rect 123569 194518 148935 194520
rect 123569 194515 123635 194518
rect 148869 194515 148935 194518
rect 167729 194578 167795 194581
rect 201718 194578 201724 194580
rect 167729 194576 201724 194578
rect 167729 194520 167734 194576
rect 167790 194520 201724 194576
rect 167729 194518 201724 194520
rect 167729 194515 167795 194518
rect 201718 194516 201724 194518
rect 201788 194516 201794 194580
rect 102726 194380 102732 194444
rect 102796 194442 102802 194444
rect 130101 194442 130167 194445
rect 102796 194440 130167 194442
rect 102796 194384 130106 194440
rect 130162 194384 130167 194440
rect 102796 194382 130167 194384
rect 102796 194380 102802 194382
rect 130101 194379 130167 194382
rect 144637 194442 144703 194445
rect 147254 194442 147260 194444
rect 144637 194440 147260 194442
rect 144637 194384 144642 194440
rect 144698 194384 147260 194440
rect 144637 194382 147260 194384
rect 144637 194379 144703 194382
rect 147254 194380 147260 194382
rect 147324 194380 147330 194444
rect 173014 194380 173020 194444
rect 173084 194442 173090 194444
rect 173433 194442 173499 194445
rect 173084 194440 173499 194442
rect 173084 194384 173438 194440
rect 173494 194384 173499 194440
rect 173084 194382 173499 194384
rect 173084 194380 173090 194382
rect 173433 194379 173499 194382
rect 174629 194442 174695 194445
rect 208577 194442 208643 194445
rect 174629 194440 208643 194442
rect 174629 194384 174634 194440
rect 174690 194384 208582 194440
rect 208638 194384 208643 194440
rect 174629 194382 208643 194384
rect 174629 194379 174695 194382
rect 208577 194379 208643 194382
rect 103237 194306 103303 194309
rect 134885 194306 134951 194309
rect 103237 194304 134951 194306
rect 103237 194248 103242 194304
rect 103298 194248 134890 194304
rect 134946 194248 134951 194304
rect 103237 194246 134951 194248
rect 103237 194243 103303 194246
rect 134885 194243 134951 194246
rect 142245 194308 142311 194309
rect 142245 194304 142292 194308
rect 142356 194306 142362 194308
rect 174537 194306 174603 194309
rect 208485 194306 208551 194309
rect 142245 194248 142250 194304
rect 142245 194244 142292 194248
rect 142356 194246 142402 194306
rect 174537 194304 208551 194306
rect 174537 194248 174542 194304
rect 174598 194248 208490 194304
rect 208546 194248 208551 194304
rect 174537 194246 208551 194248
rect 142356 194244 142362 194246
rect 142245 194243 142311 194244
rect 174537 194243 174603 194246
rect 208485 194243 208551 194246
rect 105997 194170 106063 194173
rect 138749 194170 138815 194173
rect 105997 194168 138815 194170
rect 105997 194112 106002 194168
rect 106058 194112 138754 194168
rect 138810 194112 138815 194168
rect 105997 194110 138815 194112
rect 105997 194107 106063 194110
rect 138749 194107 138815 194110
rect 172646 194108 172652 194172
rect 172716 194170 172722 194172
rect 207197 194170 207263 194173
rect 172716 194168 207263 194170
rect 172716 194112 207202 194168
rect 207258 194112 207263 194168
rect 172716 194110 207263 194112
rect 172716 194108 172722 194110
rect 207197 194107 207263 194110
rect 101673 194034 101739 194037
rect 134333 194034 134399 194037
rect 173617 194036 173683 194037
rect 101673 194032 134399 194034
rect 101673 193976 101678 194032
rect 101734 193976 134338 194032
rect 134394 193976 134399 194032
rect 101673 193974 134399 193976
rect 101673 193971 101739 193974
rect 134333 193971 134399 193974
rect 173566 193972 173572 194036
rect 173636 194034 173683 194036
rect 173636 194032 173728 194034
rect 173678 193976 173728 194032
rect 173636 193974 173728 193976
rect 173636 193972 173683 193974
rect 175590 193972 175596 194036
rect 175660 194034 175666 194036
rect 209998 194034 210004 194036
rect 175660 193974 210004 194034
rect 175660 193972 175666 193974
rect 209998 193972 210004 193974
rect 210068 193972 210074 194036
rect 173617 193971 173683 193972
rect 100334 193836 100340 193900
rect 100404 193898 100410 193900
rect 128353 193898 128419 193901
rect 100404 193896 128419 193898
rect 100404 193840 128358 193896
rect 128414 193840 128419 193896
rect 100404 193838 128419 193840
rect 100404 193836 100410 193838
rect 128353 193835 128419 193838
rect 182265 193898 182331 193901
rect 209814 193898 209820 193900
rect 182265 193896 209820 193898
rect 182265 193840 182270 193896
rect 182326 193840 209820 193896
rect 182265 193838 209820 193840
rect 182265 193835 182331 193838
rect 209814 193836 209820 193838
rect 209884 193836 209890 193900
rect 168741 193354 168807 193357
rect 168741 193352 175106 193354
rect 168741 193296 168746 193352
rect 168802 193296 175106 193352
rect 168741 193294 175106 193296
rect 168741 193291 168807 193294
rect 168005 193218 168071 193221
rect 175046 193218 175106 193294
rect 201902 193218 201908 193220
rect 168005 193216 174922 193218
rect 168005 193160 168010 193216
rect 168066 193160 174922 193216
rect 168005 193158 174922 193160
rect 175046 193158 201908 193218
rect 168005 193155 168071 193158
rect 169753 193082 169819 193085
rect 169753 193080 174738 193082
rect 169753 193024 169758 193080
rect 169814 193024 174738 193080
rect 169753 193022 174738 193024
rect 169753 193019 169819 193022
rect 174678 192810 174738 193022
rect 174862 192946 174922 193158
rect 201902 193156 201908 193158
rect 201972 193156 201978 193220
rect 175917 193082 175983 193085
rect 198774 193082 198780 193084
rect 175917 193080 198780 193082
rect 175917 193024 175922 193080
rect 175978 193024 198780 193080
rect 175917 193022 198780 193024
rect 175917 193019 175983 193022
rect 198774 193020 198780 193022
rect 198844 193020 198850 193084
rect 201534 192946 201540 192948
rect 174862 192886 201540 192946
rect 201534 192884 201540 192886
rect 201604 192884 201610 192948
rect 202873 192810 202939 192813
rect 174678 192808 202939 192810
rect 174678 192752 202878 192808
rect 202934 192752 202939 192808
rect 174678 192750 202939 192752
rect 202873 192747 202939 192750
rect 152733 192674 152799 192677
rect 186078 192674 186084 192676
rect 152733 192672 186084 192674
rect 152733 192616 152738 192672
rect 152794 192616 186084 192672
rect 152733 192614 186084 192616
rect 152733 192611 152799 192614
rect 186078 192612 186084 192614
rect 186148 192612 186154 192676
rect 103094 192476 103100 192540
rect 103164 192538 103170 192540
rect 131021 192538 131087 192541
rect 103164 192536 131087 192538
rect 103164 192480 131026 192536
rect 131082 192480 131087 192536
rect 103164 192478 131087 192480
rect 103164 192476 103170 192478
rect 131021 192475 131087 192478
rect 153837 192538 153903 192541
rect 209313 192538 209379 192541
rect 153837 192536 209379 192538
rect 153837 192480 153842 192536
rect 153898 192480 209318 192536
rect 209374 192480 209379 192536
rect 153837 192478 209379 192480
rect 153837 192475 153903 192478
rect 209313 192475 209379 192478
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect 168373 192266 168439 192269
rect 175917 192266 175983 192269
rect 168373 192264 175983 192266
rect 168373 192208 168378 192264
rect 168434 192208 175922 192264
rect 175978 192208 175983 192264
rect 168373 192206 175983 192208
rect 168373 192203 168439 192206
rect 175917 192203 175983 192206
rect 170029 192130 170095 192133
rect 174537 192130 174603 192133
rect 170029 192128 174603 192130
rect 170029 192072 170034 192128
rect 170090 192072 174542 192128
rect 174598 192072 174603 192128
rect 170029 192070 174603 192072
rect 170029 192067 170095 192070
rect 174537 192067 174603 192070
rect 101857 191722 101923 191725
rect 134006 191722 134012 191724
rect 101857 191720 134012 191722
rect 101857 191664 101862 191720
rect 101918 191664 134012 191720
rect 101857 191662 134012 191664
rect 101857 191659 101923 191662
rect 134006 191660 134012 191662
rect 134076 191660 134082 191724
rect 101765 191586 101831 191589
rect 132953 191586 133019 191589
rect 101765 191584 133019 191586
rect 101765 191528 101770 191584
rect 101826 191528 132958 191584
rect 133014 191528 133019 191584
rect 101765 191526 133019 191528
rect 101765 191523 101831 191526
rect 132953 191523 133019 191526
rect 102041 191450 102107 191453
rect 135478 191450 135484 191452
rect 102041 191448 135484 191450
rect 102041 191392 102046 191448
rect 102102 191392 135484 191448
rect 102041 191390 135484 191392
rect 102041 191387 102107 191390
rect 135478 191388 135484 191390
rect 135548 191388 135554 191452
rect 100661 191314 100727 191317
rect 134190 191314 134196 191316
rect 100661 191312 134196 191314
rect 100661 191256 100666 191312
rect 100722 191256 134196 191312
rect 100661 191254 134196 191256
rect 100661 191251 100727 191254
rect 134190 191252 134196 191254
rect 134260 191252 134266 191316
rect 106089 191178 106155 191181
rect 139710 191178 139716 191180
rect 106089 191176 139716 191178
rect 106089 191120 106094 191176
rect 106150 191120 139716 191176
rect 106089 191118 139716 191120
rect 106089 191115 106155 191118
rect 139710 191116 139716 191118
rect 139780 191116 139786 191180
rect 168557 191178 168623 191181
rect 185342 191178 185348 191180
rect 168557 191176 185348 191178
rect 168557 191120 168562 191176
rect 168618 191120 185348 191176
rect 168557 191118 185348 191120
rect 168557 191115 168623 191118
rect 185342 191116 185348 191118
rect 185412 191116 185418 191180
rect 101949 191042 102015 191045
rect 135662 191042 135668 191044
rect 101949 191040 135668 191042
rect 101949 190984 101954 191040
rect 102010 190984 135668 191040
rect 101949 190982 135668 190984
rect 101949 190979 102015 190982
rect 135662 190980 135668 190982
rect 135732 190980 135738 191044
rect 164918 190980 164924 191044
rect 164988 191042 164994 191044
rect 205633 191042 205699 191045
rect 164988 191040 205699 191042
rect 164988 190984 205638 191040
rect 205694 190984 205699 191040
rect 164988 190982 205699 190984
rect 164988 190980 164994 190982
rect 205633 190979 205699 190982
rect 107469 190090 107535 190093
rect 138422 190090 138428 190092
rect 107469 190088 138428 190090
rect 107469 190032 107474 190088
rect 107530 190032 138428 190088
rect 107469 190030 138428 190032
rect 107469 190027 107535 190030
rect 138422 190028 138428 190030
rect 138492 190028 138498 190092
rect 172278 190028 172284 190092
rect 172348 190090 172354 190092
rect 206185 190090 206251 190093
rect 172348 190088 206251 190090
rect 172348 190032 206190 190088
rect 206246 190032 206251 190088
rect 172348 190030 206251 190032
rect 172348 190028 172354 190030
rect 206185 190027 206251 190030
rect 100518 189892 100524 189956
rect 100588 189954 100594 189956
rect 133321 189954 133387 189957
rect 100588 189952 133387 189954
rect 100588 189896 133326 189952
rect 133382 189896 133387 189952
rect 100588 189894 133387 189896
rect 100588 189892 100594 189894
rect 133321 189891 133387 189894
rect 177113 189954 177179 189957
rect 211245 189954 211311 189957
rect 177113 189952 211311 189954
rect 177113 189896 177118 189952
rect 177174 189896 211250 189952
rect 211306 189896 211311 189952
rect 177113 189894 211311 189896
rect 177113 189891 177179 189894
rect 211245 189891 211311 189894
rect 104198 189756 104204 189820
rect 104268 189818 104274 189820
rect 136950 189818 136956 189820
rect 104268 189758 136956 189818
rect 104268 189756 104274 189758
rect 136950 189756 136956 189758
rect 137020 189756 137026 189820
rect 175641 189818 175707 189821
rect 210233 189818 210299 189821
rect 175641 189816 210299 189818
rect 175641 189760 175646 189816
rect 175702 189760 210238 189816
rect 210294 189760 210299 189816
rect 175641 189758 210299 189760
rect 175641 189755 175707 189758
rect 210233 189755 210299 189758
rect 104709 189682 104775 189685
rect 138238 189682 138244 189684
rect 104709 189680 138244 189682
rect 104709 189624 104714 189680
rect 104770 189624 138244 189680
rect 104709 189622 138244 189624
rect 104709 189619 104775 189622
rect 138238 189620 138244 189622
rect 138308 189620 138314 189684
rect 158110 189620 158116 189684
rect 158180 189682 158186 189684
rect 212533 189682 212599 189685
rect 158180 189680 212599 189682
rect 158180 189624 212538 189680
rect 212594 189624 212599 189680
rect 158180 189622 212599 189624
rect 158180 189620 158186 189622
rect 212533 189619 212599 189622
rect -960 188866 480 188956
rect 3417 188866 3483 188869
rect -960 188864 3483 188866
rect -960 188808 3422 188864
rect 3478 188808 3483 188864
rect -960 188806 3483 188808
rect -960 188716 480 188806
rect 3417 188803 3483 188806
rect 108430 187172 108436 187236
rect 108500 187234 108506 187236
rect 138565 187234 138631 187237
rect 108500 187232 138631 187234
rect 108500 187176 138570 187232
rect 138626 187176 138631 187232
rect 108500 187174 138631 187176
rect 108500 187172 108506 187174
rect 138565 187171 138631 187174
rect 108246 187036 108252 187100
rect 108316 187098 108322 187100
rect 139945 187098 140011 187101
rect 108316 187096 140011 187098
rect 108316 187040 139950 187096
rect 140006 187040 140011 187096
rect 108316 187038 140011 187040
rect 108316 187036 108322 187038
rect 139945 187035 140011 187038
rect 157006 187036 157012 187100
rect 157076 187098 157082 187100
rect 204253 187098 204319 187101
rect 157076 187096 204319 187098
rect 157076 187040 204258 187096
rect 204314 187040 204319 187096
rect 157076 187038 204319 187040
rect 157076 187036 157082 187038
rect 204253 187035 204319 187038
rect 107561 186962 107627 186965
rect 139526 186962 139532 186964
rect 107561 186960 139532 186962
rect 107561 186904 107566 186960
rect 107622 186904 139532 186960
rect 107561 186902 139532 186904
rect 107561 186899 107627 186902
rect 139526 186900 139532 186902
rect 139596 186900 139602 186964
rect 152958 186900 152964 186964
rect 153028 186962 153034 186964
rect 218053 186962 218119 186965
rect 153028 186960 218119 186962
rect 153028 186904 218058 186960
rect 218114 186904 218119 186960
rect 153028 186902 218119 186904
rect 153028 186900 153034 186902
rect 218053 186899 218119 186902
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3509 162890 3575 162893
rect -960 162888 3575 162890
rect -960 162832 3514 162888
rect 3570 162832 3575 162888
rect -960 162830 3575 162832
rect -960 162740 480 162830
rect 3509 162827 3575 162830
rect 169150 155620 169156 155684
rect 169220 155682 169226 155684
rect 203241 155682 203307 155685
rect 169220 155680 203307 155682
rect 169220 155624 203246 155680
rect 203302 155624 203307 155680
rect 169220 155622 203307 155624
rect 169220 155620 169226 155622
rect 203241 155619 203307 155622
rect 169334 155484 169340 155548
rect 169404 155546 169410 155548
rect 203149 155546 203215 155549
rect 169404 155544 203215 155546
rect 169404 155488 203154 155544
rect 203210 155488 203215 155544
rect 169404 155486 203215 155488
rect 169404 155484 169410 155486
rect 203149 155483 203215 155486
rect 176326 155348 176332 155412
rect 176396 155410 176402 155412
rect 216857 155410 216923 155413
rect 176396 155408 216923 155410
rect 176396 155352 216862 155408
rect 216918 155352 216923 155408
rect 176396 155350 216923 155352
rect 176396 155348 176402 155350
rect 216857 155347 216923 155350
rect 161238 155212 161244 155276
rect 161308 155274 161314 155276
rect 203333 155274 203399 155277
rect 161308 155272 203399 155274
rect 161308 155216 203338 155272
rect 203394 155216 203399 155272
rect 161308 155214 203399 155216
rect 161308 155212 161314 155214
rect 203333 155211 203399 155214
rect 579981 152690 580047 152693
rect 583520 152690 584960 152780
rect 579981 152688 584960 152690
rect 579981 152632 579986 152688
rect 580042 152632 584960 152688
rect 579981 152630 584960 152632
rect 579981 152627 580047 152630
rect 583520 152540 584960 152630
rect 148910 152356 148916 152420
rect 148980 152418 148986 152420
rect 186037 152418 186103 152421
rect 148980 152416 186103 152418
rect 148980 152360 186042 152416
rect 186098 152360 186103 152416
rect 148980 152358 186103 152360
rect 148980 152356 148986 152358
rect 186037 152355 186103 152358
rect 124070 151676 124076 151740
rect 124140 151738 124146 151740
rect 138473 151738 138539 151741
rect 124140 151736 138539 151738
rect 124140 151680 138478 151736
rect 138534 151680 138539 151736
rect 124140 151678 138539 151680
rect 124140 151676 124146 151678
rect 138473 151675 138539 151678
rect 122741 151602 122807 151605
rect 141049 151602 141115 151605
rect 122741 151600 141115 151602
rect 122741 151544 122746 151600
rect 122802 151544 141054 151600
rect 141110 151544 141115 151600
rect 122741 151542 141115 151544
rect 122741 151539 122807 151542
rect 141049 151539 141115 151542
rect 108798 151404 108804 151468
rect 108868 151466 108874 151468
rect 137461 151466 137527 151469
rect 108868 151464 137527 151466
rect 108868 151408 137466 151464
rect 137522 151408 137527 151464
rect 108868 151406 137527 151408
rect 108868 151404 108874 151406
rect 137461 151403 137527 151406
rect 167177 151466 167243 151469
rect 190494 151466 190500 151468
rect 167177 151464 190500 151466
rect 167177 151408 167182 151464
rect 167238 151408 190500 151464
rect 167177 151406 190500 151408
rect 167177 151403 167243 151406
rect 190494 151404 190500 151406
rect 190564 151404 190570 151468
rect 105445 151330 105511 151333
rect 136766 151330 136772 151332
rect 105445 151328 136772 151330
rect 105445 151272 105450 151328
rect 105506 151272 136772 151328
rect 105445 151270 136772 151272
rect 105445 151267 105511 151270
rect 136766 151268 136772 151270
rect 136836 151268 136842 151332
rect 153653 151330 153719 151333
rect 187734 151330 187740 151332
rect 153653 151328 187740 151330
rect 153653 151272 153658 151328
rect 153714 151272 187740 151328
rect 153653 151270 187740 151272
rect 153653 151267 153719 151270
rect 187734 151268 187740 151270
rect 187804 151268 187810 151332
rect 105353 151194 105419 151197
rect 138054 151194 138060 151196
rect 105353 151192 138060 151194
rect 105353 151136 105358 151192
rect 105414 151136 138060 151192
rect 105353 151134 138060 151136
rect 105353 151131 105419 151134
rect 138054 151132 138060 151134
rect 138124 151132 138130 151196
rect 154430 151132 154436 151196
rect 154500 151194 154506 151196
rect 200941 151194 201007 151197
rect 154500 151192 201007 151194
rect 154500 151136 200946 151192
rect 201002 151136 201007 151192
rect 154500 151134 201007 151136
rect 154500 151132 154506 151134
rect 200941 151131 201007 151134
rect 102777 151058 102843 151061
rect 136582 151058 136588 151060
rect 102777 151056 136588 151058
rect 102777 151000 102782 151056
rect 102838 151000 136588 151056
rect 102777 150998 136588 151000
rect 102777 150995 102843 150998
rect 136582 150996 136588 150998
rect 136652 150996 136658 151060
rect 162342 150996 162348 151060
rect 162412 151058 162418 151060
rect 214649 151058 214715 151061
rect 162412 151056 214715 151058
rect 162412 151000 214654 151056
rect 214710 151000 214715 151056
rect 162412 150998 214715 151000
rect 162412 150996 162418 150998
rect 214649 150995 214715 150998
rect 185853 150514 185919 150517
rect 191966 150514 191972 150516
rect 185853 150512 191972 150514
rect 185853 150456 185858 150512
rect 185914 150456 191972 150512
rect 185853 150454 191972 150456
rect 185853 150451 185919 150454
rect 191966 150452 191972 150454
rect 192036 150452 192042 150516
rect 174169 150378 174235 150381
rect 202086 150378 202092 150380
rect 174169 150376 202092 150378
rect 174169 150320 174174 150376
rect 174230 150320 202092 150376
rect 174169 150318 202092 150320
rect 174169 150315 174235 150318
rect 202086 150316 202092 150318
rect 202156 150316 202162 150380
rect 207606 150316 207612 150380
rect 207676 150378 207682 150380
rect 207749 150378 207815 150381
rect 207676 150376 207815 150378
rect 207676 150320 207754 150376
rect 207810 150320 207815 150376
rect 207676 150318 207815 150320
rect 207676 150316 207682 150318
rect 207749 150315 207815 150318
rect 176510 150180 176516 150244
rect 176580 150242 176586 150244
rect 204437 150242 204503 150245
rect 176580 150240 204503 150242
rect 176580 150184 204442 150240
rect 204498 150184 204503 150240
rect 176580 150182 204503 150184
rect 176580 150180 176586 150182
rect 204437 150179 204503 150182
rect 174353 150106 174419 150109
rect 203006 150106 203012 150108
rect 174353 150104 203012 150106
rect 174353 150048 174358 150104
rect 174414 150048 203012 150104
rect 174353 150046 203012 150048
rect 174353 150043 174419 150046
rect 203006 150044 203012 150046
rect 203076 150044 203082 150108
rect -960 149834 480 149924
rect 173750 149908 173756 149972
rect 173820 149970 173826 149972
rect 202822 149970 202828 149972
rect 173820 149910 202828 149970
rect 173820 149908 173826 149910
rect 202822 149908 202828 149910
rect 202892 149908 202898 149972
rect 3141 149834 3207 149837
rect -960 149832 3207 149834
rect -960 149776 3146 149832
rect 3202 149776 3207 149832
rect -960 149774 3207 149776
rect -960 149684 480 149774
rect 3141 149771 3207 149774
rect 113398 149772 113404 149836
rect 113468 149834 113474 149836
rect 140865 149834 140931 149837
rect 113468 149832 140931 149834
rect 113468 149776 140870 149832
rect 140926 149776 140931 149832
rect 113468 149774 140931 149776
rect 113468 149772 113474 149774
rect 140865 149771 140931 149774
rect 176653 149834 176719 149837
rect 205766 149834 205772 149836
rect 176653 149832 205772 149834
rect 176653 149776 176658 149832
rect 176714 149776 205772 149832
rect 176653 149774 205772 149776
rect 176653 149771 176719 149774
rect 205766 149772 205772 149774
rect 205836 149772 205842 149836
rect 101397 149698 101463 149701
rect 135294 149698 135300 149700
rect 101397 149696 135300 149698
rect 101397 149640 101402 149696
rect 101458 149640 135300 149696
rect 101397 149638 135300 149640
rect 101397 149635 101463 149638
rect 135294 149636 135300 149638
rect 135364 149636 135370 149700
rect 175457 149698 175523 149701
rect 205582 149698 205588 149700
rect 175457 149696 205588 149698
rect 175457 149640 175462 149696
rect 175518 149640 205588 149696
rect 175457 149638 205588 149640
rect 175457 149635 175523 149638
rect 205582 149636 205588 149638
rect 205652 149636 205658 149700
rect 167085 149562 167151 149565
rect 187734 149562 187740 149564
rect 167085 149560 187740 149562
rect 167085 149504 167090 149560
rect 167146 149504 187740 149560
rect 167085 149502 187740 149504
rect 167085 149499 167151 149502
rect 187734 149500 187740 149502
rect 187804 149500 187810 149564
rect 203374 149092 203380 149156
rect 203444 149154 203450 149156
rect 203609 149154 203675 149157
rect 203444 149152 203675 149154
rect 203444 149096 203614 149152
rect 203670 149096 203675 149152
rect 203444 149094 203675 149096
rect 203444 149092 203450 149094
rect 203609 149091 203675 149094
rect 136173 149018 136239 149021
rect 188429 149018 188495 149021
rect 136173 149016 188495 149018
rect 136173 148960 136178 149016
rect 136234 148960 188434 149016
rect 188490 148960 188495 149016
rect 136173 148958 188495 148960
rect 136173 148955 136239 148958
rect 188429 148955 188495 148958
rect 104382 148820 104388 148884
rect 104452 148882 104458 148884
rect 135713 148882 135779 148885
rect 104452 148880 135779 148882
rect 104452 148824 135718 148880
rect 135774 148824 135779 148880
rect 104452 148822 135779 148824
rect 104452 148820 104458 148822
rect 135713 148819 135779 148822
rect 120758 148684 120764 148748
rect 120828 148746 120834 148748
rect 153561 148746 153627 148749
rect 120828 148744 153627 148746
rect 120828 148688 153566 148744
rect 153622 148688 153627 148744
rect 120828 148686 153627 148688
rect 120828 148684 120834 148686
rect 153561 148683 153627 148686
rect 115422 148548 115428 148612
rect 115492 148610 115498 148612
rect 149237 148610 149303 148613
rect 115492 148608 149303 148610
rect 115492 148552 149242 148608
rect 149298 148552 149303 148608
rect 115492 148550 149303 148552
rect 115492 148548 115498 148550
rect 149237 148547 149303 148550
rect 157885 148610 157951 148613
rect 188245 148610 188311 148613
rect 157885 148608 188311 148610
rect 157885 148552 157890 148608
rect 157946 148552 188250 148608
rect 188306 148552 188311 148608
rect 157885 148550 188311 148552
rect 157885 148547 157951 148550
rect 188245 148547 188311 148550
rect 117814 148412 117820 148476
rect 117884 148474 117890 148476
rect 151997 148474 152063 148477
rect 117884 148472 152063 148474
rect 117884 148416 152002 148472
rect 152058 148416 152063 148472
rect 117884 148414 152063 148416
rect 117884 148412 117890 148414
rect 151997 148411 152063 148414
rect 166993 148474 167059 148477
rect 202045 148474 202111 148477
rect 166993 148472 202111 148474
rect 166993 148416 166998 148472
rect 167054 148416 202050 148472
rect 202106 148416 202111 148472
rect 166993 148414 202111 148416
rect 166993 148411 167059 148414
rect 202045 148411 202111 148414
rect 113582 148276 113588 148340
rect 113652 148338 113658 148340
rect 148593 148338 148659 148341
rect 113652 148336 148659 148338
rect 113652 148280 148598 148336
rect 148654 148280 148659 148336
rect 113652 148278 148659 148280
rect 113652 148276 113658 148278
rect 148593 148275 148659 148278
rect 151721 148338 151787 148341
rect 200481 148338 200547 148341
rect 151721 148336 200547 148338
rect 151721 148280 151726 148336
rect 151782 148280 200486 148336
rect 200542 148280 200547 148336
rect 151721 148278 200547 148280
rect 151721 148275 151787 148278
rect 200481 148275 200547 148278
rect 122230 148140 122236 148204
rect 122300 148202 122306 148204
rect 151905 148202 151971 148205
rect 122300 148200 151971 148202
rect 122300 148144 151910 148200
rect 151966 148144 151971 148200
rect 122300 148142 151971 148144
rect 122300 148140 122306 148142
rect 151905 148139 151971 148142
rect 122005 148066 122071 148069
rect 142286 148066 142292 148068
rect 122005 148064 142292 148066
rect 122005 148008 122010 148064
rect 122066 148008 142292 148064
rect 122005 148006 142292 148008
rect 122005 148003 122071 148006
rect 142286 148004 142292 148006
rect 142356 148004 142362 148068
rect 122046 147732 122052 147796
rect 122116 147794 122122 147796
rect 122557 147794 122623 147797
rect 122116 147792 122623 147794
rect 122116 147736 122562 147792
rect 122618 147736 122623 147792
rect 122116 147734 122623 147736
rect 122116 147732 122122 147734
rect 122557 147731 122623 147734
rect 120441 147658 120507 147661
rect 139342 147658 139348 147660
rect 120441 147656 139348 147658
rect 120441 147600 120446 147656
rect 120502 147600 139348 147656
rect 120441 147598 139348 147600
rect 120441 147595 120507 147598
rect 139342 147596 139348 147598
rect 139412 147596 139418 147660
rect 170305 147658 170371 147661
rect 192150 147658 192156 147660
rect 170305 147656 192156 147658
rect 170305 147600 170310 147656
rect 170366 147600 192156 147656
rect 170305 147598 192156 147600
rect 170305 147595 170371 147598
rect 192150 147596 192156 147598
rect 192220 147596 192226 147660
rect 112294 147460 112300 147524
rect 112364 147522 112370 147524
rect 132217 147522 132283 147525
rect 112364 147520 132283 147522
rect 112364 147464 132222 147520
rect 132278 147464 132283 147520
rect 112364 147462 132283 147464
rect 112364 147460 112370 147462
rect 132217 147459 132283 147462
rect 171133 147522 171199 147525
rect 194726 147522 194732 147524
rect 171133 147520 194732 147522
rect 171133 147464 171138 147520
rect 171194 147464 194732 147520
rect 171133 147462 194732 147464
rect 171133 147459 171199 147462
rect 194726 147460 194732 147462
rect 194796 147460 194802 147524
rect 196433 147522 196499 147525
rect 196566 147522 196572 147524
rect 196433 147520 196572 147522
rect 196433 147464 196438 147520
rect 196494 147464 196572 147520
rect 196433 147462 196572 147464
rect 196433 147459 196499 147462
rect 196566 147460 196572 147462
rect 196636 147460 196642 147524
rect 110822 147324 110828 147388
rect 110892 147386 110898 147388
rect 131849 147386 131915 147389
rect 110892 147384 131915 147386
rect 110892 147328 131854 147384
rect 131910 147328 131915 147384
rect 110892 147326 131915 147328
rect 110892 147324 110898 147326
rect 131849 147323 131915 147326
rect 169937 147386 170003 147389
rect 193806 147386 193812 147388
rect 169937 147384 193812 147386
rect 169937 147328 169942 147384
rect 169998 147328 193812 147384
rect 169937 147326 193812 147328
rect 169937 147323 170003 147326
rect 193806 147324 193812 147326
rect 193876 147324 193882 147388
rect 115054 147188 115060 147252
rect 115124 147250 115130 147252
rect 137093 147250 137159 147253
rect 115124 147248 137159 147250
rect 115124 147192 137098 147248
rect 137154 147192 137159 147248
rect 115124 147190 137159 147192
rect 115124 147188 115130 147190
rect 137093 147187 137159 147190
rect 170121 147250 170187 147253
rect 196198 147250 196204 147252
rect 170121 147248 196204 147250
rect 170121 147192 170126 147248
rect 170182 147192 196204 147248
rect 170121 147190 196204 147192
rect 170121 147187 170187 147190
rect 196198 147188 196204 147190
rect 196268 147188 196274 147252
rect 112662 147052 112668 147116
rect 112732 147114 112738 147116
rect 143574 147114 143580 147116
rect 112732 147054 143580 147114
rect 112732 147052 112738 147054
rect 143574 147052 143580 147054
rect 143644 147052 143650 147116
rect 171317 147114 171383 147117
rect 197854 147114 197860 147116
rect 171317 147112 197860 147114
rect 171317 147056 171322 147112
rect 171378 147056 197860 147112
rect 171317 147054 197860 147056
rect 171317 147051 171383 147054
rect 197854 147052 197860 147054
rect 197924 147052 197930 147116
rect 110965 146978 111031 146981
rect 142470 146978 142476 146980
rect 110965 146976 142476 146978
rect 110965 146920 110970 146976
rect 111026 146920 142476 146976
rect 110965 146918 142476 146920
rect 110965 146915 111031 146918
rect 142470 146916 142476 146918
rect 142540 146916 142546 146980
rect 157190 146916 157196 146980
rect 157260 146978 157266 146980
rect 189901 146978 189967 146981
rect 157260 146976 189967 146978
rect 157260 146920 189906 146976
rect 189962 146920 189967 146976
rect 157260 146918 189967 146920
rect 157260 146916 157266 146918
rect 189901 146915 189967 146918
rect 113950 146780 113956 146844
rect 114020 146842 114026 146844
rect 130653 146842 130719 146845
rect 114020 146840 130719 146842
rect 114020 146784 130658 146840
rect 130714 146784 130719 146840
rect 114020 146782 130719 146784
rect 114020 146780 114026 146782
rect 130653 146779 130719 146782
rect 179413 146842 179479 146845
rect 197670 146842 197676 146844
rect 179413 146840 197676 146842
rect 179413 146784 179418 146840
rect 179474 146784 197676 146840
rect 179413 146782 197676 146784
rect 179413 146779 179479 146782
rect 197670 146780 197676 146782
rect 197740 146780 197746 146844
rect 198733 146842 198799 146845
rect 199510 146842 199516 146844
rect 198733 146840 199516 146842
rect 198733 146784 198738 146840
rect 198794 146784 199516 146840
rect 198733 146782 199516 146784
rect 198733 146779 198799 146782
rect 199510 146780 199516 146782
rect 199580 146780 199586 146844
rect 122741 146708 122807 146709
rect 122741 146704 122788 146708
rect 122852 146706 122858 146708
rect 122741 146648 122746 146704
rect 122741 146644 122788 146648
rect 122852 146646 122898 146706
rect 122852 146644 122858 146646
rect 122741 146643 122807 146644
rect 109350 146236 109356 146300
rect 109420 146298 109426 146300
rect 129825 146298 129891 146301
rect 109420 146296 129891 146298
rect 109420 146240 129830 146296
rect 129886 146240 129891 146296
rect 109420 146238 129891 146240
rect 109420 146236 109426 146238
rect 129825 146235 129891 146238
rect 199326 146236 199332 146300
rect 199396 146298 199402 146300
rect 199745 146298 199811 146301
rect 199396 146296 199811 146298
rect 199396 146240 199750 146296
rect 199806 146240 199811 146296
rect 199396 146238 199811 146240
rect 199396 146236 199402 146238
rect 199745 146235 199811 146238
rect 109534 146100 109540 146164
rect 109604 146162 109610 146164
rect 135805 146162 135871 146165
rect 109604 146160 135871 146162
rect 109604 146104 135810 146160
rect 135866 146104 135871 146160
rect 109604 146102 135871 146104
rect 109604 146100 109610 146102
rect 135805 146099 135871 146102
rect 176469 146162 176535 146165
rect 197670 146162 197676 146164
rect 176469 146160 197676 146162
rect 176469 146104 176474 146160
rect 176530 146104 197676 146160
rect 176469 146102 197676 146104
rect 176469 146099 176535 146102
rect 197670 146100 197676 146102
rect 197740 146100 197746 146164
rect 116158 145964 116164 146028
rect 116228 146026 116234 146028
rect 147070 146026 147076 146028
rect 116228 145966 147076 146026
rect 116228 145964 116234 145966
rect 147070 145964 147076 145966
rect 147140 145964 147146 146028
rect 172513 146026 172579 146029
rect 196014 146026 196020 146028
rect 172513 146024 196020 146026
rect 172513 145968 172518 146024
rect 172574 145968 196020 146024
rect 172513 145966 196020 145968
rect 172513 145963 172579 145966
rect 196014 145964 196020 145966
rect 196084 145964 196090 146028
rect 115790 145828 115796 145892
rect 115860 145890 115866 145892
rect 149053 145890 149119 145893
rect 115860 145888 149119 145890
rect 115860 145832 149058 145888
rect 149114 145832 149119 145888
rect 115860 145830 149119 145832
rect 115860 145828 115866 145830
rect 149053 145827 149119 145830
rect 173893 145890 173959 145893
rect 199142 145890 199148 145892
rect 173893 145888 199148 145890
rect 173893 145832 173898 145888
rect 173954 145832 199148 145888
rect 173893 145830 199148 145832
rect 173893 145827 173959 145830
rect 199142 145828 199148 145830
rect 199212 145828 199218 145892
rect 119654 145692 119660 145756
rect 119724 145754 119730 145756
rect 153469 145754 153535 145757
rect 119724 145752 153535 145754
rect 119724 145696 153474 145752
rect 153530 145696 153535 145752
rect 119724 145694 153535 145696
rect 119724 145692 119730 145694
rect 153469 145691 153535 145694
rect 171777 145754 171843 145757
rect 199469 145754 199535 145757
rect 171777 145752 199535 145754
rect 171777 145696 171782 145752
rect 171838 145696 199474 145752
rect 199530 145696 199535 145752
rect 171777 145694 199535 145696
rect 171777 145691 171843 145694
rect 199469 145691 199535 145694
rect 112846 145556 112852 145620
rect 112916 145618 112922 145620
rect 147765 145618 147831 145621
rect 112916 145616 147831 145618
rect 112916 145560 147770 145616
rect 147826 145560 147831 145616
rect 112916 145558 147831 145560
rect 112916 145556 112922 145558
rect 147765 145555 147831 145558
rect 163037 145618 163103 145621
rect 196893 145618 196959 145621
rect 163037 145616 196959 145618
rect 163037 145560 163042 145616
rect 163098 145560 196898 145616
rect 196954 145560 196959 145616
rect 163037 145558 196959 145560
rect 163037 145555 163103 145558
rect 196893 145555 196959 145558
rect 111190 145420 111196 145484
rect 111260 145482 111266 145484
rect 131113 145482 131179 145485
rect 111260 145480 131179 145482
rect 111260 145424 131118 145480
rect 131174 145424 131179 145480
rect 111260 145422 131179 145424
rect 111260 145420 111266 145422
rect 131113 145419 131179 145422
rect 180333 144802 180399 144805
rect 193990 144802 193996 144804
rect 180333 144800 193996 144802
rect 180333 144744 180338 144800
rect 180394 144744 193996 144800
rect 180333 144742 193996 144744
rect 180333 144739 180399 144742
rect 193990 144740 193996 144742
rect 194060 144740 194066 144804
rect 114134 144604 114140 144668
rect 114204 144666 114210 144668
rect 138657 144666 138723 144669
rect 114204 144664 138723 144666
rect 114204 144608 138662 144664
rect 138718 144608 138723 144664
rect 114204 144606 138723 144608
rect 114204 144604 114210 144606
rect 138657 144603 138723 144606
rect 164325 144666 164391 144669
rect 189574 144666 189580 144668
rect 164325 144664 189580 144666
rect 164325 144608 164330 144664
rect 164386 144608 189580 144664
rect 164325 144606 189580 144608
rect 164325 144603 164391 144606
rect 189574 144604 189580 144606
rect 189644 144604 189650 144668
rect 120809 144530 120875 144533
rect 147673 144530 147739 144533
rect 120809 144528 147739 144530
rect 120809 144472 120814 144528
rect 120870 144472 147678 144528
rect 147734 144472 147739 144528
rect 120809 144470 147739 144472
rect 120809 144467 120875 144470
rect 147673 144467 147739 144470
rect 168005 144530 168071 144533
rect 198958 144530 198964 144532
rect 168005 144528 198964 144530
rect 168005 144472 168010 144528
rect 168066 144472 198964 144528
rect 168005 144470 198964 144472
rect 168005 144467 168071 144470
rect 198958 144468 198964 144470
rect 199028 144468 199034 144532
rect 111558 144332 111564 144396
rect 111628 144394 111634 144396
rect 142521 144394 142587 144397
rect 111628 144392 142587 144394
rect 111628 144336 142526 144392
rect 142582 144336 142587 144392
rect 111628 144334 142587 144336
rect 111628 144332 111634 144334
rect 142521 144331 142587 144334
rect 162485 144394 162551 144397
rect 193438 144394 193444 144396
rect 162485 144392 193444 144394
rect 162485 144336 162490 144392
rect 162546 144336 193444 144392
rect 162485 144334 193444 144336
rect 162485 144331 162551 144334
rect 193438 144332 193444 144334
rect 193508 144332 193514 144396
rect 116342 144196 116348 144260
rect 116412 144258 116418 144260
rect 148174 144258 148180 144260
rect 116412 144198 148180 144258
rect 116412 144196 116418 144198
rect 148174 144196 148180 144198
rect 148244 144196 148250 144260
rect 156137 144258 156203 144261
rect 189206 144258 189212 144260
rect 156137 144256 189212 144258
rect 156137 144200 156142 144256
rect 156198 144200 189212 144256
rect 156137 144198 189212 144200
rect 156137 144195 156203 144198
rect 189206 144196 189212 144198
rect 189276 144196 189282 144260
rect 115289 144122 115355 144125
rect 148593 144122 148659 144125
rect 115289 144120 148659 144122
rect 115289 144064 115294 144120
rect 115350 144064 148598 144120
rect 148654 144064 148659 144120
rect 115289 144062 148659 144064
rect 115289 144059 115355 144062
rect 148593 144059 148659 144062
rect 160829 144122 160895 144125
rect 193622 144122 193628 144124
rect 160829 144120 193628 144122
rect 160829 144064 160834 144120
rect 160890 144064 193628 144120
rect 160829 144062 193628 144064
rect 160829 144059 160895 144062
rect 193622 144060 193628 144062
rect 193692 144060 193698 144124
rect 116710 143924 116716 143988
rect 116780 143986 116786 143988
rect 116853 143986 116919 143989
rect 116780 143984 116919 143986
rect 116780 143928 116858 143984
rect 116914 143928 116919 143984
rect 116780 143926 116919 143928
rect 116780 143924 116786 143926
rect 116853 143923 116919 143926
rect 185669 143442 185735 143445
rect 187182 143442 187188 143444
rect 185669 143440 187188 143442
rect 185669 143384 185674 143440
rect 185730 143384 187188 143440
rect 185669 143382 187188 143384
rect 185669 143379 185735 143382
rect 187182 143380 187188 143382
rect 187252 143380 187258 143444
rect 111374 143244 111380 143308
rect 111444 143306 111450 143308
rect 125225 143306 125291 143309
rect 111444 143304 125291 143306
rect 111444 143248 125230 143304
rect 125286 143248 125291 143304
rect 111444 143246 125291 143248
rect 111444 143244 111450 143246
rect 125225 143243 125291 143246
rect 120993 143170 121059 143173
rect 121310 143170 121316 143172
rect 120993 143168 121316 143170
rect 120993 143112 120998 143168
rect 121054 143112 121316 143168
rect 120993 143110 121316 143112
rect 120993 143107 121059 143110
rect 121310 143108 121316 143110
rect 121380 143108 121386 143172
rect 185393 143170 185459 143173
rect 197077 143170 197143 143173
rect 185393 143168 197143 143170
rect 185393 143112 185398 143168
rect 185454 143112 197082 143168
rect 197138 143112 197143 143168
rect 185393 143110 197143 143112
rect 185393 143107 185459 143110
rect 197077 143107 197143 143110
rect 121126 142972 121132 143036
rect 121196 143034 121202 143036
rect 143073 143034 143139 143037
rect 121196 143032 143139 143034
rect 121196 142976 143078 143032
rect 143134 142976 143139 143032
rect 121196 142974 143139 142976
rect 121196 142972 121202 142974
rect 143073 142971 143139 142974
rect 165245 143034 165311 143037
rect 189625 143034 189691 143037
rect 165245 143032 189691 143034
rect 165245 142976 165250 143032
rect 165306 142976 189630 143032
rect 189686 142976 189691 143032
rect 165245 142974 189691 142976
rect 165245 142971 165311 142974
rect 189625 142971 189691 142974
rect 115606 142836 115612 142900
rect 115676 142898 115682 142900
rect 123569 142898 123635 142901
rect 115676 142896 123635 142898
rect 115676 142840 123574 142896
rect 123630 142840 123635 142896
rect 115676 142838 123635 142840
rect 115676 142836 115682 142838
rect 123569 142835 123635 142838
rect 130326 142836 130332 142900
rect 130396 142898 130402 142900
rect 159633 142898 159699 142901
rect 130396 142896 159699 142898
rect 130396 142840 159638 142896
rect 159694 142840 159699 142896
rect 130396 142838 159699 142840
rect 130396 142836 130402 142838
rect 159633 142835 159699 142838
rect 163589 142898 163655 142901
rect 190821 142898 190887 142901
rect 163589 142896 190887 142898
rect 163589 142840 163594 142896
rect 163650 142840 190826 142896
rect 190882 142840 190887 142896
rect 163589 142838 190887 142840
rect 163589 142835 163655 142838
rect 190821 142835 190887 142838
rect 118366 142700 118372 142764
rect 118436 142762 118442 142764
rect 151353 142762 151419 142765
rect 118436 142760 151419 142762
rect 118436 142704 151358 142760
rect 151414 142704 151419 142760
rect 118436 142702 151419 142704
rect 118436 142700 118442 142702
rect 151353 142699 151419 142702
rect 161933 142762 161999 142765
rect 190085 142762 190151 142765
rect 161933 142760 190151 142762
rect 161933 142704 161938 142760
rect 161994 142704 190090 142760
rect 190146 142704 190151 142760
rect 161933 142702 190151 142704
rect 161933 142699 161999 142702
rect 190085 142699 190151 142702
rect 121310 142564 121316 142628
rect 121380 142626 121386 142628
rect 185669 142626 185735 142629
rect 121380 142624 185735 142626
rect 121380 142568 185674 142624
rect 185730 142568 185735 142624
rect 121380 142566 185735 142568
rect 121380 142564 121386 142566
rect 185669 142563 185735 142566
rect 111006 142428 111012 142492
rect 111076 142490 111082 142492
rect 185393 142490 185459 142493
rect 111076 142488 185459 142490
rect 111076 142432 185398 142488
rect 185454 142432 185459 142488
rect 111076 142430 185459 142432
rect 111076 142428 111082 142430
rect 185393 142427 185459 142430
rect 126973 142354 127039 142357
rect 127801 142354 127867 142357
rect 467097 142354 467163 142357
rect 126973 142352 467163 142354
rect 126973 142296 126978 142352
rect 127034 142296 127806 142352
rect 127862 142296 467102 142352
rect 467158 142296 467163 142352
rect 126973 142294 467163 142296
rect 126973 142291 127039 142294
rect 127801 142291 127867 142294
rect 467097 142291 467163 142294
rect 116485 142218 116551 142221
rect 123937 142218 124003 142221
rect 580349 142218 580415 142221
rect 116485 142216 580415 142218
rect 116485 142160 116490 142216
rect 116546 142160 123942 142216
rect 123998 142160 580354 142216
rect 580410 142160 580415 142216
rect 116485 142158 580415 142160
rect 116485 142155 116551 142158
rect 123937 142155 124003 142158
rect 580349 142155 580415 142158
rect 115013 142082 115079 142085
rect 125593 142082 125659 142085
rect 115013 142080 125659 142082
rect 115013 142024 115018 142080
rect 115074 142024 125598 142080
rect 125654 142024 125659 142080
rect 115013 142022 125659 142024
rect 115013 142019 115079 142022
rect 125593 142019 125659 142022
rect 157333 142082 157399 142085
rect 190177 142082 190243 142085
rect 157333 142080 190243 142082
rect 157333 142024 157338 142080
rect 157394 142024 190182 142080
rect 190238 142024 190243 142080
rect 157333 142022 190243 142024
rect 157333 142019 157399 142022
rect 190177 142019 190243 142022
rect 116894 141884 116900 141948
rect 116964 141946 116970 141948
rect 123385 141946 123451 141949
rect 116964 141944 123451 141946
rect 116964 141888 123390 141944
rect 123446 141888 123451 141944
rect 116964 141886 123451 141888
rect 116964 141884 116970 141886
rect 123385 141883 123451 141886
rect 124581 141946 124647 141949
rect 125133 141946 125199 141949
rect 124581 141944 125199 141946
rect 124581 141888 124586 141944
rect 124642 141888 125138 141944
rect 125194 141888 125199 141944
rect 124581 141886 125199 141888
rect 124581 141883 124647 141886
rect 125133 141883 125199 141886
rect 112846 141612 112852 141676
rect 112916 141674 112922 141676
rect 140037 141674 140103 141677
rect 112916 141672 140103 141674
rect 112916 141616 140042 141672
rect 140098 141616 140103 141672
rect 112916 141614 140103 141616
rect 112916 141612 112922 141614
rect 140037 141611 140103 141614
rect 121126 141476 121132 141540
rect 121196 141538 121202 141540
rect 153285 141538 153351 141541
rect 121196 141536 153351 141538
rect 121196 141480 153290 141536
rect 153346 141480 153351 141536
rect 121196 141478 153351 141480
rect 121196 141476 121202 141478
rect 153285 141475 153351 141478
rect 174537 141538 174603 141541
rect 185894 141538 185900 141540
rect 174537 141536 185900 141538
rect 174537 141480 174542 141536
rect 174598 141480 185900 141536
rect 174537 141478 185900 141480
rect 174537 141475 174603 141478
rect 185894 141476 185900 141478
rect 185964 141476 185970 141540
rect 118182 141340 118188 141404
rect 118252 141402 118258 141404
rect 154021 141402 154087 141405
rect 118252 141400 154087 141402
rect 118252 141344 154026 141400
rect 154082 141344 154087 141400
rect 118252 141342 154087 141344
rect 118252 141340 118258 141342
rect 154021 141339 154087 141342
rect 157149 141402 157215 141405
rect 190729 141402 190795 141405
rect 157149 141400 190795 141402
rect 157149 141344 157154 141400
rect 157210 141344 190734 141400
rect 190790 141344 190795 141400
rect 157149 141342 190795 141344
rect 157149 141339 157215 141342
rect 190729 141339 190795 141342
rect 126513 141266 126579 141269
rect 464337 141266 464403 141269
rect 126513 141264 464403 141266
rect 126513 141208 126518 141264
rect 126574 141208 464342 141264
rect 464398 141208 464403 141264
rect 126513 141206 464403 141208
rect 126513 141203 126579 141206
rect 464337 141203 464403 141206
rect 124581 141130 124647 141133
rect 574737 141130 574803 141133
rect 124581 141128 574803 141130
rect 124581 141072 124586 141128
rect 124642 141072 574742 141128
rect 574798 141072 574803 141128
rect 124581 141070 574803 141072
rect 124581 141067 124647 141070
rect 574737 141067 574803 141070
rect 128445 140994 128511 140997
rect 580809 140994 580875 140997
rect 128445 140992 580875 140994
rect 128445 140936 128450 140992
rect 128506 140936 580814 140992
rect 580870 140936 580875 140992
rect 128445 140934 580875 140936
rect 128445 140931 128511 140934
rect 580809 140931 580875 140934
rect 127065 140858 127131 140861
rect 580625 140858 580691 140861
rect 127065 140856 580691 140858
rect 127065 140800 127070 140856
rect 127126 140800 580630 140856
rect 580686 140800 580691 140856
rect 127065 140798 580691 140800
rect 127065 140795 127131 140798
rect 580625 140795 580691 140798
rect 118785 140724 118851 140725
rect 118734 140722 118740 140724
rect 118694 140662 118740 140722
rect 118804 140720 118851 140724
rect 118846 140664 118851 140720
rect 118734 140660 118740 140662
rect 118804 140660 118851 140664
rect 120942 140660 120948 140724
rect 121012 140722 121018 140724
rect 127893 140722 127959 140725
rect 121012 140720 127959 140722
rect 121012 140664 127898 140720
rect 127954 140664 127959 140720
rect 121012 140662 127959 140664
rect 121012 140660 121018 140662
rect 118785 140659 118851 140660
rect 127893 140659 127959 140662
rect 119429 140586 119495 140589
rect 127709 140586 127775 140589
rect 119429 140584 127775 140586
rect 119429 140528 119434 140584
rect 119490 140528 127714 140584
rect 127770 140528 127775 140584
rect 119429 140526 127775 140528
rect 119429 140523 119495 140526
rect 127709 140523 127775 140526
rect 182817 140586 182883 140589
rect 187509 140586 187575 140589
rect 182817 140584 187575 140586
rect 182817 140528 182822 140584
rect 182878 140528 187514 140584
rect 187570 140528 187575 140584
rect 182817 140526 187575 140528
rect 182817 140523 182883 140526
rect 187509 140523 187575 140526
rect 119470 140388 119476 140452
rect 119540 140450 119546 140452
rect 128077 140450 128143 140453
rect 129089 140452 129155 140453
rect 129038 140450 129044 140452
rect 119540 140448 128143 140450
rect 119540 140392 128082 140448
rect 128138 140392 128143 140448
rect 119540 140390 128143 140392
rect 128998 140390 129044 140450
rect 129108 140448 129155 140452
rect 129150 140392 129155 140448
rect 119540 140388 119546 140390
rect 128077 140387 128143 140390
rect 129038 140388 129044 140390
rect 129108 140388 129155 140392
rect 129089 140387 129155 140388
rect 183185 140450 183251 140453
rect 191598 140450 191604 140452
rect 183185 140448 191604 140450
rect 183185 140392 183190 140448
rect 183246 140392 191604 140448
rect 183185 140390 191604 140392
rect 183185 140387 183251 140390
rect 191598 140388 191604 140390
rect 191668 140388 191674 140452
rect 124857 140316 124923 140317
rect 124806 140314 124812 140316
rect 124766 140254 124812 140314
rect 124876 140312 124923 140316
rect 124918 140256 124923 140312
rect 124806 140252 124812 140254
rect 124876 140252 124923 140256
rect 126830 140252 126836 140316
rect 126900 140314 126906 140316
rect 139853 140314 139919 140317
rect 126900 140312 139919 140314
rect 126900 140256 139858 140312
rect 139914 140256 139919 140312
rect 126900 140254 139919 140256
rect 126900 140252 126906 140254
rect 124857 140251 124923 140252
rect 139853 140251 139919 140254
rect 183001 140314 183067 140317
rect 190862 140314 190868 140316
rect 183001 140312 190868 140314
rect 183001 140256 183006 140312
rect 183062 140256 190868 140312
rect 183001 140254 190868 140256
rect 183001 140251 183067 140254
rect 190862 140252 190868 140254
rect 190932 140252 190938 140316
rect 119521 140178 119587 140181
rect 146518 140178 146524 140180
rect 119521 140176 146524 140178
rect 119521 140120 119526 140176
rect 119582 140120 146524 140176
rect 119521 140118 146524 140120
rect 119521 140115 119587 140118
rect 146518 140116 146524 140118
rect 146588 140116 146594 140180
rect 186262 140116 186268 140180
rect 186332 140178 186338 140180
rect 186497 140178 186563 140181
rect 186332 140176 186563 140178
rect 186332 140120 186502 140176
rect 186558 140120 186563 140176
rect 186332 140118 186563 140120
rect 186332 140116 186338 140118
rect 186497 140115 186563 140118
rect 146886 140042 146892 140044
rect 118650 139982 146892 140042
rect 116485 139906 116551 139909
rect 118650 139906 118710 139982
rect 146886 139980 146892 139982
rect 146956 139980 146962 140044
rect 169753 140042 169819 140045
rect 189390 140042 189396 140044
rect 169753 140040 189396 140042
rect 169753 139984 169758 140040
rect 169814 139984 189396 140040
rect 169753 139982 189396 139984
rect 169753 139979 169819 139982
rect 189390 139980 189396 139982
rect 189460 139980 189466 140044
rect 116485 139904 118710 139906
rect 116485 139848 116490 139904
rect 116546 139848 118710 139904
rect 116485 139846 118710 139848
rect 162577 139906 162643 139909
rect 195237 139906 195303 139909
rect 162577 139904 195303 139906
rect 162577 139848 162582 139904
rect 162638 139848 195242 139904
rect 195298 139848 195303 139904
rect 162577 139846 195303 139848
rect 116485 139843 116551 139846
rect 162577 139843 162643 139846
rect 195237 139843 195303 139846
rect 116526 139708 116532 139772
rect 116596 139770 116602 139772
rect 123385 139770 123451 139773
rect 116596 139768 123451 139770
rect 116596 139712 123390 139768
rect 123446 139712 123451 139768
rect 116596 139710 123451 139712
rect 116596 139708 116602 139710
rect 123385 139707 123451 139710
rect 164601 139770 164667 139773
rect 197486 139770 197492 139772
rect 164601 139768 197492 139770
rect 164601 139712 164606 139768
rect 164662 139712 197492 139768
rect 164601 139710 197492 139712
rect 164601 139707 164667 139710
rect 197486 139708 197492 139710
rect 197556 139708 197562 139772
rect 124489 139636 124555 139637
rect 124438 139634 124444 139636
rect 124398 139574 124444 139634
rect 124508 139632 124555 139636
rect 124550 139576 124555 139632
rect 124438 139572 124444 139574
rect 124508 139572 124555 139576
rect 125358 139572 125364 139636
rect 125428 139634 125434 139636
rect 125501 139634 125567 139637
rect 125428 139632 125567 139634
rect 125428 139576 125506 139632
rect 125562 139576 125567 139632
rect 125428 139574 125567 139576
rect 125428 139572 125434 139574
rect 124489 139571 124555 139572
rect 125501 139571 125567 139574
rect 127382 139572 127388 139636
rect 127452 139634 127458 139636
rect 127525 139634 127591 139637
rect 127452 139632 127591 139634
rect 127452 139576 127530 139632
rect 127586 139576 127591 139632
rect 127452 139574 127591 139576
rect 127452 139572 127458 139574
rect 127525 139571 127591 139574
rect 129457 139634 129523 139637
rect 188286 139634 188292 139636
rect 129457 139632 188292 139634
rect 129457 139576 129462 139632
rect 129518 139576 188292 139632
rect 129457 139574 188292 139576
rect 129457 139571 129523 139574
rect 188286 139572 188292 139574
rect 188356 139572 188362 139636
rect 8937 139498 9003 139501
rect 181253 139498 181319 139501
rect 187509 139498 187575 139501
rect 191782 139498 191788 139500
rect 8937 139496 181319 139498
rect 8937 139440 8942 139496
rect 8998 139440 181258 139496
rect 181314 139440 181319 139496
rect 8937 139438 181319 139440
rect 8937 139435 9003 139438
rect 181253 139435 181319 139438
rect 185350 139438 186514 139498
rect 111190 139300 111196 139364
rect 111260 139362 111266 139364
rect 115054 139362 115060 139364
rect 111260 139302 115060 139362
rect 111260 139300 111266 139302
rect 115054 139300 115060 139302
rect 115124 139300 115130 139364
rect 122966 139300 122972 139364
rect 123036 139362 123042 139364
rect 123109 139362 123175 139365
rect 123036 139360 123175 139362
rect 123036 139304 123114 139360
rect 123170 139304 123175 139360
rect 123036 139302 123175 139304
rect 123036 139300 123042 139302
rect 123109 139299 123175 139302
rect 123845 139362 123911 139365
rect 124070 139362 124076 139364
rect 123845 139360 124076 139362
rect 123845 139304 123850 139360
rect 123906 139304 124076 139360
rect 123845 139302 124076 139304
rect 123845 139299 123911 139302
rect 124070 139300 124076 139302
rect 124140 139300 124146 139364
rect 124254 139300 124260 139364
rect 124324 139362 124330 139364
rect 129181 139362 129247 139365
rect 131941 139362 132007 139365
rect 124324 139360 129247 139362
rect 124324 139304 129186 139360
rect 129242 139304 129247 139360
rect 124324 139302 129247 139304
rect 124324 139300 124330 139302
rect 129181 139299 129247 139302
rect 129414 139360 132007 139362
rect 129414 139304 131946 139360
rect 132002 139304 132007 139360
rect 129414 139302 132007 139304
rect 117998 139164 118004 139228
rect 118068 139226 118074 139228
rect 129414 139226 129474 139302
rect 131941 139299 132007 139302
rect 166717 139362 166783 139365
rect 173433 139362 173499 139365
rect 184105 139362 184171 139365
rect 184381 139362 184447 139365
rect 185350 139362 185410 139438
rect 166717 139360 167010 139362
rect 166717 139304 166722 139360
rect 166778 139304 167010 139360
rect 166717 139302 167010 139304
rect 166717 139299 166783 139302
rect 118068 139166 129474 139226
rect 118068 139164 118074 139166
rect 110873 139090 110939 139093
rect 124438 139090 124444 139092
rect 110873 139088 124444 139090
rect 110873 139032 110878 139088
rect 110934 139032 124444 139088
rect 110873 139030 124444 139032
rect 110873 139027 110939 139030
rect 124438 139028 124444 139030
rect 124508 139028 124514 139092
rect 114001 138954 114067 138957
rect 124254 138954 124260 138956
rect 114001 138952 124260 138954
rect 114001 138896 114006 138952
rect 114062 138896 124260 138952
rect 114001 138894 124260 138896
rect 114001 138891 114067 138894
rect 124254 138892 124260 138894
rect 124324 138892 124330 138956
rect 109534 138756 109540 138820
rect 109604 138818 109610 138820
rect 125358 138818 125364 138820
rect 109604 138758 125364 138818
rect 109604 138756 109610 138758
rect 125358 138756 125364 138758
rect 125428 138756 125434 138820
rect 112529 138682 112595 138685
rect 129038 138682 129044 138684
rect 112529 138680 129044 138682
rect 112529 138624 112534 138680
rect 112590 138624 129044 138680
rect 112529 138622 129044 138624
rect 112529 138619 112595 138622
rect 129038 138620 129044 138622
rect 129108 138620 129114 138684
rect 166950 138682 167010 139302
rect 173433 139360 180810 139362
rect 173433 139304 173438 139360
rect 173494 139304 180810 139360
rect 173433 139302 180810 139304
rect 173433 139299 173499 139302
rect 180750 138818 180810 139302
rect 184105 139360 184306 139362
rect 184105 139304 184110 139360
rect 184166 139304 184306 139360
rect 184105 139302 184306 139304
rect 184105 139299 184171 139302
rect 184246 138954 184306 139302
rect 184381 139360 185410 139362
rect 184381 139304 184386 139360
rect 184442 139304 185410 139360
rect 184381 139302 185410 139304
rect 185485 139362 185551 139365
rect 186221 139362 186287 139365
rect 186454 139362 186514 139438
rect 187509 139496 191788 139498
rect 187509 139440 187514 139496
rect 187570 139440 191788 139496
rect 187509 139438 191788 139440
rect 187509 139435 187575 139438
rect 191782 139436 191788 139438
rect 191852 139436 191858 139500
rect 193765 139362 193831 139365
rect 583520 139362 584960 139452
rect 185485 139360 185594 139362
rect 185485 139304 185490 139360
rect 185546 139304 185594 139360
rect 184381 139299 184447 139302
rect 185485 139299 185594 139304
rect 186221 139360 186330 139362
rect 186221 139304 186226 139360
rect 186282 139304 186330 139360
rect 186221 139299 186330 139304
rect 186454 139360 193831 139362
rect 186454 139304 193770 139360
rect 193826 139304 193831 139360
rect 186454 139302 193831 139304
rect 193765 139299 193831 139302
rect 583342 139302 584960 139362
rect 185534 139090 185594 139299
rect 186270 139226 186330 139299
rect 193673 139226 193739 139229
rect 186270 139224 193739 139226
rect 186270 139168 193678 139224
rect 193734 139168 193739 139224
rect 186270 139166 193739 139168
rect 583342 139226 583402 139302
rect 583520 139226 584960 139302
rect 583342 139212 584960 139226
rect 583342 139166 583586 139212
rect 193673 139163 193739 139166
rect 194041 139090 194107 139093
rect 185534 139088 194107 139090
rect 185534 139032 194046 139088
rect 194102 139032 194107 139088
rect 185534 139030 194107 139032
rect 194041 139027 194107 139030
rect 191281 138954 191347 138957
rect 184246 138952 191347 138954
rect 184246 138896 191286 138952
rect 191342 138896 191347 138952
rect 184246 138894 191347 138896
rect 191281 138891 191347 138894
rect 192477 138818 192543 138821
rect 180750 138816 192543 138818
rect 180750 138760 192482 138816
rect 192538 138760 192543 138816
rect 180750 138758 192543 138760
rect 192477 138755 192543 138758
rect 200849 138682 200915 138685
rect 166950 138680 200915 138682
rect 166950 138624 200854 138680
rect 200910 138624 200915 138680
rect 166950 138622 200915 138624
rect 200849 138619 200915 138622
rect 120993 138546 121059 138549
rect 121310 138546 121316 138548
rect 120993 138544 121316 138546
rect 120993 138488 120998 138544
rect 121054 138488 121316 138544
rect 120993 138486 121316 138488
rect 120993 138483 121059 138486
rect 121310 138484 121316 138486
rect 121380 138484 121386 138548
rect 114093 138410 114159 138413
rect 124806 138410 124812 138412
rect 114093 138408 124812 138410
rect 114093 138352 114098 138408
rect 114154 138352 124812 138408
rect 114093 138350 124812 138352
rect 114093 138347 114159 138350
rect 124806 138348 124812 138350
rect 124876 138348 124882 138412
rect 127382 138274 127388 138276
rect 118650 138214 127388 138274
rect 116669 138138 116735 138141
rect 118650 138138 118710 138214
rect 127382 138212 127388 138214
rect 127452 138212 127458 138276
rect 185342 138212 185348 138276
rect 185412 138274 185418 138276
rect 186630 138274 186636 138276
rect 185412 138214 186636 138274
rect 185412 138212 185418 138214
rect 186630 138212 186636 138214
rect 186700 138212 186706 138276
rect 116669 138136 118710 138138
rect 116669 138080 116674 138136
rect 116730 138080 118710 138136
rect 116669 138078 118710 138080
rect 121729 138138 121795 138141
rect 122782 138138 122788 138140
rect 121729 138136 122788 138138
rect 121729 138080 121734 138136
rect 121790 138080 122788 138136
rect 121729 138078 122788 138080
rect 116669 138075 116735 138078
rect 121729 138075 121795 138078
rect 122782 138076 122788 138078
rect 122852 138076 122858 138140
rect 185894 138076 185900 138140
rect 185964 138138 185970 138140
rect 186446 138138 186452 138140
rect 185964 138078 186452 138138
rect 185964 138076 185970 138078
rect 186446 138076 186452 138078
rect 186516 138076 186522 138140
rect 187049 138138 187115 138141
rect 187182 138138 187188 138140
rect 187049 138136 187188 138138
rect 187049 138080 187054 138136
rect 187110 138080 187188 138136
rect 187049 138078 187188 138080
rect 187049 138075 187115 138078
rect 187182 138076 187188 138078
rect 187252 138076 187258 138140
rect 188286 138076 188292 138140
rect 188356 138138 188362 138140
rect 583526 138138 583586 139166
rect 188356 138078 583586 138138
rect 188356 138076 188362 138078
rect 113766 137940 113772 138004
rect 113836 138002 113842 138004
rect 123886 138002 123892 138004
rect 113836 137942 123892 138002
rect 113836 137940 113842 137942
rect 123886 137940 123892 137942
rect 123956 137940 123962 138004
rect 184054 137940 184060 138004
rect 184124 138002 184130 138004
rect 187049 138002 187115 138005
rect 184124 138000 187115 138002
rect 184124 137944 187054 138000
rect 187110 137944 187115 138000
rect 184124 137942 187115 137944
rect 184124 137940 184130 137942
rect 187049 137939 187115 137942
rect 108113 137866 108179 137869
rect 126830 137866 126836 137868
rect 108113 137864 126836 137866
rect 108113 137808 108118 137864
rect 108174 137808 126836 137864
rect 108113 137806 126836 137808
rect 108113 137803 108179 137806
rect 126830 137804 126836 137806
rect 126900 137804 126906 137868
rect 185342 137804 185348 137868
rect 185412 137866 185418 137868
rect 187417 137866 187483 137869
rect 185412 137864 187483 137866
rect 185412 137808 187422 137864
rect 187478 137808 187483 137864
rect 185412 137806 187483 137808
rect 185412 137804 185418 137806
rect 187417 137803 187483 137806
rect 199326 137260 199332 137324
rect 199396 137322 199402 137324
rect 199745 137322 199811 137325
rect 199396 137320 199811 137322
rect 199396 137264 199750 137320
rect 199806 137264 199811 137320
rect 199396 137262 199811 137264
rect 199396 137260 199402 137262
rect 199745 137259 199811 137262
rect 187325 137186 187391 137189
rect 199561 137186 199627 137189
rect 187325 137184 199627 137186
rect 187325 137128 187330 137184
rect 187386 137128 199566 137184
rect 199622 137128 199627 137184
rect 187325 137126 199627 137128
rect 187325 137123 187391 137126
rect 199561 137123 199627 137126
rect -960 136778 480 136868
rect 3233 136778 3299 136781
rect -960 136776 3299 136778
rect -960 136720 3238 136776
rect 3294 136720 3299 136776
rect -960 136718 3299 136720
rect -960 136628 480 136718
rect 3233 136715 3299 136718
rect 119337 136642 119403 136645
rect 121821 136642 121887 136645
rect 119337 136640 121887 136642
rect 119337 136584 119342 136640
rect 119398 136584 121826 136640
rect 121882 136584 121887 136640
rect 119337 136582 121887 136584
rect 119337 136579 119403 136582
rect 121821 136579 121887 136582
rect 203558 136580 203564 136644
rect 203628 136642 203634 136644
rect 203701 136642 203767 136645
rect 203628 136640 203767 136642
rect 203628 136584 203706 136640
rect 203762 136584 203767 136640
rect 203628 136582 203767 136584
rect 203628 136580 203634 136582
rect 203701 136579 203767 136582
rect 186446 136036 186452 136100
rect 186516 136098 186522 136100
rect 201953 136098 202019 136101
rect 186516 136096 202019 136098
rect 186516 136040 201958 136096
rect 202014 136040 202019 136096
rect 186516 136038 202019 136040
rect 186516 136036 186522 136038
rect 201953 136035 202019 136038
rect 186630 135900 186636 135964
rect 186700 135962 186706 135964
rect 203701 135962 203767 135965
rect 186700 135960 203767 135962
rect 186700 135904 203706 135960
rect 203762 135904 203767 135960
rect 186700 135902 203767 135904
rect 186700 135900 186706 135902
rect 203701 135899 203767 135902
rect 121729 132562 121795 132565
rect 122782 132562 122788 132564
rect 121729 132560 122788 132562
rect 121729 132504 121734 132560
rect 121790 132504 122788 132560
rect 121729 132502 122788 132504
rect 121729 132499 121795 132502
rect 122782 132500 122788 132502
rect 122852 132500 122858 132564
rect 121821 132426 121887 132429
rect 122782 132426 122788 132428
rect 121821 132424 122788 132426
rect 121821 132368 121826 132424
rect 121882 132368 122788 132424
rect 121821 132366 122788 132368
rect 121821 132363 121887 132366
rect 122782 132364 122788 132366
rect 122852 132364 122858 132428
rect 580809 126034 580875 126037
rect 583520 126034 584960 126124
rect 580809 126032 584960 126034
rect 580809 125976 580814 126032
rect 580870 125976 584960 126032
rect 580809 125974 584960 125976
rect 580809 125971 580875 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 121821 122906 121887 122909
rect 122782 122906 122788 122908
rect 121821 122904 122788 122906
rect 121821 122848 121826 122904
rect 121882 122848 122788 122904
rect 121821 122846 122788 122848
rect 121821 122843 121887 122846
rect 122782 122844 122788 122846
rect 122852 122844 122858 122908
rect 121821 122770 121887 122773
rect 122782 122770 122788 122772
rect 121821 122768 122788 122770
rect 121821 122712 121826 122768
rect 121882 122712 122788 122768
rect 121821 122710 122788 122712
rect 121821 122707 121887 122710
rect 122782 122708 122788 122710
rect 122852 122708 122858 122772
rect 121821 113250 121887 113253
rect 122782 113250 122788 113252
rect 121821 113248 122788 113250
rect 121821 113192 121826 113248
rect 121882 113192 122788 113248
rect 121821 113190 122788 113192
rect 121821 113187 121887 113190
rect 122782 113188 122788 113190
rect 122852 113188 122858 113252
rect 121821 113114 121887 113117
rect 122782 113114 122788 113116
rect 121821 113112 122788 113114
rect 121821 113056 121826 113112
rect 121882 113056 122788 113112
rect 121821 113054 122788 113056
rect 121821 113051 121887 113054
rect 122782 113052 122788 113054
rect 122852 113052 122858 113116
rect 580625 112842 580691 112845
rect 583520 112842 584960 112932
rect 580625 112840 584960 112842
rect 580625 112784 580630 112840
rect 580686 112784 584960 112840
rect 580625 112782 584960 112784
rect 580625 112779 580691 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3049 110666 3115 110669
rect -960 110664 3115 110666
rect -960 110608 3054 110664
rect 3110 110608 3115 110664
rect -960 110606 3115 110608
rect -960 110516 480 110606
rect 3049 110603 3115 110606
rect 121821 103594 121887 103597
rect 122782 103594 122788 103596
rect 121821 103592 122788 103594
rect 121821 103536 121826 103592
rect 121882 103536 122788 103592
rect 121821 103534 122788 103536
rect 121821 103531 121887 103534
rect 122782 103532 122788 103534
rect 122852 103532 122858 103596
rect 121821 103458 121887 103461
rect 122782 103458 122788 103460
rect 121821 103456 122788 103458
rect 121821 103400 121826 103456
rect 121882 103400 122788 103456
rect 121821 103398 122788 103400
rect 121821 103395 121887 103398
rect 122782 103396 122788 103398
rect 122852 103396 122858 103460
rect 188337 100874 188403 100877
rect 189073 100874 189139 100877
rect 188337 100872 189139 100874
rect 188337 100816 188342 100872
rect 188398 100816 189078 100872
rect 189134 100816 189139 100872
rect 188337 100814 189139 100816
rect 188337 100811 188403 100814
rect 189073 100811 189139 100814
rect 187233 99514 187299 99517
rect 188613 99514 188679 99517
rect 187233 99512 188679 99514
rect 187233 99456 187238 99512
rect 187294 99456 188618 99512
rect 188674 99456 188679 99512
rect 187233 99454 188679 99456
rect 187233 99451 187299 99454
rect 188613 99451 188679 99454
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect 188337 98834 188403 98837
rect 188981 98834 189047 98837
rect 188337 98832 189047 98834
rect 188337 98776 188342 98832
rect 188398 98776 188986 98832
rect 189042 98776 189047 98832
rect 188337 98774 189047 98776
rect 188337 98771 188403 98774
rect 188981 98771 189047 98774
rect 187233 98698 187299 98701
rect 188245 98698 188311 98701
rect 187233 98696 188311 98698
rect 187233 98640 187238 98696
rect 187294 98640 188250 98696
rect 188306 98640 188311 98696
rect 187233 98638 188311 98640
rect 187233 98635 187299 98638
rect 188245 98635 188311 98638
rect -960 97610 480 97700
rect -960 97550 674 97610
rect -960 97474 480 97550
rect 614 97474 674 97550
rect -960 97460 674 97474
rect 246 97414 674 97460
rect 246 96930 306 97414
rect 246 96870 6930 96930
rect 6870 96658 6930 96870
rect 118734 96658 118740 96660
rect 6870 96598 118740 96658
rect 118734 96596 118740 96598
rect 118804 96596 118810 96660
rect 121821 93938 121887 93941
rect 122782 93938 122788 93940
rect 121821 93936 122788 93938
rect 121821 93880 121826 93936
rect 121882 93880 122788 93936
rect 121821 93878 122788 93880
rect 121821 93875 121887 93878
rect 122782 93876 122788 93878
rect 122852 93876 122858 93940
rect 186078 93740 186084 93804
rect 186148 93802 186154 93804
rect 188521 93802 188587 93805
rect 186148 93800 188587 93802
rect 186148 93744 188526 93800
rect 188582 93744 188587 93800
rect 186148 93742 188587 93744
rect 186148 93740 186154 93742
rect 188521 93739 188587 93742
rect 117773 92442 117839 92445
rect 122782 92442 122788 92444
rect 117773 92440 122788 92442
rect 117773 92384 117778 92440
rect 117834 92384 122788 92440
rect 117773 92382 122788 92384
rect 117773 92379 117839 92382
rect 122782 92380 122788 92382
rect 122852 92380 122858 92444
rect 186078 90340 186084 90404
rect 186148 90402 186154 90404
rect 195421 90402 195487 90405
rect 186148 90400 195487 90402
rect 186148 90344 195426 90400
rect 195482 90344 195487 90400
rect 186148 90342 195487 90344
rect 186148 90340 186154 90342
rect 195421 90339 195487 90342
rect 579981 86186 580047 86189
rect 583520 86186 584960 86276
rect 579981 86184 584960 86186
rect 579981 86128 579986 86184
rect 580042 86128 584960 86184
rect 579981 86126 584960 86128
rect 579981 86123 580047 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3509 84690 3575 84693
rect -960 84688 3575 84690
rect -960 84632 3514 84688
rect 3570 84632 3575 84688
rect -960 84630 3575 84632
rect -960 84540 480 84630
rect 3509 84627 3575 84630
rect 186078 84628 186084 84692
rect 186148 84690 186154 84692
rect 186814 84690 186820 84692
rect 186148 84630 186820 84690
rect 186148 84628 186154 84630
rect 186814 84628 186820 84630
rect 186884 84628 186890 84692
rect 186446 82044 186452 82108
rect 186516 82106 186522 82108
rect 196801 82106 196867 82109
rect 186516 82104 196867 82106
rect 186516 82048 196806 82104
rect 196862 82048 196867 82104
rect 186516 82046 196867 82048
rect 186516 82044 186522 82046
rect 196801 82043 196867 82046
rect 103973 81970 104039 81973
rect 125542 81970 125548 81972
rect 103973 81968 125548 81970
rect 103973 81912 103978 81968
rect 104034 81912 125548 81968
rect 103973 81910 125548 81912
rect 103973 81907 104039 81910
rect 125542 81908 125548 81910
rect 125612 81908 125618 81972
rect 203057 81970 203123 81973
rect 186086 81968 203123 81970
rect 186086 81912 203062 81968
rect 203118 81912 203123 81968
rect 186086 81910 203123 81912
rect 185710 81772 185716 81836
rect 185780 81834 185786 81836
rect 186086 81834 186146 81910
rect 203057 81907 203123 81910
rect 185780 81774 186146 81834
rect 185780 81772 185786 81774
rect 186262 81772 186268 81836
rect 186332 81834 186338 81836
rect 195329 81834 195395 81837
rect 186332 81832 195395 81834
rect 186332 81776 195334 81832
rect 195390 81776 195395 81832
rect 186332 81774 195395 81776
rect 186332 81772 186338 81774
rect 195329 81771 195395 81774
rect 184054 81636 184060 81700
rect 184124 81698 184130 81700
rect 193949 81698 194015 81701
rect 184124 81696 194015 81698
rect 184124 81640 193954 81696
rect 194010 81640 194015 81696
rect 184124 81638 194015 81640
rect 184124 81636 184130 81638
rect 193949 81635 194015 81638
rect 181294 81500 181300 81564
rect 181364 81562 181370 81564
rect 186262 81562 186268 81564
rect 181364 81502 186268 81562
rect 181364 81500 181370 81502
rect 186262 81500 186268 81502
rect 186332 81500 186338 81564
rect 201217 81428 201283 81429
rect 185342 81364 185348 81428
rect 185412 81426 185418 81428
rect 186814 81426 186820 81428
rect 185412 81366 186820 81426
rect 185412 81364 185418 81366
rect 186814 81364 186820 81366
rect 186884 81364 186890 81428
rect 201166 81426 201172 81428
rect 201126 81366 201172 81426
rect 201236 81424 201283 81428
rect 201278 81368 201283 81424
rect 201166 81364 201172 81366
rect 201236 81364 201283 81368
rect 201217 81363 201283 81364
rect 176326 81228 176332 81292
rect 176396 81290 176402 81292
rect 197670 81290 197676 81292
rect 176396 81230 197676 81290
rect 176396 81228 176402 81230
rect 197670 81228 197676 81230
rect 197740 81228 197746 81292
rect 117865 81154 117931 81157
rect 129222 81154 129228 81156
rect 117865 81152 129228 81154
rect 117865 81096 117870 81152
rect 117926 81096 129228 81152
rect 117865 81094 129228 81096
rect 117865 81091 117931 81094
rect 129222 81092 129228 81094
rect 129292 81092 129298 81156
rect 170438 81092 170444 81156
rect 170508 81154 170514 81156
rect 192150 81154 192156 81156
rect 170508 81094 192156 81154
rect 170508 81092 170514 81094
rect 192150 81092 192156 81094
rect 192220 81092 192226 81156
rect 122373 81018 122439 81021
rect 146886 81018 146892 81020
rect 122373 81016 146892 81018
rect 122373 80960 122378 81016
rect 122434 80960 146892 81016
rect 122373 80958 146892 80960
rect 122373 80955 122439 80958
rect 146886 80956 146892 80958
rect 146956 80956 146962 81020
rect 174670 80956 174676 81020
rect 174740 81018 174746 81020
rect 199142 81018 199148 81020
rect 174740 80958 199148 81018
rect 174740 80956 174746 80958
rect 199142 80956 199148 80958
rect 199212 80956 199218 81020
rect 116393 80882 116459 80885
rect 149830 80882 149836 80884
rect 116393 80880 149836 80882
rect 116393 80824 116398 80880
rect 116454 80824 149836 80880
rect 116393 80822 149836 80824
rect 116393 80819 116459 80822
rect 149830 80820 149836 80822
rect 149900 80820 149906 80884
rect 196198 80882 196204 80884
rect 179370 80822 196204 80882
rect 121126 80684 121132 80748
rect 121196 80746 121202 80748
rect 121196 80686 138030 80746
rect 121196 80684 121202 80686
rect 129222 80548 129228 80612
rect 129292 80610 129298 80612
rect 130009 80610 130075 80613
rect 129292 80608 130075 80610
rect 129292 80552 130014 80608
rect 130070 80552 130075 80608
rect 129292 80550 130075 80552
rect 129292 80548 129298 80550
rect 130009 80547 130075 80550
rect 137970 80338 138030 80686
rect 170622 80684 170628 80748
rect 170692 80746 170698 80748
rect 179370 80746 179430 80822
rect 196198 80820 196204 80822
rect 196268 80820 196274 80884
rect 211521 80746 211587 80749
rect 523125 80746 523191 80749
rect 170692 80686 179430 80746
rect 180750 80744 523191 80746
rect 180750 80688 211526 80744
rect 211582 80688 523130 80744
rect 523186 80688 523191 80744
rect 180750 80686 523191 80688
rect 170692 80684 170698 80686
rect 178033 80610 178099 80613
rect 180750 80610 180810 80686
rect 211521 80683 211587 80686
rect 523125 80683 523191 80686
rect 178033 80608 180810 80610
rect 178033 80552 178038 80608
rect 178094 80552 180810 80608
rect 178033 80550 180810 80552
rect 178033 80547 178099 80550
rect 137970 80278 151508 80338
rect 129733 80202 129799 80205
rect 151302 80202 151308 80204
rect 129733 80200 140882 80202
rect 129733 80144 129738 80200
rect 129794 80144 140882 80200
rect 129733 80142 140882 80144
rect 129733 80139 129799 80142
rect 132450 80006 132924 80066
rect 128537 79930 128603 79933
rect 132450 79930 132510 80006
rect 132631 79930 132697 79933
rect 128537 79928 132510 79930
rect 128537 79872 128542 79928
rect 128598 79872 132510 79928
rect 128537 79870 132510 79872
rect 132588 79928 132697 79930
rect 132588 79872 132636 79928
rect 132692 79872 132697 79928
rect 128537 79867 128603 79870
rect 132588 79867 132697 79872
rect 132588 79522 132648 79867
rect 132864 79797 132924 80006
rect 140822 79967 140882 80142
rect 141558 80142 145298 80202
rect 133183 79964 133249 79967
rect 133551 79964 133617 79967
rect 134195 79964 134261 79967
rect 133183 79962 133384 79964
rect 133183 79930 133188 79962
rect 133094 79906 133188 79930
rect 133244 79906 133384 79962
rect 133094 79870 133384 79906
rect 133551 79962 133752 79964
rect 133551 79906 133556 79962
rect 133612 79906 133752 79962
rect 134060 79962 134261 79964
rect 134060 79932 134200 79962
rect 133551 79904 133752 79906
rect 133551 79901 133617 79904
rect 132861 79792 132927 79797
rect 132861 79736 132866 79792
rect 132922 79736 132927 79792
rect 132861 79731 132927 79736
rect 133094 79661 133154 79870
rect 133229 79794 133295 79797
rect 133413 79794 133479 79797
rect 133692 79794 133752 79904
rect 134006 79868 134012 79932
rect 134076 79906 134200 79932
rect 134256 79906 134261 79962
rect 134076 79904 134261 79906
rect 134076 79870 134120 79904
rect 134195 79901 134261 79904
rect 134931 79962 134997 79967
rect 134931 79906 134936 79962
rect 134992 79906 134997 79962
rect 135667 79962 135733 79967
rect 135943 79964 136009 79967
rect 134931 79901 134997 79906
rect 135299 79930 135365 79933
rect 135478 79930 135484 79932
rect 135299 79928 135484 79930
rect 134747 79894 134813 79899
rect 134076 79868 134082 79870
rect 134747 79838 134752 79894
rect 134808 79838 134813 79894
rect 134747 79833 134813 79838
rect 133229 79792 133338 79794
rect 133229 79736 133234 79792
rect 133290 79736 133338 79792
rect 133229 79731 133338 79736
rect 133413 79792 133752 79794
rect 133413 79736 133418 79792
rect 133474 79736 133752 79792
rect 133413 79734 133752 79736
rect 133413 79731 133479 79734
rect 133278 79661 133338 79731
rect 133045 79656 133154 79661
rect 133045 79600 133050 79656
rect 133106 79600 133154 79656
rect 133045 79598 133154 79600
rect 133229 79656 133338 79661
rect 133229 79600 133234 79656
rect 133290 79600 133338 79656
rect 133229 79598 133338 79600
rect 133045 79595 133111 79598
rect 133229 79595 133295 79598
rect 133822 79596 133828 79660
rect 133892 79658 133898 79660
rect 134750 79658 134810 79833
rect 133892 79598 134810 79658
rect 134934 79661 134994 79901
rect 135299 79872 135304 79928
rect 135360 79872 135484 79928
rect 135299 79870 135484 79872
rect 135299 79867 135365 79870
rect 135478 79868 135484 79870
rect 135548 79868 135554 79932
rect 135667 79906 135672 79962
rect 135728 79906 135733 79962
rect 135667 79901 135733 79906
rect 135808 79962 136009 79964
rect 135808 79906 135948 79962
rect 136004 79906 136009 79962
rect 135808 79904 136009 79906
rect 134934 79656 135043 79661
rect 134934 79600 134982 79656
rect 135038 79600 135043 79656
rect 134934 79598 135043 79600
rect 133892 79596 133898 79598
rect 134977 79595 135043 79598
rect 133454 79522 133460 79524
rect 132588 79462 133460 79522
rect 133454 79460 133460 79462
rect 133524 79460 133530 79524
rect 135529 79522 135595 79525
rect 135670 79522 135730 79901
rect 135808 79794 135868 79904
rect 135943 79901 136009 79904
rect 136495 79962 136561 79967
rect 136495 79906 136500 79962
rect 136556 79906 136561 79962
rect 137323 79962 137389 79967
rect 137047 79930 137113 79933
rect 136495 79901 136561 79906
rect 137004 79928 137113 79930
rect 135989 79794 136055 79797
rect 135808 79792 136055 79794
rect 135808 79736 135994 79792
rect 136050 79736 136055 79792
rect 135808 79734 136055 79736
rect 135989 79731 136055 79734
rect 136498 79661 136558 79901
rect 137004 79872 137052 79928
rect 137108 79872 137113 79928
rect 137323 79906 137328 79962
rect 137384 79930 137389 79962
rect 138979 79962 139045 79967
rect 137686 79930 137692 79932
rect 137384 79906 137692 79930
rect 137323 79901 137692 79906
rect 137004 79867 137113 79872
rect 137326 79870 137692 79901
rect 137686 79868 137692 79870
rect 137756 79868 137762 79932
rect 137875 79894 137941 79899
rect 137004 79797 137064 79867
rect 137875 79838 137880 79894
rect 137936 79838 137941 79894
rect 138054 79868 138060 79932
rect 138124 79930 138130 79932
rect 138519 79930 138585 79933
rect 138979 79932 138984 79962
rect 139040 79932 139045 79962
rect 139715 79962 139781 79967
rect 138124 79928 138585 79930
rect 138124 79872 138524 79928
rect 138580 79872 138585 79928
rect 138124 79870 138585 79872
rect 138124 79868 138130 79870
rect 138519 79867 138585 79870
rect 138974 79868 138980 79932
rect 139044 79930 139050 79932
rect 139439 79930 139505 79933
rect 139715 79932 139720 79962
rect 139776 79932 139781 79962
rect 140267 79962 140333 79967
rect 139044 79870 139102 79930
rect 139439 79928 139640 79930
rect 139163 79894 139229 79899
rect 139044 79868 139050 79870
rect 137875 79833 137941 79838
rect 139163 79838 139168 79894
rect 139224 79838 139229 79894
rect 139439 79872 139444 79928
rect 139500 79872 139640 79928
rect 139439 79870 139640 79872
rect 139439 79867 139505 79870
rect 139163 79833 139229 79838
rect 137001 79792 137067 79797
rect 137691 79794 137757 79797
rect 137001 79736 137006 79792
rect 137062 79736 137067 79792
rect 137001 79731 137067 79736
rect 137142 79792 137757 79794
rect 137142 79736 137696 79792
rect 137752 79736 137757 79792
rect 137142 79734 137757 79736
rect 136449 79656 136558 79661
rect 136449 79600 136454 79656
rect 136510 79600 136558 79656
rect 136449 79598 136558 79600
rect 136909 79658 136975 79661
rect 136909 79656 137018 79658
rect 136909 79600 136914 79656
rect 136970 79600 137018 79656
rect 136449 79595 136515 79598
rect 136909 79595 137018 79600
rect 135529 79520 135730 79522
rect 135529 79464 135534 79520
rect 135590 79464 135730 79520
rect 135529 79462 135730 79464
rect 136265 79522 136331 79525
rect 136958 79522 137018 79595
rect 136265 79520 137018 79522
rect 136265 79464 136270 79520
rect 136326 79464 137018 79520
rect 136265 79462 137018 79464
rect 137142 79522 137202 79734
rect 137691 79731 137757 79734
rect 137277 79658 137343 79661
rect 137878 79658 137938 79833
rect 138335 79794 138401 79797
rect 137277 79656 137938 79658
rect 137277 79600 137282 79656
rect 137338 79600 137938 79656
rect 137277 79598 137938 79600
rect 138062 79792 138401 79794
rect 138062 79736 138340 79792
rect 138396 79736 138401 79792
rect 138062 79734 138401 79736
rect 138062 79658 138122 79734
rect 138335 79731 138401 79734
rect 138565 79796 138631 79797
rect 138565 79792 138612 79796
rect 138676 79794 138682 79796
rect 138565 79736 138570 79792
rect 138565 79732 138612 79736
rect 138676 79734 138722 79794
rect 138676 79732 138682 79734
rect 138565 79731 138631 79732
rect 139166 79661 139226 79833
rect 139580 79794 139640 79870
rect 139710 79868 139716 79932
rect 139780 79930 139786 79932
rect 139780 79870 139838 79930
rect 139780 79868 139786 79870
rect 140078 79868 140084 79932
rect 140148 79930 140154 79932
rect 140267 79930 140272 79962
rect 140148 79906 140272 79930
rect 140328 79906 140333 79962
rect 140148 79901 140333 79906
rect 140819 79962 140885 79967
rect 140819 79906 140824 79962
rect 140880 79906 140885 79962
rect 140819 79901 140885 79906
rect 140148 79870 140330 79901
rect 140148 79868 140154 79870
rect 140998 79868 141004 79932
rect 141068 79930 141074 79932
rect 141371 79930 141437 79933
rect 141068 79928 141437 79930
rect 141068 79872 141376 79928
rect 141432 79872 141437 79928
rect 141068 79870 141437 79872
rect 141068 79868 141074 79870
rect 141371 79867 141437 79870
rect 139894 79794 139900 79796
rect 139580 79734 139900 79794
rect 139894 79732 139900 79734
rect 139964 79732 139970 79796
rect 141558 79794 141618 80142
rect 143390 80004 143396 80068
rect 143460 80066 143466 80068
rect 143460 80006 144194 80066
rect 143460 80004 143466 80006
rect 142659 79932 142725 79933
rect 143579 79932 143645 79933
rect 142654 79930 142660 79932
rect 142291 79894 142357 79899
rect 142291 79838 142296 79894
rect 142352 79838 142357 79894
rect 142568 79870 142660 79930
rect 142654 79868 142660 79870
rect 142724 79868 142730 79932
rect 143574 79930 143580 79932
rect 143211 79894 143277 79899
rect 142659 79867 142725 79868
rect 142291 79833 142357 79838
rect 143211 79838 143216 79894
rect 143272 79838 143277 79894
rect 143488 79870 143580 79930
rect 143574 79868 143580 79870
rect 143644 79868 143650 79932
rect 144134 79930 144194 80006
rect 145238 79967 145298 80142
rect 150574 80142 151308 80202
rect 150574 79967 150634 80142
rect 151302 80140 151308 80142
rect 151372 80140 151378 80204
rect 151448 80066 151508 80278
rect 173198 80276 173204 80340
rect 173268 80338 173274 80340
rect 178309 80338 178375 80341
rect 173268 80336 178375 80338
rect 173268 80280 178314 80336
rect 178370 80280 178375 80336
rect 173268 80278 178375 80280
rect 173268 80276 173274 80278
rect 178309 80275 178375 80278
rect 183461 80338 183527 80341
rect 189022 80338 189028 80340
rect 183461 80336 189028 80338
rect 183461 80280 183466 80336
rect 183522 80280 189028 80336
rect 183461 80278 189028 80280
rect 183461 80275 183527 80278
rect 189022 80276 189028 80278
rect 189092 80276 189098 80340
rect 187734 80202 187740 80204
rect 154806 80142 160570 80202
rect 151448 80006 154084 80066
rect 154024 79967 154084 80006
rect 145051 79962 145117 79967
rect 144134 79870 144746 79930
rect 145051 79906 145056 79962
rect 145112 79906 145117 79962
rect 145051 79901 145117 79906
rect 145235 79962 145301 79967
rect 145235 79906 145240 79962
rect 145296 79906 145301 79962
rect 145971 79962 146037 79967
rect 145235 79901 145301 79906
rect 143579 79867 143645 79868
rect 143211 79833 143277 79838
rect 140086 79734 141618 79794
rect 138238 79658 138244 79660
rect 138062 79598 138244 79658
rect 137277 79595 137343 79598
rect 138238 79596 138244 79598
rect 138308 79596 138314 79660
rect 139166 79656 139275 79661
rect 139166 79600 139214 79656
rect 139270 79600 139275 79656
rect 139166 79598 139275 79600
rect 139209 79595 139275 79598
rect 139669 79658 139735 79661
rect 140086 79658 140146 79734
rect 139669 79656 140146 79658
rect 139669 79600 139674 79656
rect 139730 79600 140146 79656
rect 139669 79598 140146 79600
rect 140221 79658 140287 79661
rect 142294 79658 142354 79833
rect 140221 79656 142354 79658
rect 140221 79600 140226 79656
rect 140282 79600 142354 79656
rect 140221 79598 142354 79600
rect 143214 79658 143274 79833
rect 143763 79826 143829 79831
rect 143763 79794 143768 79826
rect 143582 79770 143768 79794
rect 143824 79770 143829 79826
rect 143582 79765 143829 79770
rect 143947 79792 144013 79797
rect 143582 79734 143826 79765
rect 143947 79736 143952 79792
rect 144008 79736 144013 79792
rect 143441 79658 143507 79661
rect 143214 79656 143507 79658
rect 143214 79600 143446 79656
rect 143502 79600 143507 79656
rect 143214 79598 143507 79600
rect 139669 79595 139735 79598
rect 140221 79595 140287 79598
rect 143441 79595 143507 79598
rect 137553 79522 137619 79525
rect 137142 79520 137619 79522
rect 137142 79464 137558 79520
rect 137614 79464 137619 79520
rect 137142 79462 137619 79464
rect 135529 79459 135595 79462
rect 136265 79459 136331 79462
rect 137553 79459 137619 79462
rect 139485 79386 139551 79389
rect 142245 79386 142311 79389
rect 139485 79384 142311 79386
rect 139485 79328 139490 79384
rect 139546 79328 142250 79384
rect 142306 79328 142311 79384
rect 139485 79326 142311 79328
rect 143582 79386 143642 79734
rect 143947 79731 144013 79736
rect 144686 79794 144746 79870
rect 144821 79794 144887 79797
rect 144686 79792 144887 79794
rect 144686 79736 144826 79792
rect 144882 79736 144887 79792
rect 144686 79734 144887 79736
rect 144821 79731 144887 79734
rect 143950 79522 144010 79731
rect 144269 79660 144335 79661
rect 144269 79656 144316 79660
rect 144380 79658 144386 79660
rect 144545 79658 144611 79661
rect 144269 79600 144274 79656
rect 144269 79596 144316 79600
rect 144380 79598 144426 79658
rect 144545 79656 144792 79658
rect 144545 79600 144550 79656
rect 144606 79600 144792 79656
rect 144545 79598 144792 79600
rect 144380 79596 144386 79598
rect 144269 79595 144335 79596
rect 144545 79595 144611 79598
rect 144732 79525 144792 79598
rect 145054 79525 145114 79901
rect 145598 79868 145604 79932
rect 145668 79930 145674 79932
rect 145971 79930 145976 79962
rect 145668 79906 145976 79930
rect 146032 79906 146037 79962
rect 145668 79901 146037 79906
rect 146155 79962 146221 79967
rect 146155 79906 146160 79962
rect 146216 79906 146221 79962
rect 146707 79962 146773 79967
rect 146707 79930 146712 79962
rect 146155 79901 146221 79906
rect 146388 79906 146712 79930
rect 146768 79906 146773 79962
rect 147811 79962 147877 79967
rect 146388 79901 146773 79906
rect 145668 79870 146034 79901
rect 145668 79868 145674 79870
rect 145925 79794 145991 79797
rect 145606 79792 145991 79794
rect 145606 79736 145930 79792
rect 145986 79736 145991 79792
rect 145606 79734 145991 79736
rect 144545 79522 144611 79525
rect 143950 79520 144611 79522
rect 143950 79464 144550 79520
rect 144606 79464 144611 79520
rect 143950 79462 144611 79464
rect 144545 79459 144611 79462
rect 144729 79520 144795 79525
rect 144729 79464 144734 79520
rect 144790 79464 144795 79520
rect 144729 79459 144795 79464
rect 145054 79520 145163 79525
rect 145054 79464 145102 79520
rect 145158 79464 145163 79520
rect 145054 79462 145163 79464
rect 145097 79459 145163 79462
rect 145414 79460 145420 79524
rect 145484 79522 145490 79524
rect 145606 79522 145666 79734
rect 145925 79731 145991 79734
rect 146158 79525 146218 79901
rect 146388 79870 146770 79901
rect 146388 79658 146448 79870
rect 147070 79868 147076 79932
rect 147140 79930 147146 79932
rect 147259 79930 147325 79933
rect 147811 79932 147816 79962
rect 147872 79932 147877 79962
rect 148179 79962 148245 79967
rect 148179 79932 148184 79962
rect 148240 79932 148245 79962
rect 148731 79962 148797 79967
rect 147140 79928 147325 79930
rect 147140 79872 147264 79928
rect 147320 79872 147325 79928
rect 147140 79870 147325 79872
rect 147140 79868 147146 79870
rect 147259 79867 147325 79870
rect 147806 79868 147812 79932
rect 147876 79930 147882 79932
rect 147876 79870 147934 79930
rect 147876 79868 147882 79870
rect 148174 79868 148180 79932
rect 148244 79930 148250 79932
rect 148244 79870 148302 79930
rect 148547 79928 148613 79933
rect 148547 79872 148552 79928
rect 148608 79872 148613 79928
rect 148731 79906 148736 79962
rect 148792 79906 148797 79962
rect 150571 79962 150637 79967
rect 148731 79901 148797 79906
rect 149191 79930 149257 79933
rect 149830 79930 149836 79932
rect 149191 79928 149836 79930
rect 148244 79868 148250 79870
rect 148547 79867 148613 79872
rect 146518 79732 146524 79796
rect 146588 79794 146594 79796
rect 147627 79794 147693 79797
rect 148550 79794 148610 79867
rect 146588 79792 147693 79794
rect 146588 79736 147632 79792
rect 147688 79736 147693 79792
rect 146588 79734 147693 79736
rect 146588 79732 146594 79734
rect 147627 79731 147693 79734
rect 147814 79734 148610 79794
rect 146661 79658 146727 79661
rect 146388 79656 146727 79658
rect 146388 79600 146666 79656
rect 146722 79600 146727 79656
rect 146388 79598 146727 79600
rect 146661 79595 146727 79598
rect 146886 79596 146892 79660
rect 146956 79658 146962 79660
rect 147213 79658 147279 79661
rect 146956 79656 147279 79658
rect 146956 79600 147218 79656
rect 147274 79600 147279 79656
rect 146956 79598 147279 79600
rect 146956 79596 146962 79598
rect 147213 79595 147279 79598
rect 147673 79658 147739 79661
rect 147814 79658 147874 79734
rect 147673 79656 147874 79658
rect 147673 79600 147678 79656
rect 147734 79600 147874 79656
rect 147673 79598 147874 79600
rect 148409 79658 148475 79661
rect 148734 79658 148794 79901
rect 149191 79872 149196 79928
rect 149252 79872 149836 79928
rect 149191 79870 149836 79872
rect 149191 79867 149257 79870
rect 149830 79868 149836 79870
rect 149900 79868 149906 79932
rect 150571 79906 150576 79962
rect 150632 79906 150637 79962
rect 154024 79962 154133 79967
rect 150571 79901 150637 79906
rect 152687 79930 152753 79933
rect 153878 79930 153884 79932
rect 152687 79928 153884 79930
rect 150755 79894 150821 79899
rect 150755 79838 150760 79894
rect 150816 79838 150821 79894
rect 152687 79872 152692 79928
rect 152748 79872 153884 79928
rect 152687 79870 153884 79872
rect 152687 79867 152753 79870
rect 153878 79868 153884 79870
rect 153948 79868 153954 79932
rect 154024 79906 154072 79962
rect 154128 79906 154133 79962
rect 154024 79904 154133 79906
rect 154067 79901 154133 79904
rect 154435 79962 154501 79967
rect 154435 79906 154440 79962
rect 154496 79906 154501 79962
rect 154435 79901 154501 79906
rect 150755 79833 150821 79838
rect 148409 79656 148794 79658
rect 148409 79600 148414 79656
rect 148470 79600 148794 79656
rect 148409 79598 148794 79600
rect 150065 79658 150131 79661
rect 150249 79658 150315 79661
rect 150065 79656 150315 79658
rect 150065 79600 150070 79656
rect 150126 79600 150254 79656
rect 150310 79600 150315 79656
rect 150065 79598 150315 79600
rect 150758 79658 150818 79833
rect 151859 79794 151925 79797
rect 152273 79794 152339 79797
rect 151859 79792 152339 79794
rect 151859 79736 151864 79792
rect 151920 79736 152278 79792
rect 152334 79736 152339 79792
rect 151859 79734 152339 79736
rect 151859 79731 151925 79734
rect 152273 79731 152339 79734
rect 152595 79794 152661 79797
rect 152774 79794 152780 79796
rect 152595 79792 152780 79794
rect 152595 79736 152600 79792
rect 152656 79736 152780 79792
rect 152595 79734 152780 79736
rect 152595 79731 152661 79734
rect 152774 79732 152780 79734
rect 152844 79732 152850 79796
rect 153285 79792 153351 79797
rect 154297 79794 154363 79797
rect 153285 79736 153290 79792
rect 153346 79736 153351 79792
rect 153285 79731 153351 79736
rect 154254 79792 154363 79794
rect 154254 79736 154302 79792
rect 154358 79736 154363 79792
rect 154254 79731 154363 79736
rect 151261 79658 151327 79661
rect 150758 79656 151327 79658
rect 150758 79600 151266 79656
rect 151322 79600 151327 79656
rect 150758 79598 151327 79600
rect 147673 79595 147739 79598
rect 148409 79595 148475 79598
rect 150065 79595 150131 79598
rect 150249 79595 150315 79598
rect 151261 79595 151327 79598
rect 151445 79658 151511 79661
rect 153288 79658 153348 79731
rect 153469 79658 153535 79661
rect 151445 79656 151554 79658
rect 151445 79600 151450 79656
rect 151506 79600 151554 79656
rect 151445 79595 151554 79600
rect 153288 79656 153535 79658
rect 153288 79600 153474 79656
rect 153530 79600 153535 79656
rect 153288 79598 153535 79600
rect 153469 79595 153535 79598
rect 153653 79658 153719 79661
rect 153837 79658 153903 79661
rect 153653 79656 153903 79658
rect 153653 79600 153658 79656
rect 153714 79600 153842 79656
rect 153898 79600 153903 79656
rect 153653 79598 153903 79600
rect 153653 79595 153719 79598
rect 153837 79595 153903 79598
rect 145484 79462 145666 79522
rect 146109 79520 146218 79525
rect 146109 79464 146114 79520
rect 146170 79464 146218 79520
rect 146109 79462 146218 79464
rect 147857 79522 147923 79525
rect 148685 79522 148751 79525
rect 147857 79520 148751 79522
rect 147857 79464 147862 79520
rect 147918 79464 148690 79520
rect 148746 79464 148751 79520
rect 147857 79462 148751 79464
rect 145484 79460 145490 79462
rect 146109 79459 146175 79462
rect 147857 79459 147923 79462
rect 148685 79459 148751 79462
rect 150801 79522 150867 79525
rect 151494 79522 151554 79595
rect 154254 79525 154314 79731
rect 154438 79661 154498 79901
rect 154806 79831 154866 80142
rect 154987 79962 155053 79967
rect 154987 79932 154992 79962
rect 155048 79932 155053 79962
rect 155263 79962 155329 79967
rect 154982 79868 154988 79932
rect 155052 79930 155058 79932
rect 155052 79870 155110 79930
rect 155263 79906 155268 79962
rect 155324 79906 155329 79962
rect 155907 79964 155973 79967
rect 155907 79962 156030 79964
rect 155263 79901 155329 79906
rect 155539 79930 155605 79933
rect 155907 79932 155912 79962
rect 155968 79932 156030 79962
rect 155539 79928 155786 79930
rect 155052 79868 155058 79870
rect 154803 79826 154869 79831
rect 154803 79770 154808 79826
rect 154864 79770 154869 79826
rect 154803 79765 154869 79770
rect 155266 79794 155326 79901
rect 155539 79872 155544 79928
rect 155600 79872 155786 79928
rect 155539 79870 155786 79872
rect 155539 79867 155605 79870
rect 155534 79794 155540 79796
rect 155266 79734 155540 79794
rect 155534 79732 155540 79734
rect 155604 79732 155610 79796
rect 155726 79661 155786 79870
rect 155902 79868 155908 79932
rect 155972 79904 156030 79932
rect 156091 79962 156157 79967
rect 156091 79906 156096 79962
rect 156152 79906 156157 79962
rect 155972 79868 155978 79904
rect 156091 79901 156157 79906
rect 156275 79962 156341 79967
rect 156275 79906 156280 79962
rect 156336 79906 156341 79962
rect 156275 79901 156341 79906
rect 156735 79964 156801 79967
rect 157471 79964 157537 79967
rect 156735 79962 156844 79964
rect 156735 79906 156740 79962
rect 156796 79906 156844 79962
rect 157471 79962 157810 79964
rect 156735 79901 156844 79906
rect 154389 79656 154498 79661
rect 154389 79600 154394 79656
rect 154450 79600 154498 79656
rect 154389 79598 154498 79600
rect 155677 79656 155786 79661
rect 155677 79600 155682 79656
rect 155738 79600 155786 79656
rect 155677 79598 155786 79600
rect 154389 79595 154455 79598
rect 155677 79595 155743 79598
rect 150801 79520 151554 79522
rect 150801 79464 150806 79520
rect 150862 79464 151554 79520
rect 150801 79462 151554 79464
rect 154205 79520 154314 79525
rect 154205 79464 154210 79520
rect 154266 79464 154314 79520
rect 154205 79462 154314 79464
rect 156094 79522 156154 79901
rect 156278 79658 156338 79901
rect 156784 79794 156844 79901
rect 157287 79928 157353 79933
rect 157287 79872 157292 79928
rect 157348 79872 157353 79928
rect 157471 79906 157476 79962
rect 157532 79906 157810 79962
rect 158575 79962 158641 79967
rect 159311 79964 159377 79967
rect 157471 79904 157810 79906
rect 157471 79901 157537 79904
rect 157287 79867 157353 79872
rect 156646 79734 156844 79794
rect 156646 79661 156706 79734
rect 156413 79658 156479 79661
rect 156278 79656 156479 79658
rect 156278 79600 156418 79656
rect 156474 79600 156479 79656
rect 156278 79598 156479 79600
rect 156646 79656 156755 79661
rect 156646 79600 156694 79656
rect 156750 79600 156755 79656
rect 156646 79598 156755 79600
rect 156413 79595 156479 79598
rect 156689 79595 156755 79598
rect 156873 79658 156939 79661
rect 157290 79658 157350 79867
rect 156873 79656 157350 79658
rect 156873 79600 156878 79656
rect 156934 79600 157350 79656
rect 156873 79598 157350 79600
rect 157750 79658 157810 79904
rect 157926 79868 157932 79932
rect 157996 79930 158002 79932
rect 158115 79930 158181 79933
rect 158575 79930 158580 79962
rect 157996 79928 158181 79930
rect 157996 79872 158120 79928
rect 158176 79872 158181 79928
rect 157996 79870 158181 79872
rect 157996 79868 158002 79870
rect 158115 79867 158181 79870
rect 158440 79906 158580 79930
rect 158636 79906 158641 79962
rect 158440 79901 158641 79906
rect 159038 79962 159377 79964
rect 159038 79906 159316 79962
rect 159372 79906 159377 79962
rect 159038 79904 159377 79906
rect 158440 79870 158638 79901
rect 158440 79796 158500 79870
rect 158440 79734 158484 79796
rect 158478 79732 158484 79734
rect 158548 79732 158554 79796
rect 158897 79794 158963 79797
rect 158670 79792 158963 79794
rect 158670 79736 158902 79792
rect 158958 79736 158963 79792
rect 158670 79734 158963 79736
rect 158437 79658 158503 79661
rect 157750 79656 158503 79658
rect 157750 79600 158442 79656
rect 158498 79600 158503 79656
rect 157750 79598 158503 79600
rect 156873 79595 156939 79598
rect 158437 79595 158503 79598
rect 156321 79522 156387 79525
rect 156094 79520 156387 79522
rect 156094 79464 156326 79520
rect 156382 79464 156387 79520
rect 156094 79462 156387 79464
rect 150801 79459 150867 79462
rect 154205 79459 154271 79462
rect 156321 79459 156387 79462
rect 144361 79386 144427 79389
rect 147857 79388 147923 79389
rect 143582 79384 144427 79386
rect 143582 79328 144366 79384
rect 144422 79328 144427 79384
rect 143582 79326 144427 79328
rect 139485 79323 139551 79326
rect 142245 79323 142311 79326
rect 144361 79323 144427 79326
rect 147806 79324 147812 79388
rect 147876 79386 147923 79388
rect 148133 79388 148199 79389
rect 148133 79386 148180 79388
rect 147876 79384 147968 79386
rect 147918 79328 147968 79384
rect 147876 79326 147968 79328
rect 148088 79384 148180 79386
rect 148088 79328 148138 79384
rect 148088 79326 148180 79328
rect 147876 79324 147923 79326
rect 147857 79323 147923 79324
rect 148133 79324 148180 79326
rect 148244 79324 148250 79388
rect 153929 79386 153995 79389
rect 154430 79386 154436 79388
rect 153929 79384 154436 79386
rect 153929 79328 153934 79384
rect 153990 79328 154436 79384
rect 153929 79326 154436 79328
rect 148133 79323 148199 79324
rect 153929 79323 153995 79326
rect 154430 79324 154436 79326
rect 154500 79324 154506 79388
rect 119654 79188 119660 79252
rect 119724 79250 119730 79252
rect 153285 79250 153351 79253
rect 119724 79248 153351 79250
rect 119724 79192 153290 79248
rect 153346 79192 153351 79248
rect 119724 79190 153351 79192
rect 119724 79188 119730 79190
rect 153285 79187 153351 79190
rect 156045 79250 156111 79253
rect 156638 79250 156644 79252
rect 156045 79248 156644 79250
rect 156045 79192 156050 79248
rect 156106 79192 156644 79248
rect 156045 79190 156644 79192
rect 156045 79187 156111 79190
rect 156638 79188 156644 79190
rect 156708 79188 156714 79252
rect 157793 79250 157859 79253
rect 158110 79250 158116 79252
rect 157793 79248 158116 79250
rect 157793 79192 157798 79248
rect 157854 79192 158116 79248
rect 157793 79190 158116 79192
rect 157793 79187 157859 79190
rect 158110 79188 158116 79190
rect 158180 79188 158186 79252
rect 158670 79250 158730 79734
rect 158897 79731 158963 79734
rect 159038 79658 159098 79904
rect 159311 79901 159377 79904
rect 159495 79930 159561 79933
rect 159955 79932 160021 79933
rect 159950 79930 159956 79932
rect 159495 79928 159604 79930
rect 159495 79872 159500 79928
rect 159556 79872 159604 79928
rect 159495 79867 159604 79872
rect 159864 79870 159956 79930
rect 159950 79868 159956 79870
rect 160020 79868 160026 79932
rect 160323 79928 160389 79933
rect 160323 79872 160328 79928
rect 160384 79872 160389 79928
rect 159955 79867 160021 79868
rect 160323 79867 160389 79872
rect 159265 79658 159331 79661
rect 159038 79656 159331 79658
rect 159038 79600 159270 79656
rect 159326 79600 159331 79656
rect 159038 79598 159331 79600
rect 159265 79595 159331 79598
rect 158805 79522 158871 79525
rect 158805 79520 158914 79522
rect 158805 79464 158810 79520
rect 158866 79464 158914 79520
rect 158805 79459 158914 79464
rect 158854 79386 158914 79459
rect 159544 79386 159604 79867
rect 159771 79794 159837 79797
rect 159909 79794 159975 79797
rect 159771 79792 159975 79794
rect 159771 79736 159776 79792
rect 159832 79736 159914 79792
rect 159970 79736 159975 79792
rect 159771 79734 159975 79736
rect 159771 79731 159837 79734
rect 159909 79731 159975 79734
rect 160326 79661 160386 79867
rect 160510 79797 160570 80142
rect 168238 80142 187740 80202
rect 168238 79967 168298 80142
rect 187734 80140 187740 80142
rect 187804 80202 187810 80204
rect 188286 80202 188292 80204
rect 187804 80142 188292 80202
rect 187804 80140 187810 80142
rect 188286 80140 188292 80142
rect 188356 80140 188362 80204
rect 170438 80066 170444 80068
rect 170400 80004 170444 80066
rect 170508 80004 170514 80068
rect 176510 80066 176516 80068
rect 175828 80006 176516 80066
rect 161795 79962 161861 79967
rect 160875 79930 160941 79933
rect 161054 79930 161060 79932
rect 160875 79928 161060 79930
rect 160875 79872 160880 79928
rect 160936 79872 161060 79928
rect 160875 79870 161060 79872
rect 160875 79867 160941 79870
rect 161054 79868 161060 79870
rect 161124 79868 161130 79932
rect 161795 79906 161800 79962
rect 161856 79906 161861 79962
rect 165659 79962 165725 79967
rect 161795 79901 161861 79906
rect 160461 79792 160570 79797
rect 160461 79736 160466 79792
rect 160522 79736 160570 79792
rect 160461 79734 160570 79736
rect 160461 79731 160527 79734
rect 161238 79732 161244 79796
rect 161308 79794 161314 79796
rect 161427 79794 161493 79797
rect 161308 79792 161493 79794
rect 161308 79736 161432 79792
rect 161488 79736 161493 79792
rect 161308 79734 161493 79736
rect 161308 79732 161314 79734
rect 161427 79731 161493 79734
rect 161798 79661 161858 79901
rect 162158 79868 162164 79932
rect 162228 79930 162234 79932
rect 162807 79930 162873 79933
rect 162228 79928 162873 79930
rect 162228 79872 162812 79928
rect 162868 79872 162873 79928
rect 162228 79870 162873 79872
rect 162228 79868 162234 79870
rect 162807 79867 162873 79870
rect 163083 79930 163149 79933
rect 163262 79930 163268 79932
rect 163083 79928 163268 79930
rect 163083 79872 163088 79928
rect 163144 79872 163268 79928
rect 163083 79870 163268 79872
rect 163083 79867 163149 79870
rect 163262 79868 163268 79870
rect 163332 79868 163338 79932
rect 163446 79868 163452 79932
rect 163516 79930 163522 79932
rect 163911 79930 163977 79933
rect 164555 79932 164621 79933
rect 164550 79930 164556 79932
rect 163516 79928 163977 79930
rect 163516 79872 163916 79928
rect 163972 79872 163977 79928
rect 163516 79870 163977 79872
rect 163516 79868 163522 79870
rect 163911 79867 163977 79870
rect 164187 79894 164253 79899
rect 164187 79838 164192 79894
rect 164248 79838 164253 79894
rect 164464 79870 164556 79930
rect 164550 79868 164556 79870
rect 164620 79868 164626 79932
rect 164739 79928 164805 79933
rect 164739 79872 164744 79928
rect 164800 79872 164805 79928
rect 164555 79867 164621 79868
rect 164739 79867 164805 79872
rect 165015 79930 165081 79933
rect 165286 79930 165292 79932
rect 165015 79928 165292 79930
rect 165015 79872 165020 79928
rect 165076 79872 165292 79928
rect 165015 79870 165292 79872
rect 165015 79867 165081 79870
rect 165286 79868 165292 79870
rect 165356 79868 165362 79932
rect 165659 79906 165664 79962
rect 165720 79906 165725 79962
rect 166027 79962 166093 79967
rect 166027 79932 166032 79962
rect 166088 79932 166093 79962
rect 168235 79962 168301 79967
rect 165659 79901 165725 79906
rect 165475 79894 165541 79899
rect 164187 79833 164253 79838
rect 162531 79796 162597 79797
rect 162526 79794 162532 79796
rect 162440 79734 162532 79794
rect 162526 79732 162532 79734
rect 162596 79732 162602 79796
rect 162899 79792 162965 79797
rect 162899 79736 162904 79792
rect 162960 79736 162965 79792
rect 162531 79731 162597 79732
rect 162899 79731 162965 79736
rect 162902 79661 162962 79731
rect 160326 79656 160435 79661
rect 160326 79600 160374 79656
rect 160430 79600 160435 79656
rect 160326 79598 160435 79600
rect 161798 79656 161907 79661
rect 161798 79600 161846 79656
rect 161902 79600 161907 79656
rect 161798 79598 161907 79600
rect 162902 79656 163011 79661
rect 162902 79600 162950 79656
rect 163006 79600 163011 79656
rect 162902 79598 163011 79600
rect 160369 79595 160435 79598
rect 161841 79595 161907 79598
rect 162945 79595 163011 79598
rect 163630 79596 163636 79660
rect 163700 79658 163706 79660
rect 164190 79658 164250 79833
rect 164742 79794 164802 79867
rect 165475 79838 165480 79894
rect 165536 79838 165541 79894
rect 165475 79833 165541 79838
rect 165102 79794 165108 79796
rect 164742 79734 165108 79794
rect 165102 79732 165108 79734
rect 165172 79732 165178 79796
rect 165478 79661 165538 79833
rect 165662 79794 165722 79901
rect 166022 79868 166028 79932
rect 166092 79930 166098 79932
rect 166092 79870 166150 79930
rect 166092 79868 166098 79870
rect 166574 79868 166580 79932
rect 166644 79930 166650 79932
rect 166947 79930 167013 79933
rect 166644 79928 167013 79930
rect 166644 79872 166952 79928
rect 167008 79872 167013 79928
rect 166644 79870 167013 79872
rect 166644 79868 166650 79870
rect 166947 79867 167013 79870
rect 167315 79928 167381 79933
rect 167867 79932 167933 79933
rect 167862 79930 167868 79932
rect 167315 79872 167320 79928
rect 167376 79872 167381 79928
rect 167315 79867 167381 79872
rect 167776 79870 167868 79930
rect 167862 79868 167868 79870
rect 167932 79868 167938 79932
rect 168235 79906 168240 79962
rect 168296 79906 168301 79962
rect 169799 79964 169865 79967
rect 169799 79962 169908 79964
rect 168603 79930 168669 79933
rect 168235 79901 168301 79906
rect 168422 79928 168669 79930
rect 168422 79872 168608 79928
rect 168664 79872 168669 79928
rect 168422 79870 168669 79872
rect 167867 79867 167933 79868
rect 166758 79794 166764 79796
rect 165662 79734 166764 79794
rect 166758 79732 166764 79734
rect 166828 79732 166834 79796
rect 166993 79794 167059 79797
rect 167318 79794 167378 79867
rect 168422 79797 168482 79870
rect 168603 79867 168669 79870
rect 168971 79930 169037 79933
rect 169615 79930 169681 79933
rect 168971 79928 169402 79930
rect 168971 79872 168976 79928
rect 169032 79872 169402 79928
rect 168971 79870 169402 79872
rect 168971 79867 169037 79870
rect 167683 79796 167749 79797
rect 168051 79796 168117 79797
rect 167678 79794 167684 79796
rect 166993 79792 167378 79794
rect 166993 79736 166998 79792
rect 167054 79736 167378 79792
rect 166993 79734 167378 79736
rect 167592 79734 167684 79794
rect 166993 79731 167059 79734
rect 167678 79732 167684 79734
rect 167748 79732 167754 79796
rect 168046 79794 168052 79796
rect 167960 79734 168052 79794
rect 168046 79732 168052 79734
rect 168116 79732 168122 79796
rect 168373 79792 168482 79797
rect 168373 79736 168378 79792
rect 168434 79736 168482 79792
rect 168373 79734 168482 79736
rect 168695 79794 168761 79797
rect 168695 79792 169218 79794
rect 168695 79736 168700 79792
rect 168756 79736 169218 79792
rect 168695 79734 169218 79736
rect 167683 79731 167749 79732
rect 168051 79731 168117 79732
rect 168373 79731 168439 79734
rect 168695 79731 168761 79734
rect 163700 79598 164250 79658
rect 165429 79656 165538 79661
rect 165429 79600 165434 79656
rect 165490 79600 165538 79656
rect 165429 79598 165538 79600
rect 163700 79596 163706 79598
rect 165429 79595 165495 79598
rect 166390 79596 166396 79660
rect 166460 79658 166466 79660
rect 166625 79658 166691 79661
rect 166460 79656 166691 79658
rect 166460 79600 166630 79656
rect 166686 79600 166691 79656
rect 166460 79598 166691 79600
rect 166460 79596 166466 79598
rect 166625 79595 166691 79598
rect 168465 79522 168531 79525
rect 168741 79522 168807 79525
rect 168465 79520 168807 79522
rect 168465 79464 168470 79520
rect 168526 79464 168746 79520
rect 168802 79464 168807 79520
rect 168465 79462 168807 79464
rect 169158 79522 169218 79734
rect 169342 79658 169402 79870
rect 169480 79928 169681 79930
rect 169480 79872 169620 79928
rect 169676 79872 169681 79928
rect 169799 79906 169804 79962
rect 169860 79930 169908 79962
rect 170400 79933 170460 80004
rect 170719 79964 170785 79967
rect 173847 79964 173913 79967
rect 170719 79962 170828 79964
rect 170070 79930 170076 79932
rect 169860 79906 170076 79930
rect 169799 79901 170076 79906
rect 169480 79870 169681 79872
rect 169848 79870 170076 79901
rect 169480 79794 169540 79870
rect 169615 79867 169681 79870
rect 170070 79868 170076 79870
rect 170140 79868 170146 79932
rect 170351 79928 170460 79933
rect 170351 79872 170356 79928
rect 170412 79872 170460 79928
rect 170351 79870 170460 79872
rect 170535 79930 170601 79933
rect 170535 79928 170644 79930
rect 170535 79872 170540 79928
rect 170596 79872 170644 79928
rect 170719 79906 170724 79962
rect 170780 79930 170828 79962
rect 173804 79962 173913 79964
rect 170990 79930 170996 79932
rect 170780 79906 170996 79930
rect 170719 79901 170996 79906
rect 170351 79867 170417 79870
rect 170535 79867 170644 79872
rect 170768 79870 170996 79901
rect 170990 79868 170996 79870
rect 171060 79868 171066 79932
rect 171271 79930 171337 79933
rect 171910 79930 171916 79932
rect 171271 79928 171916 79930
rect 171271 79872 171276 79928
rect 171332 79872 171916 79928
rect 171271 79870 171916 79872
rect 171271 79867 171337 79870
rect 171910 79868 171916 79870
rect 171980 79868 171986 79932
rect 172094 79868 172100 79932
rect 172164 79930 172170 79932
rect 172467 79930 172533 79933
rect 172164 79928 172533 79930
rect 172164 79872 172472 79928
rect 172528 79872 172533 79928
rect 172164 79870 172533 79872
rect 172164 79868 172170 79870
rect 172467 79867 172533 79870
rect 173566 79868 173572 79932
rect 173636 79930 173642 79932
rect 173804 79930 173852 79962
rect 173636 79906 173852 79930
rect 173908 79906 173913 79962
rect 174859 79962 174925 79967
rect 173636 79901 173913 79906
rect 174215 79930 174281 79933
rect 174670 79930 174676 79932
rect 174215 79928 174676 79930
rect 173636 79870 173864 79901
rect 174215 79872 174220 79928
rect 174276 79872 174676 79928
rect 174215 79870 174676 79872
rect 173636 79868 173642 79870
rect 174215 79867 174281 79870
rect 174670 79868 174676 79870
rect 174740 79868 174746 79932
rect 174859 79906 174864 79962
rect 174920 79906 174925 79962
rect 174859 79901 174925 79906
rect 175319 79930 175385 79933
rect 175828 79930 175888 80006
rect 176510 80004 176516 80006
rect 176580 80004 176586 80068
rect 205766 80004 205772 80068
rect 205836 80066 205842 80068
rect 206645 80066 206711 80069
rect 205836 80064 206711 80066
rect 205836 80008 206650 80064
rect 206706 80008 206711 80064
rect 205836 80006 206711 80008
rect 205836 80004 205842 80006
rect 206645 80003 206711 80006
rect 176791 79962 176857 79967
rect 175319 79928 175888 79930
rect 170070 79794 170076 79796
rect 169480 79734 170076 79794
rect 170070 79732 170076 79734
rect 170140 79732 170146 79796
rect 170584 79794 170644 79867
rect 174862 79797 174922 79901
rect 175319 79872 175324 79928
rect 175380 79872 175888 79928
rect 175319 79870 175888 79872
rect 175319 79867 175385 79870
rect 175958 79868 175964 79932
rect 176028 79930 176034 79932
rect 176028 79899 176670 79930
rect 176791 79906 176796 79962
rect 176852 79930 176857 79962
rect 177849 79930 177915 79933
rect 176852 79928 177915 79930
rect 176852 79906 177854 79928
rect 176791 79901 177854 79906
rect 176028 79894 176673 79899
rect 176028 79870 176612 79894
rect 176028 79868 176034 79870
rect 176607 79838 176612 79870
rect 176668 79838 176673 79894
rect 176794 79872 177854 79901
rect 177910 79872 177915 79928
rect 176794 79870 177915 79872
rect 177849 79867 177915 79870
rect 176607 79833 176673 79838
rect 171174 79794 171180 79796
rect 170584 79734 171180 79794
rect 171174 79732 171180 79734
rect 171244 79732 171250 79796
rect 172513 79794 172579 79797
rect 171366 79792 172579 79794
rect 171366 79736 172518 79792
rect 172574 79736 172579 79792
rect 171366 79734 172579 79736
rect 169477 79658 169543 79661
rect 170121 79658 170187 79661
rect 171366 79658 171426 79734
rect 172513 79731 172579 79734
rect 173065 79794 173131 79797
rect 173065 79792 173450 79794
rect 173065 79736 173070 79792
rect 173126 79736 173450 79792
rect 173065 79734 173450 79736
rect 173065 79731 173131 79734
rect 169342 79656 169543 79658
rect 169342 79600 169482 79656
rect 169538 79600 169543 79656
rect 169342 79598 169543 79600
rect 169477 79595 169543 79598
rect 169848 79656 170187 79658
rect 169848 79600 170126 79656
rect 170182 79600 170187 79656
rect 169848 79598 170187 79600
rect 169848 79525 169908 79598
rect 170121 79595 170187 79598
rect 170262 79598 171426 79658
rect 171961 79658 172027 79661
rect 173390 79658 173450 79734
rect 174486 79732 174492 79796
rect 174556 79794 174562 79796
rect 174721 79794 174787 79797
rect 174556 79792 174787 79794
rect 174556 79736 174726 79792
rect 174782 79736 174787 79792
rect 174556 79734 174787 79736
rect 174862 79792 174971 79797
rect 174862 79736 174910 79792
rect 174966 79736 174971 79792
rect 174862 79734 174971 79736
rect 174556 79732 174562 79734
rect 174721 79731 174787 79734
rect 174905 79731 174971 79734
rect 176055 79794 176121 79797
rect 177665 79794 177731 79797
rect 180977 79794 181043 79797
rect 176055 79792 176532 79794
rect 176055 79736 176060 79792
rect 176116 79736 176532 79792
rect 176055 79734 176532 79736
rect 176055 79731 176121 79734
rect 173750 79658 173756 79660
rect 171961 79656 172714 79658
rect 171961 79600 171966 79656
rect 172022 79600 172714 79656
rect 171961 79598 172714 79600
rect 173390 79598 173756 79658
rect 169518 79522 169524 79524
rect 169158 79462 169524 79522
rect 168465 79459 168531 79462
rect 168741 79459 168807 79462
rect 169518 79460 169524 79462
rect 169588 79460 169594 79524
rect 169845 79520 169911 79525
rect 169845 79464 169850 79520
rect 169906 79464 169911 79520
rect 169845 79459 169911 79464
rect 158854 79326 159604 79386
rect 162117 79386 162183 79389
rect 170262 79386 170322 79598
rect 171961 79595 172027 79598
rect 170673 79524 170739 79525
rect 170622 79522 170628 79524
rect 170582 79462 170628 79522
rect 170692 79520 170739 79524
rect 170734 79464 170739 79520
rect 170622 79460 170628 79462
rect 170692 79460 170739 79464
rect 172654 79522 172714 79598
rect 173750 79596 173756 79598
rect 173820 79596 173826 79660
rect 173985 79658 174051 79661
rect 175038 79658 175044 79660
rect 173985 79656 175044 79658
rect 173985 79600 173990 79656
rect 174046 79600 175044 79656
rect 173985 79598 175044 79600
rect 173985 79595 174051 79598
rect 175038 79596 175044 79598
rect 175108 79596 175114 79660
rect 175549 79658 175615 79661
rect 176326 79658 176332 79660
rect 175549 79656 176332 79658
rect 175549 79600 175554 79656
rect 175610 79600 176332 79656
rect 175549 79598 176332 79600
rect 175549 79595 175615 79598
rect 176326 79596 176332 79598
rect 176396 79596 176402 79660
rect 176472 79658 176532 79734
rect 177665 79792 181043 79794
rect 177665 79736 177670 79792
rect 177726 79736 180982 79792
rect 181038 79736 181043 79792
rect 177665 79734 181043 79736
rect 177665 79731 177731 79734
rect 180977 79731 181043 79734
rect 178033 79658 178099 79661
rect 176472 79656 178099 79658
rect 176472 79600 178038 79656
rect 178094 79600 178099 79656
rect 176472 79598 178099 79600
rect 178033 79595 178099 79598
rect 177665 79522 177731 79525
rect 172654 79520 177731 79522
rect 172654 79464 177670 79520
rect 177726 79464 177731 79520
rect 172654 79462 177731 79464
rect 170673 79459 170739 79460
rect 177665 79459 177731 79462
rect 178217 79522 178283 79525
rect 186221 79524 186287 79525
rect 186221 79522 186268 79524
rect 178217 79520 186268 79522
rect 178217 79464 178222 79520
rect 178278 79464 186226 79520
rect 178217 79462 186268 79464
rect 178217 79459 178283 79462
rect 186221 79460 186268 79462
rect 186332 79460 186338 79524
rect 186221 79459 186287 79460
rect 162117 79384 170322 79386
rect 162117 79328 162122 79384
rect 162178 79328 170322 79384
rect 162117 79326 170322 79328
rect 170765 79386 170831 79389
rect 189390 79386 189396 79388
rect 170765 79384 189396 79386
rect 170765 79328 170770 79384
rect 170826 79328 189396 79384
rect 170765 79326 189396 79328
rect 162117 79323 162183 79326
rect 170765 79323 170831 79326
rect 189390 79324 189396 79326
rect 189460 79324 189466 79388
rect 159725 79250 159791 79253
rect 158670 79248 159791 79250
rect 158670 79192 159730 79248
rect 159786 79192 159791 79248
rect 158670 79190 159791 79192
rect 159725 79187 159791 79190
rect 168465 79250 168531 79253
rect 169201 79250 169267 79253
rect 190862 79250 190868 79252
rect 168465 79248 190868 79250
rect 168465 79192 168470 79248
rect 168526 79192 169206 79248
rect 169262 79192 190868 79248
rect 168465 79190 190868 79192
rect 168465 79187 168531 79190
rect 169201 79187 169267 79190
rect 190862 79188 190868 79190
rect 190932 79188 190938 79252
rect 120942 79052 120948 79116
rect 121012 79114 121018 79116
rect 155902 79114 155908 79116
rect 121012 79054 155908 79114
rect 121012 79052 121018 79054
rect 155902 79052 155908 79054
rect 155972 79114 155978 79116
rect 162117 79114 162183 79117
rect 171409 79114 171475 79117
rect 194726 79114 194732 79116
rect 155972 79054 160110 79114
rect 155972 79052 155978 79054
rect 100201 78978 100267 78981
rect 134425 78978 134491 78981
rect 100201 78976 134491 78978
rect 100201 78920 100206 78976
rect 100262 78920 134430 78976
rect 134486 78920 134491 78976
rect 100201 78918 134491 78920
rect 100201 78915 100267 78918
rect 134425 78915 134491 78918
rect 143533 78980 143599 78981
rect 143533 78976 143580 78980
rect 143644 78978 143650 78980
rect 143533 78920 143538 78976
rect 143533 78916 143580 78920
rect 143644 78918 143690 78978
rect 143644 78916 143650 78918
rect 143533 78915 143599 78916
rect 116485 78842 116551 78845
rect 151261 78842 151327 78845
rect 116485 78840 151327 78842
rect 116485 78784 116490 78840
rect 116546 78784 151266 78840
rect 151322 78784 151327 78840
rect 116485 78782 151327 78784
rect 116485 78779 116551 78782
rect 151261 78779 151327 78782
rect 158846 78780 158852 78844
rect 158916 78842 158922 78844
rect 159449 78842 159515 78845
rect 158916 78840 159515 78842
rect 158916 78784 159454 78840
rect 159510 78784 159515 78840
rect 158916 78782 159515 78784
rect 160050 78842 160110 79054
rect 162117 79112 171150 79114
rect 162117 79056 162122 79112
rect 162178 79056 171150 79112
rect 162117 79054 171150 79056
rect 162117 79051 162183 79054
rect 171090 78978 171150 79054
rect 171409 79112 194732 79114
rect 171409 79056 171414 79112
rect 171470 79056 194732 79112
rect 171409 79054 194732 79056
rect 171409 79051 171475 79054
rect 194726 79052 194732 79054
rect 194796 79052 194802 79116
rect 173198 78978 173204 78980
rect 171090 78918 173204 78978
rect 173198 78916 173204 78918
rect 173268 78916 173274 78980
rect 173893 78978 173959 78981
rect 203006 78978 203012 78980
rect 173893 78976 203012 78978
rect 173893 78920 173898 78976
rect 173954 78920 203012 78976
rect 173893 78918 203012 78920
rect 173893 78915 173959 78918
rect 203006 78916 203012 78918
rect 203076 78916 203082 78980
rect 171133 78842 171199 78845
rect 175089 78842 175155 78845
rect 160050 78782 169770 78842
rect 158916 78780 158922 78782
rect 159449 78779 159515 78782
rect 115013 78706 115079 78709
rect 149329 78706 149395 78709
rect 115013 78704 149395 78706
rect 115013 78648 115018 78704
rect 115074 78648 149334 78704
rect 149390 78648 149395 78704
rect 115013 78646 149395 78648
rect 115013 78643 115079 78646
rect 149329 78643 149395 78646
rect 158294 78644 158300 78708
rect 158364 78706 158370 78708
rect 158897 78706 158963 78709
rect 158364 78704 158963 78706
rect 158364 78648 158902 78704
rect 158958 78648 158963 78704
rect 158364 78646 158963 78648
rect 158364 78644 158370 78646
rect 158897 78643 158963 78646
rect 159541 78706 159607 78709
rect 159950 78706 159956 78708
rect 159541 78704 159956 78706
rect 159541 78648 159546 78704
rect 159602 78648 159956 78704
rect 159541 78646 159956 78648
rect 159541 78643 159607 78646
rect 159950 78644 159956 78646
rect 160020 78644 160026 78708
rect 169710 78706 169770 78782
rect 171133 78840 175155 78842
rect 171133 78784 171138 78840
rect 171194 78784 175094 78840
rect 175150 78784 175155 78840
rect 171133 78782 175155 78784
rect 171133 78779 171199 78782
rect 175089 78779 175155 78782
rect 176285 78842 176351 78845
rect 206461 78842 206527 78845
rect 176285 78840 206527 78842
rect 176285 78784 176290 78840
rect 176346 78784 206466 78840
rect 206522 78784 206527 78840
rect 176285 78782 206527 78784
rect 176285 78779 176351 78782
rect 206461 78779 206527 78782
rect 302233 78706 302299 78709
rect 169710 78704 302299 78706
rect 169710 78648 302238 78704
rect 302294 78648 302299 78704
rect 169710 78646 302299 78648
rect 302233 78643 302299 78646
rect 103145 78570 103211 78573
rect 128997 78570 129063 78573
rect 103145 78568 129063 78570
rect 103145 78512 103150 78568
rect 103206 78512 129002 78568
rect 129058 78512 129063 78568
rect 103145 78510 129063 78512
rect 103145 78507 103211 78510
rect 20713 78162 20779 78165
rect 103470 78162 103530 78510
rect 128997 78507 129063 78510
rect 134149 78572 134215 78573
rect 134149 78568 134196 78572
rect 134260 78570 134266 78572
rect 137921 78570 137987 78573
rect 138422 78570 138428 78572
rect 134149 78512 134154 78568
rect 134149 78508 134196 78512
rect 134260 78510 134306 78570
rect 137921 78568 138428 78570
rect 137921 78512 137926 78568
rect 137982 78512 138428 78568
rect 137921 78510 138428 78512
rect 134260 78508 134266 78510
rect 134149 78507 134215 78508
rect 137921 78507 137987 78510
rect 138422 78508 138428 78510
rect 138492 78508 138498 78572
rect 139342 78508 139348 78572
rect 139412 78570 139418 78572
rect 139577 78570 139643 78573
rect 139412 78568 139643 78570
rect 139412 78512 139582 78568
rect 139638 78512 139643 78568
rect 139412 78510 139643 78512
rect 139412 78508 139418 78510
rect 139577 78507 139643 78510
rect 148358 78508 148364 78572
rect 148428 78570 148434 78572
rect 149053 78570 149119 78573
rect 148428 78568 149119 78570
rect 148428 78512 149058 78568
rect 149114 78512 149119 78568
rect 148428 78510 149119 78512
rect 148428 78508 148434 78510
rect 149053 78507 149119 78510
rect 149462 78508 149468 78572
rect 149532 78570 149538 78572
rect 150433 78570 150499 78573
rect 149532 78568 150499 78570
rect 149532 78512 150438 78568
rect 150494 78512 150499 78568
rect 149532 78510 150499 78512
rect 149532 78508 149538 78510
rect 150433 78507 150499 78510
rect 170489 78570 170555 78573
rect 171041 78572 171107 78573
rect 170806 78570 170812 78572
rect 170489 78568 170812 78570
rect 170489 78512 170494 78568
rect 170550 78512 170812 78568
rect 170489 78510 170812 78512
rect 170489 78507 170555 78510
rect 170806 78508 170812 78510
rect 170876 78508 170882 78572
rect 170990 78508 170996 78572
rect 171060 78570 171107 78572
rect 171060 78568 171152 78570
rect 171102 78512 171152 78568
rect 171060 78510 171152 78512
rect 171060 78508 171107 78510
rect 176326 78508 176332 78572
rect 176396 78570 176402 78572
rect 176469 78570 176535 78573
rect 176396 78568 176535 78570
rect 176396 78512 176474 78568
rect 176530 78512 176535 78568
rect 176396 78510 176535 78512
rect 176396 78508 176402 78510
rect 171041 78507 171107 78508
rect 176469 78507 176535 78510
rect 178033 78570 178099 78573
rect 183461 78570 183527 78573
rect 178033 78568 183527 78570
rect 178033 78512 178038 78568
rect 178094 78512 183466 78568
rect 183522 78512 183527 78568
rect 178033 78510 183527 78512
rect 178033 78507 178099 78510
rect 183461 78507 183527 78510
rect 186221 78570 186287 78573
rect 187601 78570 187667 78573
rect 186221 78568 187667 78570
rect 186221 78512 186226 78568
rect 186282 78512 187606 78568
rect 187662 78512 187667 78568
rect 186221 78510 187667 78512
rect 186221 78507 186287 78510
rect 187601 78507 187667 78510
rect 128537 78434 128603 78437
rect 20713 78160 103530 78162
rect 20713 78104 20718 78160
rect 20774 78104 103530 78160
rect 20713 78102 103530 78104
rect 107518 78432 128603 78434
rect 107518 78376 128542 78432
rect 128598 78376 128603 78432
rect 107518 78374 128603 78376
rect 20713 78099 20779 78102
rect 6913 78026 6979 78029
rect 105629 78026 105695 78029
rect 107518 78026 107578 78374
rect 128537 78371 128603 78374
rect 134006 78372 134012 78436
rect 134076 78434 134082 78436
rect 134149 78434 134215 78437
rect 134076 78432 134215 78434
rect 134076 78376 134154 78432
rect 134210 78376 134215 78432
rect 134076 78374 134215 78376
rect 134076 78372 134082 78374
rect 134149 78371 134215 78374
rect 168557 78434 168623 78437
rect 202965 78434 203031 78437
rect 465165 78434 465231 78437
rect 168557 78432 465231 78434
rect 168557 78376 168562 78432
rect 168618 78376 202970 78432
rect 203026 78376 465170 78432
rect 465226 78376 465231 78432
rect 168557 78374 465231 78376
rect 168557 78371 168623 78374
rect 202965 78371 203031 78374
rect 465165 78371 465231 78374
rect 6913 78024 107578 78026
rect 6913 77968 6918 78024
rect 6974 77968 105634 78024
rect 105690 77968 107578 78024
rect 6913 77966 107578 77968
rect 108990 78238 122850 78298
rect 6913 77963 6979 77966
rect 105629 77963 105695 77966
rect 2773 77890 2839 77893
rect 107510 77890 107516 77892
rect 2773 77888 107516 77890
rect 2773 77832 2778 77888
rect 2834 77832 107516 77888
rect 2773 77830 107516 77832
rect 2773 77827 2839 77830
rect 107510 77828 107516 77830
rect 107580 77890 107586 77892
rect 108990 77890 109050 78238
rect 122790 78162 122850 78238
rect 122966 78236 122972 78300
rect 123036 78298 123042 78300
rect 124121 78298 124187 78301
rect 132493 78298 132559 78301
rect 123036 78296 124187 78298
rect 123036 78240 124126 78296
rect 124182 78240 124187 78296
rect 123036 78238 124187 78240
rect 123036 78236 123042 78238
rect 124121 78235 124187 78238
rect 124262 78296 132559 78298
rect 124262 78240 132498 78296
rect 132554 78240 132559 78296
rect 124262 78238 132559 78240
rect 124262 78162 124322 78238
rect 132493 78235 132559 78238
rect 134006 78236 134012 78300
rect 134076 78298 134082 78300
rect 134333 78298 134399 78301
rect 134076 78296 134399 78298
rect 134076 78240 134338 78296
rect 134394 78240 134399 78296
rect 134076 78238 134399 78240
rect 134076 78236 134082 78238
rect 134333 78235 134399 78238
rect 136725 78298 136791 78301
rect 137502 78298 137508 78300
rect 136725 78296 137508 78298
rect 136725 78240 136730 78296
rect 136786 78240 137508 78296
rect 136725 78238 137508 78240
rect 136725 78235 136791 78238
rect 137502 78236 137508 78238
rect 137572 78236 137578 78300
rect 140814 78236 140820 78300
rect 140884 78298 140890 78300
rect 141417 78298 141483 78301
rect 140884 78296 141483 78298
rect 140884 78240 141422 78296
rect 141478 78240 141483 78296
rect 140884 78238 141483 78240
rect 140884 78236 140890 78238
rect 141417 78235 141483 78238
rect 156229 78298 156295 78301
rect 157006 78298 157012 78300
rect 156229 78296 157012 78298
rect 156229 78240 156234 78296
rect 156290 78240 157012 78296
rect 156229 78238 157012 78240
rect 156229 78235 156295 78238
rect 157006 78236 157012 78238
rect 157076 78236 157082 78300
rect 167913 78298 167979 78301
rect 190494 78298 190500 78300
rect 167913 78296 190500 78298
rect 167913 78240 167918 78296
rect 167974 78240 190500 78296
rect 167913 78238 190500 78240
rect 167913 78235 167979 78238
rect 190494 78236 190500 78238
rect 190564 78298 190570 78300
rect 456793 78298 456859 78301
rect 190564 78296 456859 78298
rect 190564 78240 456798 78296
rect 456854 78240 456859 78296
rect 190564 78238 456859 78240
rect 190564 78236 190570 78238
rect 456793 78235 456859 78238
rect 141693 78162 141759 78165
rect 122790 78102 124322 78162
rect 128310 78160 141759 78162
rect 128310 78104 141698 78160
rect 141754 78104 141759 78160
rect 128310 78102 141759 78104
rect 107580 77830 109050 77890
rect 126973 77890 127039 77893
rect 128310 77890 128370 78102
rect 141693 78099 141759 78102
rect 149830 78100 149836 78164
rect 149900 78162 149906 78164
rect 151077 78162 151143 78165
rect 149900 78160 151143 78162
rect 149900 78104 151082 78160
rect 151138 78104 151143 78160
rect 149900 78102 151143 78104
rect 149900 78100 149906 78102
rect 151077 78099 151143 78102
rect 154849 78162 154915 78165
rect 154982 78162 154988 78164
rect 154849 78160 154988 78162
rect 154849 78104 154854 78160
rect 154910 78104 154988 78160
rect 154849 78102 154988 78104
rect 154849 78099 154915 78102
rect 154982 78100 154988 78102
rect 155052 78100 155058 78164
rect 171869 78162 171935 78165
rect 203701 78162 203767 78165
rect 471973 78162 472039 78165
rect 171869 78160 472039 78162
rect 171869 78104 171874 78160
rect 171930 78104 203706 78160
rect 203762 78104 471978 78160
rect 472034 78104 472039 78160
rect 171869 78102 472039 78104
rect 171869 78099 171935 78102
rect 203701 78099 203767 78102
rect 471973 78099 472039 78102
rect 130837 78026 130903 78029
rect 138933 78028 138999 78029
rect 138933 78026 138980 78028
rect 130837 78024 134810 78026
rect 130837 77968 130842 78024
rect 130898 77968 134810 78024
rect 130837 77966 134810 77968
rect 138888 78024 138980 78026
rect 138888 77968 138938 78024
rect 138888 77966 138980 77968
rect 130837 77963 130903 77966
rect 126973 77888 128370 77890
rect 126973 77832 126978 77888
rect 127034 77832 128370 77888
rect 126973 77830 128370 77832
rect 129641 77890 129707 77893
rect 134517 77890 134583 77893
rect 129641 77888 134583 77890
rect 129641 77832 129646 77888
rect 129702 77832 134522 77888
rect 134578 77832 134583 77888
rect 129641 77830 134583 77832
rect 134750 77890 134810 77966
rect 138933 77964 138980 77966
rect 139044 77964 139050 78028
rect 143758 77964 143764 78028
rect 143828 78026 143834 78028
rect 144453 78026 144519 78029
rect 143828 78024 144519 78026
rect 143828 77968 144458 78024
rect 144514 77968 144519 78024
rect 143828 77966 144519 77968
rect 143828 77964 143834 77966
rect 138933 77963 138999 77964
rect 144453 77963 144519 77966
rect 155718 77964 155724 78028
rect 155788 78026 155794 78028
rect 155953 78026 156019 78029
rect 155788 78024 156019 78026
rect 155788 77968 155958 78024
rect 156014 77968 156019 78024
rect 155788 77966 156019 77968
rect 155788 77964 155794 77966
rect 155953 77963 156019 77966
rect 177481 78026 177547 78029
rect 211981 78026 212047 78029
rect 580993 78026 581059 78029
rect 177481 78024 581059 78026
rect 177481 77968 177486 78024
rect 177542 77968 211986 78024
rect 212042 77968 580998 78024
rect 581054 77968 581059 78024
rect 177481 77966 581059 77968
rect 177481 77963 177547 77966
rect 211981 77963 212047 77966
rect 580993 77963 581059 77966
rect 140497 77890 140563 77893
rect 134750 77888 140563 77890
rect 134750 77832 140502 77888
rect 140558 77832 140563 77888
rect 134750 77830 140563 77832
rect 107580 77828 107586 77830
rect 126973 77827 127039 77830
rect 129641 77827 129707 77830
rect 134517 77827 134583 77830
rect 140497 77827 140563 77830
rect 140998 77828 141004 77892
rect 141068 77890 141074 77892
rect 141417 77890 141483 77893
rect 141068 77888 141483 77890
rect 141068 77832 141422 77888
rect 141478 77832 141483 77888
rect 141068 77830 141483 77832
rect 141068 77828 141074 77830
rect 141417 77827 141483 77830
rect 142153 77890 142219 77893
rect 142654 77890 142660 77892
rect 142153 77888 142660 77890
rect 142153 77832 142158 77888
rect 142214 77832 142660 77888
rect 142153 77830 142660 77832
rect 142153 77827 142219 77830
rect 142654 77828 142660 77830
rect 142724 77828 142730 77892
rect 143942 77828 143948 77892
rect 144012 77890 144018 77892
rect 144637 77890 144703 77893
rect 144012 77888 144703 77890
rect 144012 77832 144642 77888
rect 144698 77832 144703 77888
rect 144012 77830 144703 77832
rect 144012 77828 144018 77830
rect 144637 77827 144703 77830
rect 177573 77890 177639 77893
rect 211889 77890 211955 77893
rect 581085 77890 581151 77893
rect 177573 77888 581151 77890
rect 177573 77832 177578 77888
rect 177634 77832 211894 77888
rect 211950 77832 581090 77888
rect 581146 77832 581151 77888
rect 177573 77830 581151 77832
rect 177573 77827 177639 77830
rect 211889 77827 211955 77830
rect 581085 77827 581151 77830
rect 133321 77756 133387 77757
rect 133270 77754 133276 77756
rect 133230 77694 133276 77754
rect 133340 77752 133387 77756
rect 133382 77696 133387 77752
rect 133270 77692 133276 77694
rect 133340 77692 133387 77696
rect 133321 77691 133387 77692
rect 175733 77754 175799 77757
rect 176142 77754 176148 77756
rect 175733 77752 176148 77754
rect 175733 77696 175738 77752
rect 175794 77696 176148 77752
rect 175733 77694 176148 77696
rect 175733 77691 175799 77694
rect 176142 77692 176148 77694
rect 176212 77692 176218 77756
rect 187693 77754 187759 77757
rect 188102 77754 188108 77756
rect 187693 77752 188108 77754
rect 187693 77696 187698 77752
rect 187754 77696 188108 77752
rect 187693 77694 188108 77696
rect 187693 77691 187759 77694
rect 188102 77692 188108 77694
rect 188172 77692 188178 77756
rect 129549 77618 129615 77621
rect 129549 77616 133706 77618
rect 129549 77560 129554 77616
rect 129610 77560 133706 77616
rect 129549 77558 133706 77560
rect 129549 77555 129615 77558
rect 133646 77482 133706 77558
rect 135294 77556 135300 77620
rect 135364 77618 135370 77620
rect 135805 77618 135871 77621
rect 135364 77616 135871 77618
rect 135364 77560 135810 77616
rect 135866 77560 135871 77616
rect 135364 77558 135871 77560
rect 135364 77556 135370 77558
rect 135805 77555 135871 77558
rect 147990 77556 147996 77620
rect 148060 77618 148066 77620
rect 148961 77618 149027 77621
rect 148060 77616 149027 77618
rect 148060 77560 148966 77616
rect 149022 77560 149027 77616
rect 148060 77558 149027 77560
rect 148060 77556 148066 77558
rect 148961 77555 149027 77558
rect 175825 77618 175891 77621
rect 176009 77618 176075 77621
rect 175825 77616 176075 77618
rect 175825 77560 175830 77616
rect 175886 77560 176014 77616
rect 176070 77560 176075 77616
rect 175825 77558 176075 77560
rect 175825 77555 175891 77558
rect 176009 77555 176075 77558
rect 142337 77482 142403 77485
rect 133646 77480 142403 77482
rect 133646 77424 142342 77480
rect 142398 77424 142403 77480
rect 133646 77422 142403 77424
rect 142337 77419 142403 77422
rect 146886 77420 146892 77484
rect 146956 77482 146962 77484
rect 147029 77482 147095 77485
rect 148593 77484 148659 77485
rect 146956 77480 147095 77482
rect 146956 77424 147034 77480
rect 147090 77424 147095 77480
rect 146956 77422 147095 77424
rect 146956 77420 146962 77422
rect 147029 77419 147095 77422
rect 148542 77420 148548 77484
rect 148612 77482 148659 77484
rect 148612 77480 148704 77482
rect 148654 77424 148704 77480
rect 148612 77422 148704 77424
rect 148612 77420 148659 77422
rect 150014 77420 150020 77484
rect 150084 77482 150090 77484
rect 150341 77482 150407 77485
rect 150084 77480 150407 77482
rect 150084 77424 150346 77480
rect 150402 77424 150407 77480
rect 150084 77422 150407 77424
rect 150084 77420 150090 77422
rect 148593 77419 148659 77420
rect 150341 77419 150407 77422
rect 150709 77482 150775 77485
rect 151670 77482 151676 77484
rect 150709 77480 151676 77482
rect 150709 77424 150714 77480
rect 150770 77424 151676 77480
rect 150709 77422 151676 77424
rect 150709 77419 150775 77422
rect 151670 77420 151676 77422
rect 151740 77420 151746 77484
rect 152590 77420 152596 77484
rect 152660 77482 152666 77484
rect 152733 77482 152799 77485
rect 152660 77480 152799 77482
rect 152660 77424 152738 77480
rect 152794 77424 152799 77480
rect 152660 77422 152799 77424
rect 152660 77420 152666 77422
rect 152733 77419 152799 77422
rect 169661 77482 169727 77485
rect 183461 77482 183527 77485
rect 184289 77482 184355 77485
rect 169661 77480 179430 77482
rect 169661 77424 169666 77480
rect 169722 77424 179430 77480
rect 169661 77422 179430 77424
rect 169661 77419 169727 77422
rect 130009 77346 130075 77349
rect 130837 77346 130903 77349
rect 130009 77344 130903 77346
rect 130009 77288 130014 77344
rect 130070 77288 130842 77344
rect 130898 77288 130903 77344
rect 130009 77286 130903 77288
rect 130009 77283 130075 77286
rect 130837 77283 130903 77286
rect 134057 77346 134123 77349
rect 134374 77346 134380 77348
rect 134057 77344 134380 77346
rect 134057 77288 134062 77344
rect 134118 77288 134380 77344
rect 134057 77286 134380 77288
rect 134057 77283 134123 77286
rect 134374 77284 134380 77286
rect 134444 77284 134450 77348
rect 135345 77346 135411 77349
rect 135662 77346 135668 77348
rect 135345 77344 135668 77346
rect 135345 77288 135350 77344
rect 135406 77288 135668 77344
rect 135345 77286 135668 77288
rect 135345 77283 135411 77286
rect 135662 77284 135668 77286
rect 135732 77284 135738 77348
rect 147438 77284 147444 77348
rect 147508 77346 147514 77348
rect 147581 77346 147647 77349
rect 147508 77344 147647 77346
rect 147508 77288 147586 77344
rect 147642 77288 147647 77344
rect 147508 77286 147647 77288
rect 147508 77284 147514 77286
rect 147581 77283 147647 77286
rect 147806 77284 147812 77348
rect 147876 77346 147882 77348
rect 148869 77346 148935 77349
rect 149605 77348 149671 77349
rect 149605 77346 149652 77348
rect 147876 77344 148935 77346
rect 147876 77288 148874 77344
rect 148930 77288 148935 77344
rect 147876 77286 148935 77288
rect 149560 77344 149652 77346
rect 149560 77288 149610 77344
rect 149560 77286 149652 77288
rect 147876 77284 147882 77286
rect 148869 77283 148935 77286
rect 149605 77284 149652 77286
rect 149716 77284 149722 77348
rect 149830 77284 149836 77348
rect 149900 77346 149906 77348
rect 150065 77346 150131 77349
rect 149900 77344 150131 77346
rect 149900 77288 150070 77344
rect 150126 77288 150131 77344
rect 149900 77286 150131 77288
rect 149900 77284 149906 77286
rect 149605 77283 149671 77284
rect 150065 77283 150131 77286
rect 164918 77284 164924 77348
rect 164988 77346 164994 77348
rect 165337 77346 165403 77349
rect 164988 77344 165403 77346
rect 164988 77288 165342 77344
rect 165398 77288 165403 77344
rect 164988 77286 165403 77288
rect 179370 77346 179430 77422
rect 183461 77480 184355 77482
rect 183461 77424 183466 77480
rect 183522 77424 184294 77480
rect 184350 77424 184355 77480
rect 183461 77422 184355 77424
rect 183461 77419 183527 77422
rect 184289 77419 184355 77422
rect 209221 77346 209287 77349
rect 179370 77344 209287 77346
rect 179370 77288 209226 77344
rect 209282 77288 209287 77344
rect 179370 77286 209287 77288
rect 164988 77284 164994 77286
rect 165337 77283 165403 77286
rect 209221 77283 209287 77286
rect 119654 77148 119660 77212
rect 119724 77210 119730 77212
rect 154297 77210 154363 77213
rect 119724 77208 154363 77210
rect 119724 77152 154302 77208
rect 154358 77152 154363 77208
rect 119724 77150 154363 77152
rect 119724 77148 119730 77150
rect 154297 77147 154363 77150
rect 162577 77210 162643 77213
rect 162577 77208 169770 77210
rect 162577 77152 162582 77208
rect 162638 77152 169770 77208
rect 162577 77150 169770 77152
rect 162577 77147 162643 77150
rect 100753 77074 100819 77077
rect 101489 77074 101555 77077
rect 134701 77074 134767 77077
rect 100753 77072 134767 77074
rect 100753 77016 100758 77072
rect 100814 77016 101494 77072
rect 101550 77016 134706 77072
rect 134762 77016 134767 77072
rect 100753 77014 134767 77016
rect 169710 77074 169770 77150
rect 174670 77148 174676 77212
rect 174740 77210 174746 77212
rect 174813 77210 174879 77213
rect 174740 77208 174879 77210
rect 174740 77152 174818 77208
rect 174874 77152 174879 77208
rect 174740 77150 174879 77152
rect 174740 77148 174746 77150
rect 174813 77147 174879 77150
rect 209998 77148 210004 77212
rect 210068 77210 210074 77212
rect 210509 77210 210575 77213
rect 210068 77208 210575 77210
rect 210068 77152 210514 77208
rect 210570 77152 210575 77208
rect 210068 77150 210575 77152
rect 210068 77148 210074 77150
rect 210509 77147 210575 77150
rect 214741 77074 214807 77077
rect 169710 77072 215310 77074
rect 169710 77016 214746 77072
rect 214802 77016 215310 77072
rect 169710 77014 215310 77016
rect 100753 77011 100819 77014
rect 101489 77011 101555 77014
rect 134701 77011 134767 77014
rect 214741 77011 214807 77014
rect 109585 76938 109651 76941
rect 140957 76938 141023 76941
rect 109585 76936 141023 76938
rect 109585 76880 109590 76936
rect 109646 76880 140962 76936
rect 141018 76880 141023 76936
rect 109585 76878 141023 76880
rect 109585 76875 109651 76878
rect 140957 76875 141023 76878
rect 160686 76876 160692 76940
rect 160756 76938 160762 76940
rect 161289 76938 161355 76941
rect 160756 76936 161355 76938
rect 160756 76880 161294 76936
rect 161350 76880 161355 76936
rect 160756 76878 161355 76880
rect 160756 76876 160762 76878
rect 161289 76875 161355 76878
rect 164550 76876 164556 76940
rect 164620 76938 164626 76940
rect 165337 76938 165403 76941
rect 164620 76936 165403 76938
rect 164620 76880 165342 76936
rect 165398 76880 165403 76936
rect 164620 76878 165403 76880
rect 164620 76876 164626 76878
rect 165337 76875 165403 76878
rect 167862 76876 167868 76940
rect 167932 76938 167938 76940
rect 168281 76938 168347 76941
rect 167932 76936 168347 76938
rect 167932 76880 168286 76936
rect 168342 76880 168347 76936
rect 167932 76878 168347 76880
rect 167932 76876 167938 76878
rect 168281 76875 168347 76878
rect 172789 76938 172855 76941
rect 173801 76938 173867 76941
rect 199510 76938 199516 76940
rect 172789 76936 199516 76938
rect 172789 76880 172794 76936
rect 172850 76880 173806 76936
rect 173862 76880 199516 76936
rect 172789 76878 199516 76880
rect 172789 76875 172855 76878
rect 173801 76875 173867 76878
rect 199510 76876 199516 76878
rect 199580 76876 199586 76940
rect 118417 76802 118483 76805
rect 151997 76802 152063 76805
rect 152406 76802 152412 76804
rect 118417 76800 142170 76802
rect 118417 76744 118422 76800
rect 118478 76744 142170 76800
rect 118417 76742 142170 76744
rect 118417 76739 118483 76742
rect 67633 76666 67699 76669
rect 111190 76666 111196 76668
rect 67633 76664 111196 76666
rect 67633 76608 67638 76664
rect 67694 76608 111196 76664
rect 67633 76606 111196 76608
rect 67633 76603 67699 76606
rect 111190 76604 111196 76606
rect 111260 76666 111266 76668
rect 111701 76666 111767 76669
rect 111260 76664 111767 76666
rect 111260 76608 111706 76664
rect 111762 76608 111767 76664
rect 111260 76606 111767 76608
rect 111260 76604 111266 76606
rect 111701 76603 111767 76606
rect 133086 76604 133092 76668
rect 133156 76666 133162 76668
rect 133965 76666 134031 76669
rect 133156 76664 134031 76666
rect 133156 76608 133970 76664
rect 134026 76608 134031 76664
rect 133156 76606 134031 76608
rect 142110 76666 142170 76742
rect 151997 76800 152412 76802
rect 151997 76744 152002 76800
rect 152058 76744 152412 76800
rect 151997 76742 152412 76744
rect 151997 76739 152063 76742
rect 152406 76740 152412 76742
rect 152476 76740 152482 76804
rect 160870 76740 160876 76804
rect 160940 76802 160946 76804
rect 161197 76802 161263 76805
rect 160940 76800 161263 76802
rect 160940 76744 161202 76800
rect 161258 76744 161263 76800
rect 160940 76742 161263 76744
rect 160940 76740 160946 76742
rect 161197 76739 161263 76742
rect 162301 76804 162367 76805
rect 162301 76800 162348 76804
rect 162412 76802 162418 76804
rect 164969 76802 165035 76805
rect 165470 76802 165476 76804
rect 162301 76744 162306 76800
rect 162301 76740 162348 76744
rect 162412 76742 162458 76802
rect 164969 76800 165476 76802
rect 164969 76744 164974 76800
rect 165030 76744 165476 76800
rect 164969 76742 165476 76744
rect 162412 76740 162418 76742
rect 162301 76739 162367 76740
rect 164969 76739 165035 76742
rect 165470 76740 165476 76742
rect 165540 76740 165546 76804
rect 165797 76802 165863 76805
rect 167821 76804 167887 76805
rect 169293 76804 169359 76805
rect 166022 76802 166028 76804
rect 165797 76800 166028 76802
rect 165797 76744 165802 76800
rect 165858 76744 166028 76800
rect 165797 76742 166028 76744
rect 165797 76739 165863 76742
rect 166022 76740 166028 76742
rect 166092 76740 166098 76804
rect 167821 76800 167868 76804
rect 167932 76802 167938 76804
rect 167821 76744 167826 76800
rect 167821 76740 167868 76744
rect 167932 76742 167978 76802
rect 169293 76800 169340 76804
rect 169404 76802 169410 76804
rect 169293 76744 169298 76800
rect 167932 76740 167938 76742
rect 169293 76740 169340 76744
rect 169404 76742 169450 76802
rect 169404 76740 169410 76742
rect 170438 76740 170444 76804
rect 170508 76802 170514 76804
rect 170857 76802 170923 76805
rect 193806 76802 193812 76804
rect 170508 76800 193812 76802
rect 170508 76744 170862 76800
rect 170918 76744 193812 76800
rect 170508 76742 193812 76744
rect 170508 76740 170514 76742
rect 167821 76739 167887 76740
rect 169293 76739 169359 76740
rect 170857 76739 170923 76742
rect 193806 76740 193812 76742
rect 193876 76740 193882 76804
rect 146201 76666 146267 76669
rect 178033 76666 178099 76669
rect 142110 76664 178099 76666
rect 142110 76608 146206 76664
rect 146262 76608 178038 76664
rect 178094 76608 178099 76664
rect 142110 76606 178099 76608
rect 133156 76604 133162 76606
rect 133965 76603 134031 76606
rect 146201 76603 146267 76606
rect 178033 76603 178099 76606
rect 178493 76666 178559 76669
rect 179229 76666 179295 76669
rect 191966 76666 191972 76668
rect 178493 76664 191972 76666
rect 178493 76608 178498 76664
rect 178554 76608 179234 76664
rect 179290 76608 191972 76664
rect 178493 76606 191972 76608
rect 178493 76603 178559 76606
rect 179229 76603 179295 76606
rect 191966 76604 191972 76606
rect 192036 76604 192042 76668
rect 34513 76530 34579 76533
rect 100753 76530 100819 76533
rect 34513 76528 100819 76530
rect 34513 76472 34518 76528
rect 34574 76472 100758 76528
rect 100814 76472 100819 76528
rect 34513 76470 100819 76472
rect 34513 76467 34579 76470
rect 100753 76467 100819 76470
rect 151537 76530 151603 76533
rect 193121 76530 193187 76533
rect 209129 76530 209195 76533
rect 151537 76528 209195 76530
rect 151537 76472 151542 76528
rect 151598 76472 193126 76528
rect 193182 76472 209134 76528
rect 209190 76472 209195 76528
rect 151537 76470 209195 76472
rect 215250 76530 215310 77014
rect 217133 76666 217199 76669
rect 217409 76666 217475 76669
rect 260097 76666 260163 76669
rect 217133 76664 260163 76666
rect 217133 76608 217138 76664
rect 217194 76608 217414 76664
rect 217470 76608 260102 76664
rect 260158 76608 260163 76664
rect 217133 76606 260163 76608
rect 217133 76603 217199 76606
rect 217409 76603 217475 76606
rect 260097 76603 260163 76606
rect 389173 76530 389239 76533
rect 215250 76528 389239 76530
rect 215250 76472 389178 76528
rect 389234 76472 389239 76528
rect 215250 76470 389239 76472
rect 151537 76467 151603 76470
rect 193121 76467 193187 76470
rect 209129 76467 209195 76470
rect 389173 76467 389239 76470
rect 154246 76332 154252 76396
rect 154316 76394 154322 76396
rect 154481 76394 154547 76397
rect 154316 76392 154547 76394
rect 154316 76336 154486 76392
rect 154542 76336 154547 76392
rect 154316 76334 154547 76336
rect 154316 76332 154322 76334
rect 154481 76331 154547 76334
rect 169017 76394 169083 76397
rect 191598 76394 191604 76396
rect 169017 76392 191604 76394
rect 169017 76336 169022 76392
rect 169078 76336 191604 76392
rect 169017 76334 191604 76336
rect 169017 76331 169083 76334
rect 191598 76332 191604 76334
rect 191668 76332 191674 76396
rect 174629 76258 174695 76261
rect 174854 76258 174860 76260
rect 174629 76256 174860 76258
rect 174629 76200 174634 76256
rect 174690 76200 174860 76256
rect 174629 76198 174860 76200
rect 174629 76195 174695 76198
rect 174854 76196 174860 76198
rect 174924 76196 174930 76260
rect 187693 76258 187759 76261
rect 187918 76258 187924 76260
rect 187693 76256 187924 76258
rect 187693 76200 187698 76256
rect 187754 76200 187924 76256
rect 187693 76198 187924 76200
rect 187693 76195 187759 76198
rect 187918 76196 187924 76198
rect 187988 76196 187994 76260
rect 153878 76060 153884 76124
rect 153948 76122 153954 76124
rect 217133 76122 217199 76125
rect 153948 76120 217199 76122
rect 153948 76064 217138 76120
rect 217194 76064 217199 76120
rect 153948 76062 217199 76064
rect 153948 76060 153954 76062
rect 217133 76059 217199 76062
rect 170622 75924 170628 75988
rect 170692 75986 170698 75988
rect 170949 75986 171015 75989
rect 170692 75984 171015 75986
rect 170692 75928 170954 75984
rect 171010 75928 171015 75984
rect 170692 75926 171015 75928
rect 170692 75924 170698 75926
rect 170949 75923 171015 75926
rect 119654 75788 119660 75852
rect 119724 75850 119730 75852
rect 132033 75850 132099 75853
rect 119724 75848 132099 75850
rect 119724 75792 132038 75848
rect 132094 75792 132099 75848
rect 119724 75790 132099 75792
rect 119724 75788 119730 75790
rect 132033 75787 132099 75790
rect 173249 75850 173315 75853
rect 207657 75850 207723 75853
rect 208209 75850 208275 75853
rect 173249 75848 208275 75850
rect 173249 75792 173254 75848
rect 173310 75792 207662 75848
rect 207718 75792 208214 75848
rect 208270 75792 208275 75848
rect 173249 75790 208275 75792
rect 173249 75787 173315 75790
rect 207657 75787 207723 75790
rect 208209 75787 208275 75790
rect 156781 75716 156847 75717
rect 113030 75652 113036 75716
rect 113100 75714 113106 75716
rect 147438 75714 147444 75716
rect 113100 75654 147444 75714
rect 113100 75652 113106 75654
rect 147438 75652 147444 75654
rect 147508 75652 147514 75716
rect 156781 75714 156828 75716
rect 156736 75712 156828 75714
rect 156736 75656 156786 75712
rect 156736 75654 156828 75656
rect 156781 75652 156828 75654
rect 156892 75652 156898 75716
rect 180057 75714 180123 75717
rect 206553 75714 206619 75717
rect 206921 75714 206987 75717
rect 180057 75712 206987 75714
rect 180057 75656 180062 75712
rect 180118 75656 206558 75712
rect 206614 75656 206926 75712
rect 206982 75656 206987 75712
rect 180057 75654 206987 75656
rect 156781 75651 156847 75652
rect 180057 75651 180123 75654
rect 206553 75651 206619 75654
rect 206921 75651 206987 75654
rect 122414 75516 122420 75580
rect 122484 75578 122490 75580
rect 154113 75578 154179 75581
rect 122484 75576 154179 75578
rect 122484 75520 154118 75576
rect 154174 75520 154179 75576
rect 122484 75518 154179 75520
rect 122484 75516 122490 75518
rect 154113 75515 154179 75518
rect 171685 75578 171751 75581
rect 171685 75576 205650 75578
rect 171685 75520 171690 75576
rect 171746 75520 205650 75576
rect 171685 75518 205650 75520
rect 171685 75515 171751 75518
rect 115749 75442 115815 75445
rect 145598 75442 145604 75444
rect 115749 75440 145604 75442
rect 115749 75384 115754 75440
rect 115810 75384 145604 75440
rect 115749 75382 145604 75384
rect 115749 75379 115815 75382
rect 145598 75380 145604 75382
rect 145668 75380 145674 75444
rect 173433 75442 173499 75445
rect 173709 75442 173775 75445
rect 173433 75440 173775 75442
rect 173433 75384 173438 75440
rect 173494 75384 173714 75440
rect 173770 75384 173775 75440
rect 173433 75382 173775 75384
rect 173433 75379 173499 75382
rect 173709 75379 173775 75382
rect 174537 75442 174603 75445
rect 174905 75442 174971 75445
rect 202086 75442 202092 75444
rect 174537 75440 202092 75442
rect 174537 75384 174542 75440
rect 174598 75384 174910 75440
rect 174966 75384 202092 75440
rect 174537 75382 202092 75384
rect 174537 75379 174603 75382
rect 174905 75379 174971 75382
rect 202086 75380 202092 75382
rect 202156 75380 202162 75444
rect 205590 75442 205650 75518
rect 206185 75442 206251 75445
rect 482277 75442 482343 75445
rect 205590 75440 482343 75442
rect 205590 75384 206190 75440
rect 206246 75384 482282 75440
rect 482338 75384 482343 75440
rect 205590 75382 482343 75384
rect 206185 75379 206251 75382
rect 482277 75379 482343 75382
rect 112437 75306 112503 75309
rect 112662 75306 112668 75308
rect 112437 75304 112668 75306
rect 112437 75248 112442 75304
rect 112498 75248 112668 75304
rect 112437 75246 112668 75248
rect 112437 75243 112503 75246
rect 112662 75244 112668 75246
rect 112732 75244 112738 75308
rect 116945 75306 117011 75309
rect 130469 75306 130535 75309
rect 130929 75306 130995 75309
rect 116945 75304 130995 75306
rect 116945 75248 116950 75304
rect 117006 75248 130474 75304
rect 130530 75248 130934 75304
rect 130990 75248 130995 75304
rect 116945 75246 130995 75248
rect 116945 75243 117011 75246
rect 130469 75243 130535 75246
rect 130929 75243 130995 75246
rect 156597 75306 156663 75309
rect 157190 75306 157196 75308
rect 156597 75304 157196 75306
rect 156597 75248 156602 75304
rect 156658 75248 157196 75304
rect 156597 75246 157196 75248
rect 156597 75243 156663 75246
rect 157190 75244 157196 75246
rect 157260 75244 157266 75308
rect 159030 75244 159036 75308
rect 159100 75306 159106 75308
rect 159541 75306 159607 75309
rect 159100 75304 159607 75306
rect 159100 75248 159546 75304
rect 159602 75248 159607 75304
rect 159100 75246 159607 75248
rect 159100 75244 159106 75246
rect 159541 75243 159607 75246
rect 168925 75306 168991 75309
rect 185894 75306 185900 75308
rect 168925 75304 185900 75306
rect 168925 75248 168930 75304
rect 168986 75248 185900 75304
rect 168925 75246 185900 75248
rect 168925 75243 168991 75246
rect 185894 75244 185900 75246
rect 185964 75244 185970 75308
rect 206921 75306 206987 75309
rect 509877 75306 509943 75309
rect 206921 75304 509943 75306
rect 206921 75248 206926 75304
rect 206982 75248 509882 75304
rect 509938 75248 509943 75304
rect 206921 75246 509943 75248
rect 206921 75243 206987 75246
rect 509877 75243 509943 75246
rect 7557 75170 7623 75173
rect 119654 75170 119660 75172
rect 7557 75168 119660 75170
rect 7557 75112 7562 75168
rect 7618 75112 119660 75168
rect 7557 75110 119660 75112
rect 7557 75107 7623 75110
rect 119654 75108 119660 75110
rect 119724 75108 119730 75172
rect 128997 75170 129063 75173
rect 129917 75170 129983 75173
rect 128997 75168 129983 75170
rect 128997 75112 129002 75168
rect 129058 75112 129922 75168
rect 129978 75112 129983 75168
rect 128997 75110 129983 75112
rect 128997 75107 129063 75110
rect 129917 75107 129983 75110
rect 172145 75170 172211 75173
rect 186998 75170 187004 75172
rect 172145 75168 187004 75170
rect 172145 75112 172150 75168
rect 172206 75112 187004 75168
rect 172145 75110 187004 75112
rect 172145 75107 172211 75110
rect 186998 75108 187004 75110
rect 187068 75108 187074 75172
rect 208209 75170 208275 75173
rect 524413 75170 524479 75173
rect 208209 75168 524479 75170
rect 208209 75112 208214 75168
rect 208270 75112 524418 75168
rect 524474 75112 524479 75168
rect 208209 75110 524479 75112
rect 208209 75107 208275 75110
rect 524413 75107 524479 75110
rect 125542 74972 125548 75036
rect 125612 75034 125618 75036
rect 144177 75034 144243 75037
rect 125612 75032 144243 75034
rect 125612 74976 144182 75032
rect 144238 74976 144243 75032
rect 125612 74974 144243 74976
rect 125612 74972 125618 74974
rect 144177 74971 144243 74974
rect 170070 74972 170076 75036
rect 170140 75034 170146 75036
rect 180701 75034 180767 75037
rect 170140 75032 180767 75034
rect 170140 74976 180706 75032
rect 180762 74976 180767 75032
rect 170140 74974 180767 74976
rect 170140 74972 170146 74974
rect 180701 74971 180767 74974
rect 120625 74626 120691 74629
rect 122782 74626 122788 74628
rect 120625 74624 122788 74626
rect 120625 74568 120630 74624
rect 120686 74568 122788 74624
rect 120625 74566 122788 74568
rect 120625 74563 120691 74566
rect 122782 74564 122788 74566
rect 122852 74564 122858 74628
rect 117078 74428 117084 74492
rect 117148 74490 117154 74492
rect 151721 74490 151787 74493
rect 117148 74488 151787 74490
rect 117148 74432 151726 74488
rect 151782 74432 151787 74488
rect 117148 74430 151787 74432
rect 117148 74428 117154 74430
rect 151721 74427 151787 74430
rect 185894 74428 185900 74492
rect 185964 74490 185970 74492
rect 186221 74490 186287 74493
rect 185964 74488 186287 74490
rect 185964 74432 186226 74488
rect 186282 74432 186287 74488
rect 185964 74430 186287 74432
rect 185964 74428 185970 74430
rect 186221 74427 186287 74430
rect 113582 74292 113588 74356
rect 113652 74354 113658 74356
rect 148542 74354 148548 74356
rect 113652 74294 148548 74354
rect 113652 74292 113658 74294
rect 148542 74292 148548 74294
rect 148612 74354 148618 74356
rect 154389 74354 154455 74357
rect 218421 74354 218487 74357
rect 148612 74294 149346 74354
rect 148612 74292 148618 74294
rect 100385 74218 100451 74221
rect 134374 74218 134380 74220
rect 100385 74216 134380 74218
rect 100385 74160 100390 74216
rect 100446 74160 134380 74216
rect 100385 74158 134380 74160
rect 100385 74155 100451 74158
rect 134374 74156 134380 74158
rect 134444 74156 134450 74220
rect 106774 74082 106780 74084
rect 103470 74022 106780 74082
rect 54477 73946 54543 73949
rect 103470 73946 103530 74022
rect 106774 74020 106780 74022
rect 106844 74082 106850 74084
rect 107193 74082 107259 74085
rect 106844 74080 107259 74082
rect 106844 74024 107198 74080
rect 107254 74024 107259 74080
rect 106844 74022 107259 74024
rect 106844 74020 106850 74022
rect 107193 74019 107259 74022
rect 122598 74020 122604 74084
rect 122668 74082 122674 74084
rect 149145 74082 149211 74085
rect 122668 74080 149211 74082
rect 122668 74024 149150 74080
rect 149206 74024 149211 74080
rect 122668 74022 149211 74024
rect 149286 74082 149346 74294
rect 154389 74352 218487 74354
rect 154389 74296 154394 74352
rect 154450 74296 218426 74352
rect 218482 74296 218487 74352
rect 154389 74294 218487 74296
rect 154389 74291 154455 74294
rect 218421 74291 218487 74294
rect 149462 74156 149468 74220
rect 149532 74218 149538 74220
rect 211613 74218 211679 74221
rect 149532 74216 211679 74218
rect 149532 74160 211618 74216
rect 211674 74160 211679 74216
rect 149532 74158 211679 74160
rect 149532 74156 149538 74158
rect 211613 74155 211679 74158
rect 218237 74082 218303 74085
rect 218513 74082 218579 74085
rect 237373 74082 237439 74085
rect 149286 74022 157350 74082
rect 122668 74020 122674 74022
rect 149145 74019 149211 74022
rect 54477 73944 103530 73946
rect 54477 73888 54482 73944
rect 54538 73888 103530 73944
rect 54477 73886 103530 73888
rect 54477 73883 54543 73886
rect 118550 73884 118556 73948
rect 118620 73946 118626 73948
rect 151169 73946 151235 73949
rect 118620 73944 151235 73946
rect 118620 73888 151174 73944
rect 151230 73888 151235 73944
rect 118620 73886 151235 73888
rect 118620 73884 118626 73886
rect 151169 73883 151235 73886
rect 22737 73810 22803 73813
rect 100385 73810 100451 73813
rect 22737 73808 100451 73810
rect 22737 73752 22742 73808
rect 22798 73752 100390 73808
rect 100446 73752 100451 73808
rect 22737 73750 100451 73752
rect 157290 73810 157350 74022
rect 218237 74080 237439 74082
rect 218237 74024 218242 74080
rect 218298 74024 218518 74080
rect 218574 74024 237378 74080
rect 237434 74024 237439 74080
rect 218237 74022 237439 74024
rect 218237 74019 218303 74022
rect 218513 74019 218579 74022
rect 237373 74019 237439 74022
rect 172329 73946 172395 73949
rect 197854 73946 197860 73948
rect 172329 73944 197860 73946
rect 172329 73888 172334 73944
rect 172390 73888 197860 73944
rect 172329 73886 197860 73888
rect 172329 73883 172395 73886
rect 197854 73884 197860 73886
rect 197924 73884 197930 73948
rect 218421 73946 218487 73949
rect 284293 73946 284359 73949
rect 218421 73944 284359 73946
rect 218421 73888 218426 73944
rect 218482 73888 284298 73944
rect 284354 73888 284359 73944
rect 218421 73886 284359 73888
rect 218421 73883 218487 73886
rect 284293 73883 284359 73886
rect 181529 73810 181595 73813
rect 157290 73808 181595 73810
rect 157290 73752 181534 73808
rect 181590 73752 181595 73808
rect 157290 73750 181595 73752
rect 22737 73747 22803 73750
rect 100385 73747 100451 73750
rect 181529 73747 181595 73750
rect 187969 73810 188035 73813
rect 269113 73810 269179 73813
rect 187969 73808 269179 73810
rect 187969 73752 187974 73808
rect 188030 73752 269118 73808
rect 269174 73752 269179 73808
rect 187969 73750 269179 73752
rect 187969 73747 188035 73750
rect 269113 73747 269179 73750
rect 173525 73674 173591 73677
rect 196014 73674 196020 73676
rect 173525 73672 196020 73674
rect 173525 73616 173530 73672
rect 173586 73616 196020 73672
rect 173525 73614 196020 73616
rect 173525 73611 173591 73614
rect 196014 73612 196020 73614
rect 196084 73612 196090 73676
rect 153469 73538 153535 73541
rect 187969 73538 188035 73541
rect 153469 73536 188035 73538
rect 153469 73480 153474 73536
rect 153530 73480 187974 73536
rect 188030 73480 188035 73536
rect 153469 73478 188035 73480
rect 153469 73475 153535 73478
rect 187969 73475 188035 73478
rect 151670 73340 151676 73404
rect 151740 73402 151746 73404
rect 218237 73402 218303 73405
rect 151740 73400 218303 73402
rect 151740 73344 218242 73400
rect 218298 73344 218303 73400
rect 151740 73342 218303 73344
rect 151740 73340 151746 73342
rect 218237 73339 218303 73342
rect 111425 73130 111491 73133
rect 145414 73130 145420 73132
rect 111425 73128 145420 73130
rect 111425 73072 111430 73128
rect 111486 73072 145420 73128
rect 111425 73070 145420 73072
rect 111425 73067 111491 73070
rect 145414 73068 145420 73070
rect 145484 73068 145490 73132
rect 169477 73130 169543 73133
rect 203425 73130 203491 73133
rect 169477 73128 203491 73130
rect 169477 73072 169482 73128
rect 169538 73072 203430 73128
rect 203486 73072 203491 73128
rect 169477 73070 203491 73072
rect 169477 73067 169543 73070
rect 203425 73067 203491 73070
rect 115841 72994 115907 72997
rect 146518 72994 146524 72996
rect 115841 72992 146524 72994
rect 115841 72936 115846 72992
rect 115902 72936 146524 72992
rect 115841 72934 146524 72936
rect 115841 72931 115907 72934
rect 146518 72932 146524 72934
rect 146588 72932 146594 72996
rect 170949 72994 171015 72997
rect 204529 72994 204595 72997
rect 170949 72992 204595 72994
rect 170949 72936 170954 72992
rect 171010 72936 204534 72992
rect 204590 72936 204595 72992
rect 170949 72934 204595 72936
rect 170949 72931 171015 72934
rect 204529 72931 204595 72934
rect 579613 72994 579679 72997
rect 583520 72994 584960 73084
rect 579613 72992 584960 72994
rect 579613 72936 579618 72992
rect 579674 72936 584960 72992
rect 579613 72934 584960 72936
rect 579613 72931 579679 72934
rect 116669 72858 116735 72861
rect 147070 72858 147076 72860
rect 116669 72856 147076 72858
rect 116669 72800 116674 72856
rect 116730 72800 147076 72856
rect 116669 72798 147076 72800
rect 116669 72795 116735 72798
rect 147070 72796 147076 72798
rect 147140 72796 147146 72860
rect 174997 72858 175063 72861
rect 175181 72858 175247 72861
rect 206277 72858 206343 72861
rect 174997 72856 206343 72858
rect 174997 72800 175002 72856
rect 175058 72800 175186 72856
rect 175242 72800 206282 72856
rect 206338 72800 206343 72856
rect 583520 72844 584960 72934
rect 174997 72798 206343 72800
rect 174997 72795 175063 72798
rect 175181 72795 175247 72798
rect 206277 72795 206343 72798
rect 119889 72722 119955 72725
rect 148358 72722 148364 72724
rect 119889 72720 148364 72722
rect 119889 72664 119894 72720
rect 119950 72664 148364 72720
rect 119889 72662 148364 72664
rect 119889 72659 119955 72662
rect 148358 72660 148364 72662
rect 148428 72660 148434 72724
rect 205766 72722 205772 72724
rect 176610 72662 205772 72722
rect 176193 72586 176259 72589
rect 176377 72586 176443 72589
rect 176610 72586 176670 72662
rect 205766 72660 205772 72662
rect 205836 72660 205842 72724
rect 176193 72584 176670 72586
rect 176193 72528 176198 72584
rect 176254 72528 176382 72584
rect 176438 72528 176670 72584
rect 176193 72526 176670 72528
rect 176193 72523 176259 72526
rect 176377 72523 176443 72526
rect 188286 72388 188292 72452
rect 188356 72450 188362 72452
rect 460933 72450 460999 72453
rect 188356 72448 460999 72450
rect 188356 72392 460938 72448
rect 460994 72392 460999 72448
rect 188356 72390 460999 72392
rect 188356 72388 188362 72390
rect 460933 72387 460999 72390
rect -960 71634 480 71724
rect 116158 71708 116164 71772
rect 116228 71770 116234 71772
rect 151169 71770 151235 71773
rect 151353 71770 151419 71773
rect 116228 71768 151419 71770
rect 116228 71712 151174 71768
rect 151230 71712 151358 71768
rect 151414 71712 151419 71768
rect 116228 71710 151419 71712
rect 116228 71708 116234 71710
rect 151169 71707 151235 71710
rect 151353 71707 151419 71710
rect 174721 71770 174787 71773
rect 212993 71770 213059 71773
rect 174721 71768 215310 71770
rect 174721 71712 174726 71768
rect 174782 71712 212998 71768
rect 213054 71712 215310 71768
rect 174721 71710 215310 71712
rect 174721 71707 174787 71710
rect 212993 71707 213059 71710
rect 3509 71634 3575 71637
rect -960 71632 3575 71634
rect -960 71576 3514 71632
rect 3570 71576 3575 71632
rect -960 71574 3575 71576
rect -960 71484 480 71574
rect 3509 71571 3575 71574
rect 115422 71572 115428 71636
rect 115492 71634 115498 71636
rect 150341 71634 150407 71637
rect 115492 71632 150407 71634
rect 115492 71576 150346 71632
rect 150402 71576 150407 71632
rect 115492 71574 150407 71576
rect 115492 71572 115498 71574
rect 150341 71571 150407 71574
rect 173341 71634 173407 71637
rect 205081 71634 205147 71637
rect 173341 71632 205147 71634
rect 173341 71576 173346 71632
rect 173402 71576 205086 71632
rect 205142 71576 205147 71632
rect 173341 71574 205147 71576
rect 173341 71571 173407 71574
rect 205081 71571 205147 71574
rect 122046 71436 122052 71500
rect 122116 71498 122122 71500
rect 155493 71498 155559 71501
rect 122116 71496 155559 71498
rect 122116 71440 155498 71496
rect 155554 71440 155559 71496
rect 122116 71438 155559 71440
rect 122116 71436 122122 71438
rect 155493 71435 155559 71438
rect 174445 71498 174511 71501
rect 215250 71498 215310 71710
rect 478137 71498 478203 71501
rect 174445 71496 200130 71498
rect 174445 71440 174450 71496
rect 174506 71440 200130 71496
rect 174445 71438 200130 71440
rect 215250 71496 478203 71498
rect 215250 71440 478142 71496
rect 478198 71440 478203 71496
rect 215250 71438 478203 71440
rect 174445 71435 174511 71438
rect 119521 71362 119587 71365
rect 146886 71362 146892 71364
rect 119521 71360 146892 71362
rect 119521 71304 119526 71360
rect 119582 71304 146892 71360
rect 119521 71302 146892 71304
rect 119521 71299 119587 71302
rect 146886 71300 146892 71302
rect 146956 71300 146962 71364
rect 161289 71362 161355 71365
rect 184054 71362 184060 71364
rect 161289 71360 184060 71362
rect 161289 71304 161294 71360
rect 161350 71304 184060 71360
rect 161289 71302 184060 71304
rect 161289 71299 161355 71302
rect 184054 71300 184060 71302
rect 184124 71300 184130 71364
rect 200070 71362 200130 71438
rect 478137 71435 478203 71438
rect 200982 71362 200988 71364
rect 200070 71302 200988 71362
rect 200982 71300 200988 71302
rect 201052 71362 201058 71364
rect 498837 71362 498903 71365
rect 201052 71360 498903 71362
rect 201052 71304 498842 71360
rect 498898 71304 498903 71360
rect 201052 71302 498903 71304
rect 201052 71300 201058 71302
rect 498837 71299 498903 71302
rect 122598 71164 122604 71228
rect 122668 71226 122674 71228
rect 149513 71226 149579 71229
rect 122668 71224 149579 71226
rect 122668 71168 149518 71224
rect 149574 71168 149579 71224
rect 122668 71166 149579 71168
rect 122668 71164 122674 71166
rect 149513 71163 149579 71166
rect 205081 71226 205147 71229
rect 531313 71226 531379 71229
rect 205081 71224 531379 71226
rect 205081 71168 205086 71224
rect 205142 71168 531318 71224
rect 531374 71168 531379 71224
rect 205081 71166 531379 71168
rect 205081 71163 205147 71166
rect 531313 71163 531379 71166
rect 17217 71090 17283 71093
rect 106958 71090 106964 71092
rect 17217 71088 106964 71090
rect 17217 71032 17222 71088
rect 17278 71032 106964 71088
rect 17217 71030 106964 71032
rect 17217 71027 17283 71030
rect 106958 71028 106964 71030
rect 107028 71090 107034 71092
rect 107377 71090 107443 71093
rect 107028 71088 107443 71090
rect 107028 71032 107382 71088
rect 107438 71032 107443 71088
rect 107028 71030 107443 71032
rect 107028 71028 107034 71030
rect 107377 71027 107443 71030
rect 187601 71090 187667 71093
rect 548517 71090 548583 71093
rect 187601 71088 548583 71090
rect 187601 71032 187606 71088
rect 187662 71032 548522 71088
rect 548578 71032 548583 71088
rect 187601 71030 548583 71032
rect 187601 71027 187667 71030
rect 548517 71027 548583 71030
rect 153009 70546 153075 70549
rect 142110 70544 153075 70546
rect 142110 70488 153014 70544
rect 153070 70488 153075 70544
rect 142110 70486 153075 70488
rect 117814 70212 117820 70276
rect 117884 70274 117890 70276
rect 142110 70274 142170 70486
rect 153009 70483 153075 70486
rect 205909 70274 205975 70277
rect 117884 70214 142170 70274
rect 174678 70272 205975 70274
rect 174678 70216 205914 70272
rect 205970 70216 205975 70272
rect 174678 70214 205975 70216
rect 117884 70212 117890 70214
rect 113950 70076 113956 70140
rect 114020 70138 114026 70140
rect 148869 70138 148935 70141
rect 114020 70136 148935 70138
rect 114020 70080 148874 70136
rect 148930 70080 148935 70136
rect 114020 70078 148935 70080
rect 114020 70076 114026 70078
rect 148869 70075 148935 70078
rect 120758 69940 120764 70004
rect 120828 70002 120834 70004
rect 153653 70002 153719 70005
rect 154021 70002 154087 70005
rect 120828 70000 154087 70002
rect 120828 69944 153658 70000
rect 153714 69944 154026 70000
rect 154082 69944 154087 70000
rect 120828 69942 154087 69944
rect 120828 69940 120834 69942
rect 153653 69939 153719 69942
rect 154021 69939 154087 69942
rect 171501 70002 171567 70005
rect 172145 70002 172211 70005
rect 174678 70002 174738 70214
rect 205909 70211 205975 70214
rect 206001 70138 206067 70141
rect 171501 70000 174738 70002
rect 171501 69944 171506 70000
rect 171562 69944 172150 70000
rect 172206 69944 174738 70000
rect 171501 69942 174738 69944
rect 174862 70136 206067 70138
rect 174862 70080 206006 70136
rect 206062 70080 206067 70136
rect 174862 70078 206067 70080
rect 171501 69939 171567 69942
rect 172145 69939 172211 69942
rect 122230 69804 122236 69868
rect 122300 69866 122306 69868
rect 152825 69866 152891 69869
rect 122300 69864 152891 69866
rect 122300 69808 152830 69864
rect 152886 69808 152891 69864
rect 122300 69806 152891 69808
rect 122300 69804 122306 69806
rect 152825 69803 152891 69806
rect 171685 69866 171751 69869
rect 172237 69866 172303 69869
rect 174862 69866 174922 70078
rect 206001 70075 206067 70078
rect 175917 70002 175983 70005
rect 208669 70002 208735 70005
rect 175917 70000 209790 70002
rect 175917 69944 175922 70000
rect 175978 69944 208674 70000
rect 208730 69944 209790 70000
rect 175917 69942 209790 69944
rect 175917 69939 175983 69942
rect 208669 69939 208735 69942
rect 171685 69864 174922 69866
rect 171685 69808 171690 69864
rect 171746 69808 172242 69864
rect 172298 69808 174922 69864
rect 171685 69806 174922 69808
rect 171685 69803 171751 69806
rect 172237 69803 172303 69806
rect 117681 69730 117747 69733
rect 147806 69730 147812 69732
rect 117681 69728 147812 69730
rect 117681 69672 117686 69728
rect 117742 69672 147812 69728
rect 117681 69670 147812 69672
rect 117681 69667 117747 69670
rect 147806 69668 147812 69670
rect 147876 69730 147882 69732
rect 148358 69730 148364 69732
rect 147876 69670 148364 69730
rect 147876 69668 147882 69670
rect 148358 69668 148364 69670
rect 148428 69668 148434 69732
rect 209730 69594 209790 69942
rect 557533 69594 557599 69597
rect 209730 69592 557599 69594
rect 209730 69536 557538 69592
rect 557594 69536 557599 69592
rect 209730 69534 557599 69536
rect 557533 69531 557599 69534
rect 148501 69458 148567 69461
rect 148869 69458 148935 69461
rect 148501 69456 148935 69458
rect 148501 69400 148506 69456
rect 148562 69400 148874 69456
rect 148930 69400 148935 69456
rect 148501 69398 148935 69400
rect 148501 69395 148567 69398
rect 148869 69395 148935 69398
rect 103053 68916 103119 68917
rect 103053 68912 103100 68916
rect 103164 68914 103170 68916
rect 103053 68856 103058 68912
rect 103053 68852 103100 68856
rect 103164 68854 103210 68914
rect 103164 68852 103170 68854
rect 117998 68852 118004 68916
rect 118068 68914 118074 68916
rect 151997 68914 152063 68917
rect 152733 68914 152799 68917
rect 118068 68912 152799 68914
rect 118068 68856 152002 68912
rect 152058 68856 152738 68912
rect 152794 68856 152799 68912
rect 118068 68854 152799 68856
rect 118068 68852 118074 68854
rect 103053 68851 103119 68852
rect 151997 68851 152063 68854
rect 152733 68851 152799 68854
rect 160093 68914 160159 68917
rect 161013 68914 161079 68917
rect 160093 68912 161490 68914
rect 160093 68856 160098 68912
rect 160154 68856 161018 68912
rect 161074 68856 161490 68912
rect 160093 68854 161490 68856
rect 160093 68851 160159 68854
rect 161013 68851 161079 68854
rect 118182 68716 118188 68780
rect 118252 68778 118258 68780
rect 142705 68778 142771 68781
rect 118252 68776 142771 68778
rect 118252 68720 142710 68776
rect 142766 68720 142771 68776
rect 118252 68718 142771 68720
rect 161430 68778 161490 68854
rect 187918 68852 187924 68916
rect 187988 68914 187994 68916
rect 188429 68914 188495 68917
rect 187988 68912 188495 68914
rect 187988 68856 188434 68912
rect 188490 68856 188495 68912
rect 187988 68854 188495 68856
rect 187988 68852 187994 68854
rect 188429 68851 188495 68854
rect 189073 68914 189139 68917
rect 200757 68916 200823 68917
rect 189574 68914 189580 68916
rect 189073 68912 189580 68914
rect 189073 68856 189078 68912
rect 189134 68856 189580 68912
rect 189073 68854 189580 68856
rect 189073 68851 189139 68854
rect 189574 68852 189580 68854
rect 189644 68852 189650 68916
rect 200757 68912 200804 68916
rect 200868 68914 200874 68916
rect 200757 68856 200762 68912
rect 200757 68852 200804 68856
rect 200868 68854 200914 68914
rect 200868 68852 200874 68854
rect 200757 68851 200823 68852
rect 181294 68778 181300 68780
rect 161430 68718 181300 68778
rect 118252 68716 118258 68718
rect 142705 68715 142771 68718
rect 181294 68716 181300 68718
rect 181364 68716 181370 68780
rect 116342 68580 116348 68644
rect 116412 68642 116418 68644
rect 151169 68642 151235 68645
rect 116412 68640 151235 68642
rect 116412 68584 151174 68640
rect 151230 68584 151235 68640
rect 116412 68582 151235 68584
rect 116412 68580 116418 68582
rect 151169 68579 151235 68582
rect 114093 68506 114159 68509
rect 144126 68506 144132 68508
rect 114093 68504 144132 68506
rect 114093 68448 114098 68504
rect 114154 68448 144132 68504
rect 114093 68446 144132 68448
rect 114093 68443 114159 68446
rect 144126 68444 144132 68446
rect 144196 68444 144202 68508
rect 149646 68444 149652 68508
rect 149716 68506 149722 68508
rect 215569 68506 215635 68509
rect 220813 68506 220879 68509
rect 149716 68504 220879 68506
rect 149716 68448 215574 68504
rect 215630 68448 220818 68504
rect 220874 68448 220879 68504
rect 149716 68446 220879 68448
rect 149716 68444 149722 68446
rect 215569 68443 215635 68446
rect 220813 68443 220879 68446
rect 26233 68370 26299 68373
rect 102133 68370 102199 68373
rect 26233 68368 102199 68370
rect 26233 68312 26238 68368
rect 26294 68312 102138 68368
rect 102194 68312 102199 68368
rect 26233 68310 102199 68312
rect 26233 68307 26299 68310
rect 102133 68307 102199 68310
rect 147438 68308 147444 68372
rect 147508 68370 147514 68372
rect 182817 68370 182883 68373
rect 147508 68368 182883 68370
rect 147508 68312 182822 68368
rect 182878 68312 182883 68368
rect 147508 68310 182883 68312
rect 147508 68308 147514 68310
rect 182817 68307 182883 68310
rect 18597 68234 18663 68237
rect 102225 68234 102291 68237
rect 102910 68234 102916 68236
rect 18597 68232 102916 68234
rect 18597 68176 18602 68232
rect 18658 68176 102230 68232
rect 102286 68176 102916 68232
rect 18597 68174 102916 68176
rect 18597 68171 18663 68174
rect 102225 68171 102291 68174
rect 102910 68172 102916 68174
rect 102980 68172 102986 68236
rect 146518 68172 146524 68236
rect 146588 68234 146594 68236
rect 195973 68234 196039 68237
rect 146588 68232 196039 68234
rect 146588 68176 195978 68232
rect 196034 68176 196039 68232
rect 146588 68174 196039 68176
rect 146588 68172 146594 68174
rect 195973 68171 196039 68174
rect 142705 68098 142771 68101
rect 153377 68098 153443 68101
rect 153929 68098 153995 68101
rect 142705 68096 153995 68098
rect 142705 68040 142710 68096
rect 142766 68040 153382 68096
rect 153438 68040 153934 68096
rect 153990 68040 153995 68096
rect 142705 68038 153995 68040
rect 142705 68035 142771 68038
rect 153377 68035 153443 68038
rect 153929 68035 153995 68038
rect 145598 67628 145604 67692
rect 145668 67690 145674 67692
rect 147121 67690 147187 67693
rect 145668 67688 147187 67690
rect 145668 67632 147126 67688
rect 147182 67632 147187 67688
rect 145668 67630 147187 67632
rect 145668 67628 145674 67630
rect 147121 67627 147187 67630
rect 110137 67554 110203 67557
rect 144310 67554 144316 67556
rect 110137 67552 144316 67554
rect 110137 67496 110142 67552
rect 110198 67496 144316 67552
rect 110137 67494 144316 67496
rect 110137 67491 110203 67494
rect 144310 67492 144316 67494
rect 144380 67554 144386 67556
rect 149697 67554 149763 67557
rect 144380 67552 149763 67554
rect 144380 67496 149702 67552
rect 149758 67496 149763 67552
rect 144380 67494 149763 67496
rect 144380 67492 144386 67494
rect 149697 67491 149763 67494
rect 149830 67492 149836 67556
rect 149900 67554 149906 67556
rect 215753 67554 215819 67557
rect 227713 67554 227779 67557
rect 149900 67552 227779 67554
rect 149900 67496 215758 67552
rect 215814 67496 227718 67552
rect 227774 67496 227779 67552
rect 149900 67494 227779 67496
rect 149900 67492 149906 67494
rect 215753 67491 215819 67494
rect 227713 67491 227779 67494
rect 113398 67356 113404 67420
rect 113468 67418 113474 67420
rect 114134 67418 114140 67420
rect 113468 67358 114140 67418
rect 113468 67356 113474 67358
rect 114134 67356 114140 67358
rect 114204 67356 114210 67420
rect 115606 67356 115612 67420
rect 115676 67418 115682 67420
rect 147990 67418 147996 67420
rect 115676 67358 147996 67418
rect 115676 67356 115682 67358
rect 147990 67356 147996 67358
rect 148060 67356 148066 67420
rect 170622 67356 170628 67420
rect 170692 67418 170698 67420
rect 170692 67358 200130 67418
rect 170692 67356 170698 67358
rect 114142 67282 114202 67356
rect 140814 67282 140820 67284
rect 114142 67222 140820 67282
rect 140814 67220 140820 67222
rect 140884 67220 140890 67284
rect 84193 67010 84259 67013
rect 108297 67010 108363 67013
rect 108430 67010 108436 67012
rect 84193 67008 108436 67010
rect 84193 66952 84198 67008
rect 84254 66952 108302 67008
rect 108358 66952 108436 67008
rect 84193 66950 108436 66952
rect 84193 66947 84259 66950
rect 108297 66947 108363 66950
rect 108430 66948 108436 66950
rect 108500 66948 108506 67012
rect 40033 66874 40099 66877
rect 104014 66874 104020 66876
rect 40033 66872 104020 66874
rect 40033 66816 40038 66872
rect 40094 66816 104020 66872
rect 40033 66814 104020 66816
rect 40033 66811 40099 66814
rect 104014 66812 104020 66814
rect 104084 66874 104090 66876
rect 104525 66874 104591 66877
rect 104084 66872 104591 66874
rect 104084 66816 104530 66872
rect 104586 66816 104591 66872
rect 104084 66814 104591 66816
rect 200070 66874 200130 67358
rect 212809 66874 212875 66877
rect 494053 66874 494119 66877
rect 200070 66872 494119 66874
rect 200070 66816 212814 66872
rect 212870 66816 494058 66872
rect 494114 66816 494119 66872
rect 200070 66814 494119 66816
rect 104084 66812 104090 66814
rect 104525 66811 104591 66814
rect 212809 66811 212875 66814
rect 494053 66811 494119 66814
rect 106917 66194 106983 66197
rect 108246 66194 108252 66196
rect 106917 66192 108252 66194
rect 106917 66136 106922 66192
rect 106978 66136 108252 66192
rect 106917 66134 108252 66136
rect 106917 66131 106983 66134
rect 108246 66132 108252 66134
rect 108316 66194 108322 66196
rect 108941 66194 109007 66197
rect 108316 66192 109007 66194
rect 108316 66136 108946 66192
rect 109002 66136 109007 66192
rect 108316 66134 109007 66136
rect 108316 66132 108322 66134
rect 108941 66131 109007 66134
rect 124070 66132 124076 66196
rect 124140 66194 124146 66196
rect 154849 66194 154915 66197
rect 124140 66192 154915 66194
rect 124140 66136 154854 66192
rect 154910 66136 154915 66192
rect 124140 66134 154915 66136
rect 124140 66132 124146 66134
rect 154849 66131 154915 66134
rect 170806 66132 170812 66196
rect 170876 66194 170882 66196
rect 204345 66194 204411 66197
rect 204713 66194 204779 66197
rect 170876 66192 204779 66194
rect 170876 66136 204350 66192
rect 204406 66136 204718 66192
rect 204774 66136 204779 66192
rect 170876 66134 204779 66136
rect 170876 66132 170882 66134
rect 204345 66131 204411 66134
rect 204713 66131 204779 66134
rect 109534 65996 109540 66060
rect 109604 66058 109610 66060
rect 138105 66058 138171 66061
rect 138473 66058 138539 66061
rect 203609 66060 203675 66061
rect 203558 66058 203564 66060
rect 109604 66056 138539 66058
rect 109604 66000 138110 66056
rect 138166 66000 138478 66056
rect 138534 66000 138539 66056
rect 109604 65998 138539 66000
rect 203518 65998 203564 66058
rect 203628 66056 203675 66060
rect 203670 66000 203675 66056
rect 109604 65996 109610 65998
rect 138105 65995 138171 65998
rect 138473 65995 138539 65998
rect 203558 65996 203564 65998
rect 203628 65996 203675 66000
rect 203609 65995 203675 65996
rect 110822 65922 110828 65924
rect 103470 65862 110828 65922
rect 93117 65514 93183 65517
rect 103470 65514 103530 65862
rect 110822 65860 110828 65862
rect 110892 65922 110898 65924
rect 139894 65922 139900 65924
rect 110892 65862 139900 65922
rect 110892 65860 110898 65862
rect 139894 65860 139900 65862
rect 139964 65860 139970 65924
rect 108798 65724 108804 65788
rect 108868 65786 108874 65788
rect 136909 65786 136975 65789
rect 108868 65784 136975 65786
rect 108868 65728 136914 65784
rect 136970 65728 136975 65784
rect 108868 65726 136975 65728
rect 108868 65724 108874 65726
rect 136909 65723 136975 65726
rect 112846 65588 112852 65652
rect 112916 65650 112922 65652
rect 139577 65650 139643 65653
rect 140221 65650 140287 65653
rect 112916 65648 140287 65650
rect 112916 65592 139582 65648
rect 139638 65592 140226 65648
rect 140282 65592 140287 65648
rect 112916 65590 140287 65592
rect 112916 65588 112922 65590
rect 139577 65587 139643 65590
rect 140221 65587 140287 65590
rect 93117 65512 103530 65514
rect 93117 65456 93122 65512
rect 93178 65456 103530 65512
rect 93117 65454 103530 65456
rect 204713 65514 204779 65517
rect 486417 65514 486483 65517
rect 204713 65512 486483 65514
rect 204713 65456 204718 65512
rect 204774 65456 486422 65512
rect 486478 65456 486483 65512
rect 204713 65454 486483 65456
rect 93117 65451 93183 65454
rect 204713 65451 204779 65454
rect 486417 65451 486483 65454
rect 135662 64834 135668 64836
rect 103470 64774 135668 64834
rect 101397 64698 101463 64701
rect 103470 64698 103530 64774
rect 135662 64772 135668 64774
rect 135732 64772 135738 64836
rect 143574 64772 143580 64836
rect 143644 64834 143650 64836
rect 144310 64834 144316 64836
rect 143644 64774 144316 64834
rect 143644 64772 143650 64774
rect 144310 64772 144316 64774
rect 144380 64772 144386 64836
rect 104249 64700 104315 64701
rect 104198 64698 104204 64700
rect 101397 64696 103530 64698
rect 101397 64640 101402 64696
rect 101458 64640 103530 64696
rect 101397 64638 103530 64640
rect 104158 64638 104204 64698
rect 104268 64696 104315 64700
rect 104310 64640 104315 64696
rect 101397 64635 101463 64638
rect 104198 64636 104204 64638
rect 104268 64636 104315 64640
rect 104249 64635 104315 64636
rect 110321 64698 110387 64701
rect 143758 64698 143764 64700
rect 110321 64696 143764 64698
rect 110321 64640 110326 64696
rect 110382 64640 143764 64696
rect 110321 64638 143764 64640
rect 110321 64635 110387 64638
rect 143758 64636 143764 64638
rect 143828 64698 143834 64700
rect 144494 64698 144500 64700
rect 143828 64638 144500 64698
rect 143828 64636 143834 64638
rect 144494 64636 144500 64638
rect 144564 64636 144570 64700
rect 174486 64636 174492 64700
rect 174556 64698 174562 64700
rect 200614 64698 200620 64700
rect 174556 64638 200620 64698
rect 174556 64636 174562 64638
rect 200614 64636 200620 64638
rect 200684 64698 200690 64700
rect 201350 64698 201356 64700
rect 200684 64638 201356 64698
rect 200684 64636 200690 64638
rect 201350 64636 201356 64638
rect 201420 64636 201426 64700
rect 111609 64562 111675 64565
rect 143574 64562 143580 64564
rect 111609 64560 143580 64562
rect 111609 64504 111614 64560
rect 111670 64504 143580 64560
rect 111609 64502 143580 64504
rect 111609 64499 111675 64502
rect 143574 64500 143580 64502
rect 143644 64500 143650 64564
rect 163129 64562 163195 64565
rect 187141 64564 187207 64565
rect 186078 64562 186084 64564
rect 163129 64560 186084 64562
rect 163129 64504 163134 64560
rect 163190 64504 186084 64560
rect 163129 64502 186084 64504
rect 163129 64499 163195 64502
rect 186078 64500 186084 64502
rect 186148 64500 186154 64564
rect 187141 64560 187188 64564
rect 187252 64562 187258 64564
rect 187141 64504 187146 64560
rect 187141 64500 187188 64504
rect 187252 64502 187298 64562
rect 187252 64500 187258 64502
rect 187141 64499 187207 64500
rect 156638 64364 156644 64428
rect 156708 64426 156714 64428
rect 156708 64366 200130 64426
rect 156708 64364 156714 64366
rect 57237 64290 57303 64293
rect 104249 64290 104315 64293
rect 57237 64288 104315 64290
rect 57237 64232 57242 64288
rect 57298 64232 104254 64288
rect 104310 64232 104315 64288
rect 57237 64230 104315 64232
rect 200070 64290 200130 64366
rect 213913 64290 213979 64293
rect 306373 64290 306439 64293
rect 200070 64288 306439 64290
rect 200070 64232 213918 64288
rect 213974 64232 306378 64288
rect 306434 64232 306439 64288
rect 200070 64230 306439 64232
rect 57237 64227 57303 64230
rect 104249 64227 104315 64230
rect 213913 64227 213979 64230
rect 306373 64227 306439 64230
rect 38653 64154 38719 64157
rect 101397 64154 101463 64157
rect 38653 64152 101463 64154
rect 38653 64096 38658 64152
rect 38714 64096 101402 64152
rect 101458 64096 101463 64152
rect 38653 64094 101463 64096
rect 38653 64091 38719 64094
rect 101397 64091 101463 64094
rect 201350 64092 201356 64156
rect 201420 64154 201426 64156
rect 543733 64154 543799 64157
rect 201420 64152 543799 64154
rect 201420 64096 543738 64152
rect 543794 64096 543799 64152
rect 201420 64094 543799 64096
rect 201420 64092 201426 64094
rect 543733 64091 543799 64094
rect 163129 63610 163195 63613
rect 163773 63610 163839 63613
rect 163129 63608 163839 63610
rect 163129 63552 163134 63608
rect 163190 63552 163778 63608
rect 163834 63552 163839 63608
rect 163129 63550 163839 63552
rect 163129 63547 163195 63550
rect 163773 63547 163839 63550
rect 105353 63474 105419 63477
rect 138606 63474 138612 63476
rect 84150 63472 138612 63474
rect 84150 63416 105358 63472
rect 105414 63416 138612 63472
rect 84150 63414 138612 63416
rect 81433 63066 81499 63069
rect 84150 63066 84210 63414
rect 105353 63411 105419 63414
rect 138606 63412 138612 63414
rect 138676 63412 138682 63476
rect 160686 63412 160692 63476
rect 160756 63474 160762 63476
rect 216765 63474 216831 63477
rect 160756 63472 219450 63474
rect 160756 63416 216770 63472
rect 216826 63416 219450 63472
rect 160756 63414 219450 63416
rect 160756 63412 160762 63414
rect 216765 63411 216831 63414
rect 100334 63276 100340 63340
rect 100404 63338 100410 63340
rect 133454 63338 133460 63340
rect 100404 63278 133460 63338
rect 100404 63276 100410 63278
rect 133454 63276 133460 63278
rect 133524 63276 133530 63340
rect 174670 63276 174676 63340
rect 174740 63338 174746 63340
rect 215477 63338 215543 63341
rect 174740 63336 215543 63338
rect 174740 63280 215482 63336
rect 215538 63280 215543 63336
rect 174740 63278 215543 63280
rect 174740 63276 174746 63278
rect 215477 63275 215543 63278
rect 107469 63202 107535 63205
rect 138422 63202 138428 63204
rect 81433 63064 84210 63066
rect 81433 63008 81438 63064
rect 81494 63008 84210 63064
rect 81433 63006 84210 63008
rect 103470 63200 138428 63202
rect 103470 63144 107474 63200
rect 107530 63144 138428 63200
rect 103470 63142 138428 63144
rect 81433 63003 81499 63006
rect 75177 62930 75243 62933
rect 103470 62930 103530 63142
rect 107469 63139 107535 63142
rect 138422 63140 138428 63142
rect 138492 63140 138498 63204
rect 75177 62928 103530 62930
rect 75177 62872 75182 62928
rect 75238 62872 103530 62928
rect 75177 62870 103530 62872
rect 219390 62930 219450 63414
rect 372613 62930 372679 62933
rect 219390 62928 372679 62930
rect 219390 62872 372618 62928
rect 372674 62872 372679 62928
rect 219390 62870 372679 62872
rect 75177 62867 75243 62870
rect 372613 62867 372679 62870
rect 2865 62794 2931 62797
rect 100334 62794 100340 62796
rect 2865 62792 100340 62794
rect 2865 62736 2870 62792
rect 2926 62736 100340 62792
rect 2865 62734 100340 62736
rect 2865 62731 2931 62734
rect 100334 62732 100340 62734
rect 100404 62732 100410 62796
rect 148542 62732 148548 62796
rect 148612 62794 148618 62796
rect 213913 62794 213979 62797
rect 148612 62792 213979 62794
rect 148612 62736 213918 62792
rect 213974 62736 213979 62792
rect 148612 62734 213979 62736
rect 148612 62732 148618 62734
rect 213913 62731 213979 62734
rect 215477 62794 215543 62797
rect 540237 62794 540303 62797
rect 215477 62792 540303 62794
rect 215477 62736 215482 62792
rect 215538 62736 540242 62792
rect 540298 62736 540303 62792
rect 215477 62734 540303 62736
rect 215477 62731 215543 62734
rect 540237 62731 540303 62734
rect 102685 62116 102751 62117
rect 102685 62112 102732 62116
rect 102796 62114 102802 62116
rect 106089 62114 106155 62117
rect 139710 62114 139716 62116
rect 102685 62056 102690 62112
rect 102685 62052 102732 62056
rect 102796 62054 102842 62114
rect 103470 62112 139716 62114
rect 103470 62056 106094 62112
rect 106150 62056 139716 62112
rect 103470 62054 139716 62056
rect 102796 62052 102802 62054
rect 102685 62051 102751 62052
rect 93945 61570 94011 61573
rect 103470 61570 103530 62054
rect 106089 62051 106155 62054
rect 139710 62052 139716 62054
rect 139780 62052 139786 62116
rect 173566 62052 173572 62116
rect 173636 62114 173642 62116
rect 212717 62114 212783 62117
rect 213821 62114 213887 62117
rect 173636 62112 213887 62114
rect 173636 62056 212722 62112
rect 212778 62056 213826 62112
rect 213882 62056 213887 62112
rect 173636 62054 213887 62056
rect 173636 62052 173642 62054
rect 212717 62051 212783 62054
rect 213821 62051 213887 62054
rect 199101 61978 199167 61981
rect 199326 61978 199332 61980
rect 199101 61976 199332 61978
rect 199101 61920 199106 61976
rect 199162 61920 199332 61976
rect 199101 61918 199332 61920
rect 199101 61915 199167 61918
rect 199326 61916 199332 61918
rect 199396 61916 199402 61980
rect 93945 61568 103530 61570
rect 93945 61512 93950 61568
rect 94006 61512 103530 61568
rect 93945 61510 103530 61512
rect 93945 61507 94011 61510
rect 32397 61434 32463 61437
rect 102133 61434 102199 61437
rect 32397 61432 102199 61434
rect 32397 61376 32402 61432
rect 32458 61376 102138 61432
rect 102194 61376 102199 61432
rect 32397 61374 102199 61376
rect 32397 61371 32463 61374
rect 102133 61371 102199 61374
rect 213821 61434 213887 61437
rect 526437 61434 526503 61437
rect 213821 61432 526503 61434
rect 213821 61376 213826 61432
rect 213882 61376 526442 61432
rect 526498 61376 526503 61432
rect 213821 61374 526503 61376
rect 213821 61371 213887 61374
rect 526437 61371 526503 61374
rect 112253 60620 112319 60621
rect 112253 60616 112300 60620
rect 112364 60618 112370 60620
rect 112253 60560 112258 60616
rect 112253 60556 112300 60560
rect 112364 60558 112410 60618
rect 112364 60556 112370 60558
rect 163262 60556 163268 60620
rect 163332 60618 163338 60620
rect 215385 60618 215451 60621
rect 163332 60616 215451 60618
rect 163332 60560 215390 60616
rect 215446 60560 215451 60616
rect 163332 60558 215451 60560
rect 163332 60556 163338 60558
rect 112253 60555 112319 60556
rect 215385 60555 215451 60558
rect 150014 60420 150020 60484
rect 150084 60482 150090 60484
rect 187877 60482 187943 60485
rect 150084 60480 190470 60482
rect 150084 60424 187882 60480
rect 187938 60424 190470 60480
rect 150084 60422 190470 60424
rect 150084 60420 150090 60422
rect 187877 60419 187943 60422
rect 164918 60284 164924 60348
rect 164988 60346 164994 60348
rect 164988 60286 180810 60346
rect 164988 60284 164994 60286
rect 97993 59938 98059 59941
rect 111793 59938 111859 59941
rect 97993 59936 111859 59938
rect 97993 59880 97998 59936
rect 98054 59880 111798 59936
rect 111854 59880 111859 59936
rect 97993 59878 111859 59880
rect 180750 59938 180810 60286
rect 190410 60210 190470 60422
rect 231853 60210 231919 60213
rect 190410 60208 231919 60210
rect 190410 60152 231858 60208
rect 231914 60152 231919 60208
rect 190410 60150 231919 60152
rect 231853 60147 231919 60150
rect 215385 60074 215451 60077
rect 394693 60074 394759 60077
rect 215385 60072 394759 60074
rect 215385 60016 215390 60072
rect 215446 60016 394698 60072
rect 394754 60016 394759 60072
rect 215385 60014 394759 60016
rect 215385 60011 215451 60014
rect 394693 60011 394759 60014
rect 191782 59938 191788 59940
rect 180750 59878 191788 59938
rect 97993 59875 98059 59878
rect 111793 59875 111859 59878
rect 191782 59876 191788 59878
rect 191852 59938 191858 59940
rect 423765 59938 423831 59941
rect 191852 59936 423831 59938
rect 191852 59880 423770 59936
rect 423826 59880 423831 59936
rect 191852 59878 423831 59880
rect 191852 59876 191858 59878
rect 423765 59875 423831 59878
rect 580533 59666 580599 59669
rect 583520 59666 584960 59756
rect 580533 59664 584960 59666
rect 580533 59608 580538 59664
rect 580594 59608 584960 59664
rect 580533 59606 584960 59608
rect 580533 59603 580599 59606
rect 583520 59516 584960 59606
rect 104157 59258 104223 59261
rect 104382 59258 104388 59260
rect 104157 59256 104388 59258
rect 104157 59200 104162 59256
rect 104218 59200 104388 59256
rect 104157 59198 104388 59200
rect 104157 59195 104223 59198
rect 104382 59196 104388 59198
rect 104452 59196 104458 59260
rect 172094 59196 172100 59260
rect 172164 59258 172170 59260
rect 212625 59258 212691 59261
rect 213821 59258 213887 59261
rect 172164 59256 213887 59258
rect 172164 59200 212630 59256
rect 212686 59200 213826 59256
rect 213882 59200 213887 59256
rect 172164 59198 213887 59200
rect 172164 59196 172170 59198
rect 212625 59195 212691 59198
rect 213821 59195 213887 59198
rect -960 58578 480 58668
rect 3509 58578 3575 58581
rect -960 58576 3575 58578
rect -960 58520 3514 58576
rect 3570 58520 3575 58576
rect -960 58518 3575 58520
rect -960 58428 480 58518
rect 3509 58515 3575 58518
rect 49693 58578 49759 58581
rect 104157 58578 104223 58581
rect 49693 58576 104223 58578
rect 49693 58520 49698 58576
rect 49754 58520 104162 58576
rect 104218 58520 104223 58576
rect 49693 58518 104223 58520
rect 49693 58515 49759 58518
rect 104157 58515 104223 58518
rect 213821 58578 213887 58581
rect 514017 58578 514083 58581
rect 213821 58576 514083 58578
rect 213821 58520 213826 58576
rect 213882 58520 514022 58576
rect 514078 58520 514083 58576
rect 213821 58518 514083 58520
rect 213821 58515 213887 58518
rect 514017 58515 514083 58518
rect 103789 57898 103855 57901
rect 104709 57898 104775 57901
rect 138238 57898 138244 57900
rect 103789 57896 138244 57898
rect 103789 57840 103794 57896
rect 103850 57840 104714 57896
rect 104770 57840 138244 57896
rect 103789 57838 138244 57840
rect 103789 57835 103855 57838
rect 104709 57835 104775 57838
rect 138238 57836 138244 57838
rect 138308 57836 138314 57900
rect 152590 57836 152596 57900
rect 152660 57898 152666 57900
rect 214097 57898 214163 57901
rect 152660 57896 219450 57898
rect 152660 57840 214102 57896
rect 214158 57840 219450 57896
rect 152660 57838 219450 57840
rect 152660 57836 152666 57838
rect 214097 57835 214163 57838
rect 100753 57762 100819 57765
rect 101765 57762 101831 57765
rect 134190 57762 134196 57764
rect 100753 57760 134196 57762
rect 100753 57704 100758 57760
rect 100814 57704 101770 57760
rect 101826 57704 134196 57760
rect 100753 57702 134196 57704
rect 100753 57699 100819 57702
rect 101765 57699 101831 57702
rect 134190 57700 134196 57702
rect 134260 57700 134266 57764
rect 175958 57700 175964 57764
rect 176028 57762 176034 57764
rect 215293 57762 215359 57765
rect 176028 57760 215359 57762
rect 176028 57704 215298 57760
rect 215354 57704 215359 57760
rect 176028 57702 215359 57704
rect 176028 57700 176034 57702
rect 215293 57699 215359 57702
rect 169334 57564 169340 57628
rect 169404 57626 169410 57628
rect 203241 57626 203307 57629
rect 204161 57626 204227 57629
rect 169404 57624 204227 57626
rect 169404 57568 203246 57624
rect 203302 57568 204166 57624
rect 204222 57568 204227 57624
rect 169404 57566 204227 57568
rect 219390 57626 219450 57838
rect 263593 57626 263659 57629
rect 219390 57624 263659 57626
rect 219390 57568 263598 57624
rect 263654 57568 263659 57624
rect 219390 57566 263659 57568
rect 169404 57564 169410 57566
rect 203241 57563 203307 57566
rect 204161 57563 204227 57566
rect 263593 57563 263659 57566
rect 165102 57428 165108 57492
rect 165172 57490 165178 57492
rect 199653 57490 199719 57493
rect 414657 57490 414723 57493
rect 165172 57488 414723 57490
rect 165172 57432 199658 57488
rect 199714 57432 414662 57488
rect 414718 57432 414723 57488
rect 165172 57430 414723 57432
rect 165172 57428 165178 57430
rect 199653 57427 199719 57430
rect 414657 57427 414723 57430
rect 77293 57354 77359 57357
rect 103789 57354 103855 57357
rect 77293 57352 103855 57354
rect 77293 57296 77298 57352
rect 77354 57296 103794 57352
rect 103850 57296 103855 57352
rect 77293 57294 103855 57296
rect 77293 57291 77359 57294
rect 103789 57291 103855 57294
rect 196249 57354 196315 57357
rect 196566 57354 196572 57356
rect 196249 57352 196572 57354
rect 196249 57296 196254 57352
rect 196310 57296 196572 57352
rect 196249 57294 196572 57296
rect 196249 57291 196315 57294
rect 196566 57292 196572 57294
rect 196636 57292 196642 57356
rect 204161 57354 204227 57357
rect 473445 57354 473511 57357
rect 204161 57352 473511 57354
rect 204161 57296 204166 57352
rect 204222 57296 473450 57352
rect 473506 57296 473511 57352
rect 204161 57294 473511 57296
rect 204161 57291 204227 57294
rect 473445 57291 473511 57294
rect 25497 57218 25563 57221
rect 100753 57218 100819 57221
rect 25497 57216 100819 57218
rect 25497 57160 25502 57216
rect 25558 57160 100758 57216
rect 100814 57160 100819 57216
rect 25497 57158 100819 57160
rect 25497 57155 25563 57158
rect 100753 57155 100819 57158
rect 147070 57156 147076 57220
rect 147140 57218 147146 57220
rect 191925 57218 191991 57221
rect 147140 57216 191991 57218
rect 147140 57160 191930 57216
rect 191986 57160 191991 57216
rect 147140 57158 191991 57160
rect 147140 57156 147146 57158
rect 191925 57155 191991 57158
rect 215293 57218 215359 57221
rect 567837 57218 567903 57221
rect 215293 57216 567903 57218
rect 215293 57160 215298 57216
rect 215354 57160 567842 57216
rect 567898 57160 567903 57216
rect 215293 57158 567903 57160
rect 215293 57155 215359 57158
rect 567837 57155 567903 57158
rect 99414 56476 99420 56540
rect 99484 56538 99490 56540
rect 100518 56538 100524 56540
rect 99484 56478 100524 56538
rect 99484 56476 99490 56478
rect 100518 56476 100524 56478
rect 100588 56538 100594 56540
rect 133270 56538 133276 56540
rect 100588 56478 133276 56538
rect 100588 56476 100594 56478
rect 133270 56476 133276 56478
rect 133340 56476 133346 56540
rect 157926 56476 157932 56540
rect 157996 56538 158002 56540
rect 192753 56538 192819 56541
rect 193029 56538 193095 56541
rect 157996 56536 193095 56538
rect 157996 56480 192758 56536
rect 192814 56480 193034 56536
rect 193090 56480 193095 56536
rect 157996 56478 193095 56480
rect 157996 56476 158002 56478
rect 192753 56475 192819 56478
rect 193029 56475 193095 56478
rect 162342 56340 162348 56404
rect 162412 56402 162418 56404
rect 196249 56402 196315 56405
rect 162412 56400 196315 56402
rect 162412 56344 196254 56400
rect 196310 56344 196315 56400
rect 162412 56342 196315 56344
rect 162412 56340 162418 56342
rect 196249 56339 196315 56342
rect 154246 56204 154252 56268
rect 154316 56266 154322 56268
rect 187785 56266 187851 56269
rect 284385 56266 284451 56269
rect 154316 56264 284451 56266
rect 154316 56208 187790 56264
rect 187846 56208 284390 56264
rect 284446 56208 284451 56264
rect 154316 56206 284451 56208
rect 154316 56204 154322 56206
rect 187785 56203 187851 56206
rect 284385 56203 284451 56206
rect 193029 56130 193095 56133
rect 331213 56130 331279 56133
rect 193029 56128 331279 56130
rect 193029 56072 193034 56128
rect 193090 56072 331218 56128
rect 331274 56072 331279 56128
rect 193029 56070 331279 56072
rect 193029 56067 193095 56070
rect 331213 56067 331279 56070
rect 88333 55994 88399 55997
rect 113541 55994 113607 55997
rect 113766 55994 113772 55996
rect 88333 55992 113772 55994
rect 88333 55936 88338 55992
rect 88394 55936 113546 55992
rect 113602 55936 113772 55992
rect 88333 55934 113772 55936
rect 88333 55931 88399 55934
rect 113541 55931 113607 55934
rect 113766 55932 113772 55934
rect 113836 55932 113842 55996
rect 196249 55994 196315 55997
rect 382917 55994 382983 55997
rect 196249 55992 382983 55994
rect 196249 55936 196254 55992
rect 196310 55936 382922 55992
rect 382978 55936 382983 55992
rect 196249 55934 382983 55936
rect 196249 55931 196315 55934
rect 382917 55931 382983 55934
rect 12433 55858 12499 55861
rect 99414 55858 99420 55860
rect 12433 55856 99420 55858
rect 12433 55800 12438 55856
rect 12494 55800 99420 55856
rect 12433 55798 99420 55800
rect 12433 55795 12499 55798
rect 99414 55796 99420 55798
rect 99484 55796 99490 55860
rect 171910 55796 171916 55860
rect 171980 55858 171986 55860
rect 205725 55858 205791 55861
rect 499573 55858 499639 55861
rect 171980 55856 499639 55858
rect 171980 55800 205730 55856
rect 205786 55800 499578 55856
rect 499634 55800 499639 55856
rect 171980 55798 499639 55800
rect 171980 55796 171986 55798
rect 205725 55795 205791 55798
rect 499573 55795 499639 55798
rect 107561 55178 107627 55181
rect 139526 55178 139532 55180
rect 107561 55176 139532 55178
rect 107561 55120 107566 55176
rect 107622 55120 139532 55176
rect 107561 55118 139532 55120
rect 107561 55115 107627 55118
rect 139526 55116 139532 55118
rect 139596 55116 139602 55180
rect 166390 55116 166396 55180
rect 166460 55178 166466 55180
rect 200205 55178 200271 55181
rect 201401 55178 201467 55181
rect 166460 55176 201467 55178
rect 166460 55120 200210 55176
rect 200266 55120 201406 55176
rect 201462 55120 201467 55176
rect 166460 55118 201467 55120
rect 166460 55116 166466 55118
rect 200205 55115 200271 55118
rect 201401 55115 201467 55118
rect 120441 55042 120507 55045
rect 139342 55042 139348 55044
rect 120441 55040 139348 55042
rect 120441 54984 120446 55040
rect 120502 54984 139348 55040
rect 120441 54982 139348 54984
rect 120441 54979 120507 54982
rect 139342 54980 139348 54982
rect 139412 54980 139418 55044
rect 160870 54980 160876 55044
rect 160940 55042 160946 55044
rect 160940 54982 180810 55042
rect 160940 54980 160946 54982
rect 102133 54634 102199 54637
rect 107561 54634 107627 54637
rect 102133 54632 107627 54634
rect 102133 54576 102138 54632
rect 102194 54576 107566 54632
rect 107622 54576 107627 54632
rect 102133 54574 107627 54576
rect 180750 54634 180810 54982
rect 203333 54772 203399 54773
rect 203333 54770 203380 54772
rect 203252 54768 203380 54770
rect 203444 54770 203450 54772
rect 203977 54770 204043 54773
rect 203444 54768 204043 54770
rect 203252 54712 203338 54768
rect 203444 54712 203982 54768
rect 204038 54712 204043 54768
rect 203252 54710 203380 54712
rect 203333 54708 203380 54710
rect 203444 54710 204043 54712
rect 203444 54708 203450 54710
rect 203333 54707 203399 54708
rect 203977 54707 204043 54710
rect 190821 54634 190887 54637
rect 369853 54634 369919 54637
rect 180750 54632 369919 54634
rect 180750 54576 190826 54632
rect 190882 54576 369858 54632
rect 369914 54576 369919 54632
rect 180750 54574 369919 54576
rect 102133 54571 102199 54574
rect 107561 54571 107627 54574
rect 190821 54571 190887 54574
rect 369853 54571 369919 54574
rect 92473 54498 92539 54501
rect 120441 54498 120507 54501
rect 92473 54496 120507 54498
rect 92473 54440 92478 54496
rect 92534 54440 120446 54496
rect 120502 54440 120507 54496
rect 92473 54438 120507 54440
rect 92473 54435 92539 54438
rect 120441 54435 120507 54438
rect 201401 54498 201467 54501
rect 440233 54498 440299 54501
rect 201401 54496 440299 54498
rect 201401 54440 201406 54496
rect 201462 54440 440238 54496
rect 440294 54440 440299 54496
rect 201401 54438 440299 54440
rect 201401 54435 201467 54438
rect 440233 54435 440299 54438
rect 105445 53818 105511 53821
rect 137502 53818 137508 53820
rect 105445 53816 137508 53818
rect 105445 53760 105450 53816
rect 105506 53760 137508 53816
rect 105445 53758 137508 53760
rect 105445 53755 105511 53758
rect 137502 53756 137508 53758
rect 137572 53756 137578 53820
rect 161054 53756 161060 53820
rect 161124 53818 161130 53820
rect 194542 53818 194548 53820
rect 161124 53758 194548 53818
rect 161124 53756 161130 53758
rect 194542 53756 194548 53758
rect 194612 53756 194618 53820
rect 158110 53620 158116 53684
rect 158180 53682 158186 53684
rect 190729 53682 190795 53685
rect 158180 53680 190795 53682
rect 158180 53624 190734 53680
rect 190790 53624 190795 53680
rect 158180 53622 190795 53624
rect 158180 53620 158186 53622
rect 190410 53274 190470 53622
rect 190729 53619 190795 53622
rect 333973 53274 334039 53277
rect 190410 53272 334039 53274
rect 190410 53216 333978 53272
rect 334034 53216 334039 53272
rect 190410 53214 334039 53216
rect 333973 53211 334039 53214
rect 56593 53138 56659 53141
rect 105445 53138 105511 53141
rect 56593 53136 105511 53138
rect 56593 53080 56598 53136
rect 56654 53080 105450 53136
rect 105506 53080 105511 53136
rect 56593 53078 105511 53080
rect 56593 53075 56659 53078
rect 105445 53075 105511 53078
rect 146886 53076 146892 53140
rect 146956 53138 146962 53140
rect 193305 53138 193371 53141
rect 146956 53136 193371 53138
rect 146956 53080 193310 53136
rect 193366 53080 193371 53136
rect 146956 53078 193371 53080
rect 146956 53076 146962 53078
rect 193305 53075 193371 53078
rect 194542 53076 194548 53140
rect 194612 53138 194618 53140
rect 364977 53138 365043 53141
rect 194612 53136 365043 53138
rect 194612 53080 364982 53136
rect 365038 53080 365043 53136
rect 194612 53078 365043 53080
rect 194612 53076 194618 53078
rect 364977 53075 365043 53078
rect 114134 52532 114140 52596
rect 114204 52594 114210 52596
rect 120073 52594 120139 52597
rect 114204 52592 120139 52594
rect 114204 52536 120078 52592
rect 120134 52536 120139 52592
rect 114204 52534 120139 52536
rect 114204 52532 114210 52534
rect 120073 52531 120139 52534
rect 99465 52458 99531 52461
rect 100569 52458 100635 52461
rect 193213 52460 193279 52461
rect 201953 52460 202019 52461
rect 133086 52458 133092 52460
rect 99465 52456 133092 52458
rect 99465 52400 99470 52456
rect 99526 52400 100574 52456
rect 100630 52400 133092 52456
rect 99465 52398 133092 52400
rect 99465 52395 99531 52398
rect 100569 52395 100635 52398
rect 133086 52396 133092 52398
rect 133156 52396 133162 52460
rect 193213 52456 193260 52460
rect 193324 52458 193330 52460
rect 201902 52458 201908 52460
rect 193213 52400 193218 52456
rect 193213 52396 193260 52400
rect 193324 52398 193370 52458
rect 201862 52398 201908 52458
rect 201972 52456 202019 52460
rect 202014 52400 202019 52456
rect 193324 52396 193330 52398
rect 201902 52396 201908 52398
rect 201972 52396 202019 52400
rect 193213 52395 193279 52396
rect 201953 52395 202019 52396
rect 156822 52260 156828 52324
rect 156892 52322 156898 52324
rect 190637 52322 190703 52325
rect 191741 52322 191807 52325
rect 156892 52320 191807 52322
rect 156892 52264 190642 52320
rect 190698 52264 191746 52320
rect 191802 52264 191807 52320
rect 156892 52262 191807 52264
rect 156892 52260 156898 52262
rect 190637 52259 190703 52262
rect 191741 52259 191807 52262
rect 174854 52124 174860 52188
rect 174924 52186 174930 52188
rect 208577 52186 208643 52189
rect 208761 52186 208827 52189
rect 174924 52184 208827 52186
rect 174924 52128 208582 52184
rect 208638 52128 208766 52184
rect 208822 52128 208827 52184
rect 174924 52126 208827 52128
rect 174924 52124 174930 52126
rect 208577 52123 208643 52126
rect 208761 52123 208827 52126
rect 152774 51988 152780 52052
rect 152844 52050 152850 52052
rect 214005 52050 214071 52053
rect 259453 52050 259519 52053
rect 152844 52048 259519 52050
rect 152844 51992 214010 52048
rect 214066 51992 259458 52048
rect 259514 51992 259519 52048
rect 152844 51990 259519 51992
rect 152844 51988 152850 51990
rect 214005 51987 214071 51990
rect 259453 51987 259519 51990
rect 191741 51914 191807 51917
rect 320173 51914 320239 51917
rect 191741 51912 320239 51914
rect 191741 51856 191746 51912
rect 191802 51856 320178 51912
rect 320234 51856 320239 51912
rect 191741 51854 320239 51856
rect 191741 51851 191807 51854
rect 320173 51851 320239 51854
rect 17953 51778 18019 51781
rect 99465 51778 99531 51781
rect 17953 51776 99531 51778
rect 17953 51720 17958 51776
rect 18014 51720 99470 51776
rect 99526 51720 99531 51776
rect 17953 51718 99531 51720
rect 17953 51715 18019 51718
rect 99465 51715 99531 51718
rect 208761 51778 208827 51781
rect 542353 51778 542419 51781
rect 208761 51776 542419 51778
rect 208761 51720 208766 51776
rect 208822 51720 542358 51776
rect 542414 51720 542419 51776
rect 208761 51718 542419 51720
rect 208761 51715 208827 51718
rect 542353 51715 542419 51718
rect 104801 50962 104867 50965
rect 138054 50962 138060 50964
rect 84150 50960 138060 50962
rect 84150 50904 104806 50960
rect 104862 50904 138060 50960
rect 84150 50902 138060 50904
rect 78673 50418 78739 50421
rect 84150 50418 84210 50902
rect 104801 50899 104867 50902
rect 138054 50900 138060 50902
rect 138124 50900 138130 50964
rect 207054 50900 207060 50964
rect 207124 50962 207130 50964
rect 207197 50962 207263 50965
rect 207124 50960 207263 50962
rect 207124 50904 207202 50960
rect 207258 50904 207263 50960
rect 207124 50902 207263 50904
rect 207124 50900 207130 50902
rect 207197 50899 207263 50902
rect 134006 50826 134012 50828
rect 78673 50416 84210 50418
rect 78673 50360 78678 50416
rect 78734 50360 84210 50416
rect 78673 50358 84210 50360
rect 103470 50766 134012 50826
rect 78673 50355 78739 50358
rect 27705 50282 27771 50285
rect 101857 50282 101923 50285
rect 103470 50282 103530 50766
rect 134006 50764 134012 50766
rect 134076 50764 134082 50828
rect 158294 50764 158300 50828
rect 158364 50826 158370 50828
rect 158364 50766 180810 50826
rect 158364 50764 158370 50766
rect 180750 50690 180810 50766
rect 192017 50690 192083 50693
rect 338113 50690 338179 50693
rect 180750 50688 338179 50690
rect 180750 50632 192022 50688
rect 192078 50632 338118 50688
rect 338174 50632 338179 50688
rect 180750 50630 338179 50632
rect 192017 50627 192083 50630
rect 338113 50627 338179 50630
rect 161238 50492 161244 50556
rect 161308 50554 161314 50556
rect 193990 50554 193996 50556
rect 161308 50494 193996 50554
rect 161308 50492 161314 50494
rect 193990 50492 193996 50494
rect 194060 50554 194066 50556
rect 373993 50554 374059 50557
rect 194060 50552 374059 50554
rect 194060 50496 373998 50552
rect 374054 50496 374059 50552
rect 194060 50494 374059 50496
rect 194060 50492 194066 50494
rect 373993 50491 374059 50494
rect 165286 50356 165292 50420
rect 165356 50418 165362 50420
rect 198825 50418 198891 50421
rect 418797 50418 418863 50421
rect 165356 50416 418863 50418
rect 165356 50360 198830 50416
rect 198886 50360 418802 50416
rect 418858 50360 418863 50416
rect 165356 50358 418863 50360
rect 165356 50356 165362 50358
rect 198825 50355 198891 50358
rect 418797 50355 418863 50358
rect 27705 50280 103530 50282
rect 27705 50224 27710 50280
rect 27766 50224 101862 50280
rect 101918 50224 103530 50280
rect 27705 50222 103530 50224
rect 27705 50219 27771 50222
rect 101857 50219 101923 50222
rect 176142 50220 176148 50284
rect 176212 50282 176218 50284
rect 209814 50282 209820 50284
rect 176212 50222 209820 50282
rect 176212 50220 176218 50222
rect 209814 50220 209820 50222
rect 209884 50282 209890 50284
rect 556153 50282 556219 50285
rect 209884 50280 556219 50282
rect 209884 50224 556158 50280
rect 556214 50224 556219 50280
rect 209884 50222 556219 50224
rect 209884 50220 209890 50222
rect 556153 50219 556219 50222
rect 99465 49602 99531 49605
rect 100661 49602 100727 49605
rect 133822 49602 133828 49604
rect 99465 49600 133828 49602
rect 99465 49544 99470 49600
rect 99526 49544 100666 49600
rect 100722 49544 133828 49600
rect 99465 49542 133828 49544
rect 99465 49539 99531 49542
rect 100661 49539 100727 49542
rect 133822 49540 133828 49542
rect 133892 49540 133898 49604
rect 162526 49540 162532 49604
rect 162596 49602 162602 49604
rect 196157 49602 196223 49605
rect 196709 49602 196775 49605
rect 162596 49600 196775 49602
rect 162596 49544 196162 49600
rect 196218 49544 196714 49600
rect 196770 49544 196775 49600
rect 162596 49542 196775 49544
rect 162596 49540 162602 49542
rect 196157 49539 196223 49542
rect 196709 49539 196775 49542
rect 176326 49404 176332 49468
rect 176396 49466 176402 49468
rect 204437 49466 204503 49469
rect 204713 49466 204779 49469
rect 176396 49464 204779 49466
rect 176396 49408 204442 49464
rect 204498 49408 204718 49464
rect 204774 49408 204779 49464
rect 176396 49406 204779 49408
rect 176396 49404 176402 49406
rect 204437 49403 204503 49406
rect 204713 49403 204779 49406
rect 196709 49058 196775 49061
rect 387793 49058 387859 49061
rect 196709 49056 387859 49058
rect 196709 49000 196714 49056
rect 196770 49000 387798 49056
rect 387854 49000 387859 49056
rect 196709 48998 387859 49000
rect 196709 48995 196775 48998
rect 387793 48995 387859 48998
rect 30373 48922 30439 48925
rect 99465 48922 99531 48925
rect 30373 48920 99531 48922
rect 30373 48864 30378 48920
rect 30434 48864 99470 48920
rect 99526 48864 99531 48920
rect 30373 48862 99531 48864
rect 30373 48859 30439 48862
rect 99465 48859 99531 48862
rect 204713 48922 204779 48925
rect 565813 48922 565879 48925
rect 204713 48920 565879 48922
rect 204713 48864 204718 48920
rect 204774 48864 565818 48920
rect 565874 48864 565879 48920
rect 204713 48862 565879 48864
rect 204713 48859 204779 48862
rect 565813 48859 565879 48862
rect 100753 48242 100819 48245
rect 101949 48242 102015 48245
rect 135478 48242 135484 48244
rect 100753 48240 135484 48242
rect 100753 48184 100758 48240
rect 100814 48184 101954 48240
rect 102010 48184 135484 48240
rect 100753 48182 135484 48184
rect 100753 48179 100819 48182
rect 101949 48179 102015 48182
rect 135478 48180 135484 48182
rect 135548 48180 135554 48244
rect 170990 48180 170996 48244
rect 171060 48242 171066 48244
rect 209865 48242 209931 48245
rect 211061 48242 211127 48245
rect 171060 48240 211127 48242
rect 171060 48184 209870 48240
rect 209926 48184 211066 48240
rect 211122 48184 211127 48240
rect 171060 48182 211127 48184
rect 171060 48180 171066 48182
rect 209865 48179 209931 48182
rect 211061 48179 211127 48182
rect 163446 48044 163452 48108
rect 163516 48106 163522 48108
rect 197445 48106 197511 48109
rect 198457 48106 198523 48109
rect 163516 48104 198523 48106
rect 163516 48048 197450 48104
rect 197506 48048 198462 48104
rect 198518 48048 198523 48104
rect 163516 48046 198523 48048
rect 163516 48044 163522 48046
rect 197445 48043 197511 48046
rect 198457 48043 198523 48046
rect 169518 47908 169524 47972
rect 169588 47970 169594 47972
rect 203149 47970 203215 47973
rect 204161 47970 204227 47973
rect 169588 47968 204227 47970
rect 169588 47912 203154 47968
rect 203210 47912 204166 47968
rect 204222 47912 204227 47968
rect 169588 47910 204227 47912
rect 169588 47908 169594 47910
rect 203149 47907 203215 47910
rect 204161 47907 204227 47910
rect 198457 47834 198523 47837
rect 405733 47834 405799 47837
rect 198457 47832 405799 47834
rect 198457 47776 198462 47832
rect 198518 47776 405738 47832
rect 405794 47776 405799 47832
rect 198457 47774 405799 47776
rect 198457 47771 198523 47774
rect 405733 47771 405799 47774
rect 204161 47698 204227 47701
rect 466453 47698 466519 47701
rect 204161 47696 466519 47698
rect 204161 47640 204166 47696
rect 204222 47640 466458 47696
rect 466514 47640 466519 47696
rect 204161 47638 466519 47640
rect 204161 47635 204227 47638
rect 466453 47635 466519 47638
rect 39297 47562 39363 47565
rect 100753 47562 100819 47565
rect 39297 47560 100819 47562
rect 39297 47504 39302 47560
rect 39358 47504 100758 47560
rect 100814 47504 100819 47560
rect 39297 47502 100819 47504
rect 39297 47499 39363 47502
rect 100753 47499 100819 47502
rect 211061 47562 211127 47565
rect 490005 47562 490071 47565
rect 211061 47560 490071 47562
rect 211061 47504 211066 47560
rect 211122 47504 490010 47560
rect 490066 47504 490071 47560
rect 211061 47502 490071 47504
rect 211061 47499 211127 47502
rect 490005 47499 490071 47502
rect 100753 46882 100819 46885
rect 102041 46882 102107 46885
rect 135294 46882 135300 46884
rect 100753 46880 135300 46882
rect 100753 46824 100758 46880
rect 100814 46824 102046 46880
rect 102102 46824 135300 46880
rect 100753 46822 135300 46824
rect 100753 46819 100819 46822
rect 102041 46819 102107 46822
rect 135294 46820 135300 46822
rect 135364 46820 135370 46884
rect 152406 46820 152412 46884
rect 152476 46882 152482 46884
rect 218053 46882 218119 46885
rect 152476 46880 219450 46882
rect 152476 46824 218058 46880
rect 218114 46824 219450 46880
rect 152476 46822 219450 46824
rect 152476 46820 152482 46822
rect 218053 46819 218119 46822
rect 167678 46684 167684 46748
rect 167748 46746 167754 46748
rect 207197 46746 207263 46749
rect 207606 46746 207612 46748
rect 167748 46686 200130 46746
rect 167748 46684 167754 46686
rect 167862 46548 167868 46612
rect 167932 46610 167938 46612
rect 167932 46550 180810 46610
rect 167932 46548 167938 46550
rect 44265 46202 44331 46205
rect 100753 46202 100819 46205
rect 44265 46200 100819 46202
rect 44265 46144 44270 46200
rect 44326 46144 100758 46200
rect 100814 46144 100819 46200
rect 44265 46142 100819 46144
rect 180750 46202 180810 46550
rect 200070 46338 200130 46686
rect 207197 46744 207612 46746
rect 207197 46688 207202 46744
rect 207258 46688 207612 46744
rect 207197 46686 207612 46688
rect 207197 46683 207263 46686
rect 207606 46684 207612 46686
rect 207676 46684 207682 46748
rect 219390 46474 219450 46822
rect 251173 46474 251239 46477
rect 219390 46472 251239 46474
rect 219390 46416 251178 46472
rect 251234 46416 251239 46472
rect 219390 46414 251239 46416
rect 251173 46411 251239 46414
rect 202045 46338 202111 46341
rect 454033 46338 454099 46341
rect 200070 46336 454099 46338
rect 200070 46280 202050 46336
rect 202106 46280 454038 46336
rect 454094 46280 454099 46336
rect 200070 46278 454099 46280
rect 202045 46275 202111 46278
rect 454033 46275 454099 46278
rect 580441 46338 580507 46341
rect 583520 46338 584960 46428
rect 580441 46336 584960 46338
rect 580441 46280 580446 46336
rect 580502 46280 584960 46336
rect 580441 46278 584960 46280
rect 580441 46275 580507 46278
rect 201718 46202 201724 46204
rect 180750 46142 201724 46202
rect 44265 46139 44331 46142
rect 100753 46139 100819 46142
rect 201718 46140 201724 46142
rect 201788 46202 201794 46204
rect 455413 46202 455479 46205
rect 201788 46200 455479 46202
rect 201788 46144 455418 46200
rect 455474 46144 455479 46200
rect 583520 46188 584960 46278
rect 201788 46142 455479 46144
rect 201788 46140 201794 46142
rect 455413 46139 455479 46142
rect -960 45522 480 45612
rect 207606 45596 207612 45660
rect 207676 45658 207682 45660
rect 207933 45658 207999 45661
rect 207676 45656 207999 45658
rect 207676 45600 207938 45656
rect 207994 45600 207999 45656
rect 207676 45598 207999 45600
rect 207676 45596 207682 45598
rect 207933 45595 207999 45598
rect -960 45462 674 45522
rect -960 45386 480 45462
rect 614 45386 674 45462
rect 175038 45460 175044 45524
rect 175108 45522 175114 45524
rect 208485 45522 208551 45525
rect 175108 45520 208551 45522
rect 175108 45464 208490 45520
rect 208546 45464 208551 45520
rect 175108 45462 208551 45464
rect 175108 45460 175114 45462
rect 208485 45459 208551 45462
rect -960 45372 674 45386
rect 246 45326 674 45372
rect 246 44842 306 45326
rect 148358 45324 148364 45388
rect 148428 45386 148434 45388
rect 209865 45386 209931 45389
rect 148428 45384 209931 45386
rect 148428 45328 209870 45384
rect 209926 45328 209931 45384
rect 148428 45326 209931 45328
rect 148428 45324 148434 45326
rect 209865 45323 209931 45326
rect 162158 45188 162164 45252
rect 162228 45250 162234 45252
rect 196065 45250 196131 45253
rect 390553 45250 390619 45253
rect 162228 45248 390619 45250
rect 162228 45192 196070 45248
rect 196126 45192 390558 45248
rect 390614 45192 390619 45248
rect 162228 45190 390619 45192
rect 162228 45188 162234 45190
rect 196065 45187 196131 45190
rect 390553 45187 390619 45190
rect 166574 45052 166580 45116
rect 166644 45114 166650 45116
rect 198774 45114 198780 45116
rect 166644 45054 198780 45114
rect 166644 45052 166650 45054
rect 198774 45052 198780 45054
rect 198844 45114 198850 45116
rect 444373 45114 444439 45117
rect 198844 45112 444439 45114
rect 198844 45056 444378 45112
rect 444434 45056 444439 45112
rect 198844 45054 444439 45056
rect 198844 45052 198850 45054
rect 444373 45051 444439 45054
rect 173750 44916 173756 44980
rect 173820 44978 173826 44980
rect 203006 44978 203012 44980
rect 173820 44918 203012 44978
rect 173820 44916 173826 44918
rect 203006 44916 203012 44918
rect 203076 44978 203082 44980
rect 520917 44978 520983 44981
rect 203076 44976 520983 44978
rect 203076 44920 520922 44976
rect 520978 44920 520983 44976
rect 203076 44918 520983 44920
rect 203076 44916 203082 44918
rect 520917 44915 520983 44918
rect 208485 44842 208551 44845
rect 535453 44842 535519 44845
rect 246 44782 6930 44842
rect 6870 44298 6930 44782
rect 208485 44840 535519 44842
rect 208485 44784 208490 44840
rect 208546 44784 535458 44840
rect 535514 44784 535519 44840
rect 208485 44782 535519 44784
rect 208485 44779 208551 44782
rect 535453 44779 535519 44782
rect 116526 44298 116532 44300
rect 6870 44238 116532 44298
rect 116526 44236 116532 44238
rect 116596 44236 116602 44300
rect 102225 44162 102291 44165
rect 102777 44162 102843 44165
rect 137686 44162 137692 44164
rect 102225 44160 137692 44162
rect 102225 44104 102230 44160
rect 102286 44104 102782 44160
rect 102838 44104 137692 44160
rect 102225 44102 137692 44104
rect 102225 44099 102291 44102
rect 102777 44099 102843 44102
rect 137686 44100 137692 44102
rect 137756 44100 137762 44164
rect 154430 44100 154436 44164
rect 154500 44162 154506 44164
rect 209313 44162 209379 44165
rect 154500 44160 209790 44162
rect 154500 44104 209318 44160
rect 209374 44104 209790 44160
rect 154500 44102 209790 44104
rect 154500 44100 154506 44102
rect 209313 44099 209379 44102
rect 166758 43964 166764 44028
rect 166828 44026 166834 44028
rect 200481 44026 200547 44029
rect 201401 44026 201467 44029
rect 166828 44024 201467 44026
rect 166828 43968 200486 44024
rect 200542 43968 201406 44024
rect 201462 43968 201467 44024
rect 166828 43966 201467 43968
rect 166828 43964 166834 43966
rect 200481 43963 200547 43966
rect 201401 43963 201467 43966
rect 163630 43828 163636 43892
rect 163700 43890 163706 43892
rect 197302 43890 197308 43892
rect 163700 43830 197308 43890
rect 163700 43828 163706 43830
rect 197302 43828 197308 43830
rect 197372 43890 197378 43892
rect 209730 43890 209790 44102
rect 276105 43890 276171 43893
rect 197372 43830 200130 43890
rect 209730 43888 276171 43890
rect 209730 43832 276110 43888
rect 276166 43832 276171 43888
rect 209730 43830 276171 43832
rect 197372 43828 197378 43830
rect 200070 43754 200130 43830
rect 276105 43827 276171 43830
rect 408493 43754 408559 43757
rect 200070 43752 408559 43754
rect 200070 43696 408498 43752
rect 408554 43696 408559 43752
rect 200070 43694 408559 43696
rect 408493 43691 408559 43694
rect 201401 43618 201467 43621
rect 427813 43618 427879 43621
rect 201401 43616 427879 43618
rect 201401 43560 201406 43616
rect 201462 43560 427818 43616
rect 427874 43560 427879 43616
rect 201401 43558 427879 43560
rect 201401 43555 201467 43558
rect 427813 43555 427879 43558
rect 63493 43482 63559 43485
rect 102225 43482 102291 43485
rect 63493 43480 102291 43482
rect 63493 43424 63498 43480
rect 63554 43424 102230 43480
rect 102286 43424 102291 43480
rect 63493 43422 102291 43424
rect 63493 43419 63559 43422
rect 102225 43419 102291 43422
rect 168046 43420 168052 43484
rect 168116 43482 168122 43484
rect 201534 43482 201540 43484
rect 168116 43422 201540 43482
rect 168116 43420 168122 43422
rect 201534 43420 201540 43422
rect 201604 43482 201610 43484
rect 458173 43482 458239 43485
rect 201604 43480 458239 43482
rect 201604 43424 458178 43480
rect 458234 43424 458239 43480
rect 201604 43422 458239 43424
rect 201604 43420 201610 43422
rect 458173 43419 458239 43422
rect 155534 38524 155540 38588
rect 155604 38586 155610 38588
rect 211153 38586 211219 38589
rect 212441 38586 212507 38589
rect 155604 38584 212507 38586
rect 155604 38528 211158 38584
rect 211214 38528 212446 38584
rect 212502 38528 212507 38584
rect 155604 38526 212507 38528
rect 155604 38524 155610 38526
rect 211153 38523 211219 38526
rect 212441 38523 212507 38526
rect 212441 37906 212507 37909
rect 293953 37906 294019 37909
rect 212441 37904 294019 37906
rect 212441 37848 212446 37904
rect 212502 37848 293958 37904
rect 294014 37848 294019 37904
rect 212441 37846 294019 37848
rect 212441 37843 212507 37846
rect 293953 37843 294019 37846
rect 176510 37164 176516 37228
rect 176580 37226 176586 37228
rect 216857 37226 216923 37229
rect 217225 37226 217291 37229
rect 176580 37224 217291 37226
rect 176580 37168 216862 37224
rect 216918 37168 217230 37224
rect 217286 37168 217291 37224
rect 176580 37166 217291 37168
rect 176580 37164 176586 37166
rect 216857 37163 216923 37166
rect 217225 37163 217291 37166
rect 157006 37028 157012 37092
rect 157076 37090 157082 37092
rect 157076 37030 180810 37090
rect 157076 37028 157082 37030
rect 180750 36682 180810 37030
rect 195421 36682 195487 36685
rect 307017 36682 307083 36685
rect 180750 36680 307083 36682
rect 180750 36624 195426 36680
rect 195482 36624 307022 36680
rect 307078 36624 307083 36680
rect 180750 36622 307083 36624
rect 195421 36619 195487 36622
rect 307017 36619 307083 36622
rect 217225 36546 217291 36549
rect 552013 36546 552079 36549
rect 217225 36544 552079 36546
rect 217225 36488 217230 36544
rect 217286 36488 552018 36544
rect 552074 36488 552079 36544
rect 217225 36486 552079 36488
rect 217225 36483 217291 36486
rect 552013 36483 552079 36486
rect 157190 35804 157196 35868
rect 157260 35866 157266 35868
rect 204253 35866 204319 35869
rect 157260 35864 204319 35866
rect 157260 35808 204258 35864
rect 204314 35808 204319 35864
rect 157260 35806 204319 35808
rect 157260 35804 157266 35806
rect 204253 35803 204319 35806
rect 144494 35124 144500 35188
rect 144564 35186 144570 35188
rect 156045 35186 156111 35189
rect 144564 35184 156111 35186
rect 144564 35128 156050 35184
rect 156106 35128 156111 35184
rect 144564 35126 156111 35128
rect 144564 35124 144570 35126
rect 156045 35123 156111 35126
rect 204253 35186 204319 35189
rect 311157 35186 311223 35189
rect 204253 35184 311223 35186
rect 204253 35128 204258 35184
rect 204314 35128 311162 35184
rect 311218 35128 311223 35184
rect 204253 35126 311223 35128
rect 204253 35123 204319 35126
rect 311157 35123 311223 35126
rect 151302 34444 151308 34508
rect 151372 34506 151378 34508
rect 189993 34506 190059 34509
rect 190361 34506 190427 34509
rect 151372 34504 190427 34506
rect 151372 34448 189998 34504
rect 190054 34448 190366 34504
rect 190422 34448 190427 34504
rect 151372 34446 190427 34448
rect 151372 34444 151378 34446
rect 189993 34443 190059 34446
rect 190361 34443 190427 34446
rect 189993 33826 190059 33829
rect 234705 33826 234771 33829
rect 189993 33824 234771 33826
rect 189993 33768 189998 33824
rect 190054 33768 234710 33824
rect 234766 33768 234771 33824
rect 189993 33766 234771 33768
rect 189993 33763 190059 33766
rect 234705 33763 234771 33766
rect 580349 33146 580415 33149
rect 583520 33146 584960 33236
rect 580349 33144 584960 33146
rect 580349 33088 580354 33144
rect 580410 33088 584960 33144
rect 580349 33086 584960 33088
rect 580349 33083 580415 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3509 32466 3575 32469
rect -960 32464 3575 32466
rect -960 32408 3514 32464
rect 3570 32408 3575 32464
rect -960 32406 3575 32408
rect -960 32316 480 32406
rect 3509 32403 3575 32406
rect 148174 30908 148180 30972
rect 148244 30970 148250 30972
rect 212625 30970 212691 30973
rect 148244 30968 212691 30970
rect 148244 30912 212630 30968
rect 212686 30912 212691 30968
rect 148244 30910 212691 30912
rect 148244 30908 148250 30910
rect 212625 30907 212691 30910
rect 165470 26148 165476 26212
rect 165540 26210 165546 26212
rect 205633 26210 205699 26213
rect 165540 26208 205699 26210
rect 165540 26152 205638 26208
rect 205694 26152 205699 26208
rect 165540 26150 205699 26152
rect 165540 26148 165546 26150
rect 205633 26147 205699 26150
rect 205633 25530 205699 25533
rect 418153 25530 418219 25533
rect 205633 25528 418219 25530
rect 205633 25472 205638 25528
rect 205694 25472 418158 25528
rect 418214 25472 418219 25528
rect 205633 25470 418219 25472
rect 205633 25467 205699 25470
rect 418153 25467 418219 25470
rect 145414 22612 145420 22676
rect 145484 22674 145490 22676
rect 171869 22674 171935 22677
rect 145484 22672 171935 22674
rect 145484 22616 171874 22672
rect 171930 22616 171935 22672
rect 145484 22614 171935 22616
rect 145484 22612 145490 22614
rect 171869 22611 171935 22614
rect 158478 21932 158484 21996
rect 158548 21994 158554 21996
rect 158548 21934 209790 21994
rect 158548 21932 158554 21934
rect 158846 21796 158852 21860
rect 158916 21858 158922 21860
rect 207013 21858 207079 21861
rect 158916 21856 207306 21858
rect 158916 21800 207018 21856
rect 207074 21800 207306 21856
rect 158916 21798 207306 21800
rect 158916 21796 158922 21798
rect 207013 21795 207079 21798
rect 159030 21660 159036 21724
rect 159100 21722 159106 21724
rect 159100 21662 200130 21722
rect 159100 21660 159106 21662
rect 200070 21314 200130 21662
rect 207246 21450 207306 21798
rect 209730 21586 209790 21934
rect 212533 21586 212599 21589
rect 336733 21586 336799 21589
rect 209730 21584 336799 21586
rect 209730 21528 212538 21584
rect 212594 21528 336738 21584
rect 336794 21528 336799 21584
rect 209730 21526 336799 21528
rect 212533 21523 212599 21526
rect 336733 21523 336799 21526
rect 350533 21450 350599 21453
rect 207246 21448 350599 21450
rect 207246 21392 350538 21448
rect 350594 21392 350599 21448
rect 207246 21390 350599 21392
rect 350533 21387 350599 21390
rect 207105 21314 207171 21317
rect 354673 21314 354739 21317
rect 200070 21312 354739 21314
rect 200070 21256 207110 21312
rect 207166 21256 354678 21312
rect 354734 21256 354739 21312
rect 200070 21254 354739 21256
rect 207105 21251 207171 21254
rect 354673 21251 354739 21254
rect 580165 19818 580231 19821
rect 583520 19818 584960 19908
rect 580165 19816 584960 19818
rect 580165 19760 580170 19816
rect 580226 19760 584960 19816
rect 580165 19758 584960 19760
rect 580165 19755 580231 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 155718 17852 155724 17916
rect 155788 17914 155794 17916
rect 209773 17914 209839 17917
rect 211061 17914 211127 17917
rect 155788 17912 211127 17914
rect 155788 17856 209778 17912
rect 209834 17856 211066 17912
rect 211122 17856 211127 17912
rect 155788 17854 211127 17856
rect 155788 17852 155794 17854
rect 209773 17851 209839 17854
rect 211061 17851 211127 17854
rect 211061 17234 211127 17237
rect 300853 17234 300919 17237
rect 211061 17232 300919 17234
rect 211061 17176 211066 17232
rect 211122 17176 300858 17232
rect 300914 17176 300919 17232
rect 211061 17174 300919 17176
rect 211061 17171 211127 17174
rect 300853 17171 300919 17174
rect 3417 10298 3483 10301
rect 111006 10298 111012 10300
rect 3417 10296 111012 10298
rect 3417 10240 3422 10296
rect 3478 10240 111012 10296
rect 3417 10238 111012 10240
rect 3417 10235 3483 10238
rect 111006 10236 111012 10238
rect 111076 10236 111082 10300
rect 144310 8876 144316 8940
rect 144380 8938 144386 8940
rect 160185 8938 160251 8941
rect 144380 8936 160251 8938
rect 144380 8880 160190 8936
rect 160246 8880 160251 8936
rect 144380 8878 160251 8880
rect 144380 8876 144386 8878
rect 160185 8875 160251 8878
rect 580257 6626 580323 6629
rect 583520 6626 584960 6716
rect 580257 6624 584960 6626
rect -960 6490 480 6580
rect 580257 6568 580262 6624
rect 580318 6568 584960 6624
rect 580257 6566 584960 6568
rect 580257 6563 580323 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 144126 6156 144132 6220
rect 144196 6218 144202 6220
rect 158897 6218 158963 6221
rect 144196 6216 158963 6218
rect 144196 6160 158902 6216
rect 158958 6160 158963 6216
rect 144196 6158 158963 6160
rect 144196 6156 144202 6158
rect 158897 6155 158963 6158
<< via3 >>
rect 187740 274620 187804 274684
rect 109540 265236 109604 265300
rect 197676 265236 197740 265300
rect 115796 265100 115860 265164
rect 198964 265100 199028 265164
rect 112852 264964 112916 265028
rect 197492 264964 197556 265028
rect 121132 263876 121196 263940
rect 121316 263740 121380 263804
rect 118372 263604 118436 263668
rect 114140 262788 114204 262852
rect 193628 262652 193692 262716
rect 111564 262516 111628 262580
rect 193444 262516 193508 262580
rect 189212 262304 189276 262308
rect 189212 262248 189262 262304
rect 189262 262248 189276 262304
rect 189212 262244 189276 262248
rect 111380 261156 111444 261220
rect 109356 261020 109420 261084
rect 111196 260884 111260 260948
rect 116900 259932 116964 259996
rect 116716 259524 116780 259588
rect 186084 259524 186148 259588
rect 186084 212468 186148 212532
rect 187188 212468 187252 212532
rect 132172 201180 132236 201244
rect 139900 201180 139964 201244
rect 131620 201044 131684 201108
rect 138796 201044 138860 201108
rect 117084 200772 117148 200836
rect 151492 200908 151556 200972
rect 131804 200772 131868 200836
rect 136588 200772 136652 200836
rect 153332 200636 153396 200700
rect 106780 200500 106844 200564
rect 140084 200500 140148 200564
rect 207060 200500 207124 200564
rect 122420 200364 122484 200428
rect 151676 200364 151740 200428
rect 122604 200228 122668 200292
rect 133460 199956 133524 200020
rect 140084 200092 140148 200156
rect 133644 199858 133648 199884
rect 133648 199858 133704 199884
rect 133704 199858 133708 199884
rect 133644 199820 133708 199858
rect 134196 199820 134260 199884
rect 135300 199820 135364 199884
rect 136404 199858 136408 199884
rect 136408 199858 136464 199884
rect 136464 199858 136468 199884
rect 136404 199820 136468 199858
rect 137140 199858 137144 199884
rect 137144 199858 137200 199884
rect 137200 199858 137204 199884
rect 137140 199820 137204 199858
rect 137508 199858 137512 199884
rect 137512 199858 137568 199884
rect 137568 199858 137572 199884
rect 137508 199820 137572 199858
rect 138060 199820 138124 199884
rect 138796 199858 138800 199884
rect 138800 199858 138856 199884
rect 138856 199858 138860 199884
rect 138796 199820 138860 199858
rect 139532 199858 139536 199884
rect 139536 199858 139592 199884
rect 139592 199858 139596 199884
rect 139532 199820 139596 199858
rect 139900 199858 139904 199884
rect 139904 199858 139960 199884
rect 139960 199858 139964 199884
rect 139900 199820 139964 199858
rect 141004 199820 141068 199884
rect 142292 199820 142356 199884
rect 141556 199684 141620 199748
rect 143028 199820 143092 199884
rect 131804 199608 131868 199612
rect 131804 199552 131818 199608
rect 131818 199552 131868 199608
rect 131804 199548 131868 199552
rect 141188 199548 141252 199612
rect 141924 199548 141988 199612
rect 142844 199548 142908 199612
rect 131620 199472 131684 199476
rect 131620 199416 131634 199472
rect 131634 199416 131684 199472
rect 131620 199412 131684 199416
rect 132172 199472 132236 199476
rect 132172 199416 132186 199472
rect 132186 199416 132236 199472
rect 132172 199412 132236 199416
rect 137140 199412 137204 199476
rect 142844 199412 142908 199476
rect 146708 199858 146712 199884
rect 146712 199858 146768 199884
rect 146768 199858 146772 199884
rect 146708 199820 146772 199858
rect 147260 199858 147264 199884
rect 147264 199858 147320 199884
rect 147320 199858 147324 199884
rect 147260 199820 147324 199858
rect 146524 199548 146588 199612
rect 148180 199820 148244 199884
rect 154804 200092 154868 200156
rect 151492 199880 151556 199884
rect 151492 199824 151496 199880
rect 151496 199824 151552 199880
rect 151552 199824 151556 199880
rect 151492 199820 151556 199824
rect 152964 199820 153028 199884
rect 153148 199820 153212 199884
rect 153516 199858 153520 199884
rect 153520 199858 153576 199884
rect 153576 199858 153580 199884
rect 153516 199820 153580 199858
rect 153884 199820 153948 199884
rect 155172 199820 155236 199884
rect 151676 199684 151740 199748
rect 153332 199548 153396 199612
rect 168420 200228 168484 200292
rect 166396 200092 166460 200156
rect 156644 199858 156648 199884
rect 156648 199858 156704 199884
rect 156704 199858 156708 199884
rect 156644 199820 156708 199858
rect 157748 199858 157752 199884
rect 157752 199858 157808 199884
rect 157808 199858 157812 199884
rect 157748 199820 157812 199858
rect 157196 199722 157200 199748
rect 157200 199722 157256 199748
rect 157256 199722 157260 199748
rect 157196 199684 157260 199722
rect 157564 199684 157628 199748
rect 154620 199472 154684 199476
rect 154620 199416 154634 199472
rect 154634 199416 154684 199472
rect 154620 199412 154684 199416
rect 118556 199276 118620 199340
rect 160140 199820 160204 199884
rect 161060 199820 161124 199884
rect 161244 199744 161308 199748
rect 161244 199688 161258 199744
rect 161258 199688 161308 199744
rect 161244 199684 161308 199688
rect 161428 199722 161478 199748
rect 161478 199722 161492 199748
rect 161428 199684 161492 199722
rect 161796 199820 161860 199884
rect 163084 199820 163148 199884
rect 163820 199820 163884 199884
rect 163452 199744 163516 199748
rect 163452 199688 163502 199744
rect 163502 199688 163516 199744
rect 163452 199684 163516 199688
rect 163636 199722 163640 199748
rect 163640 199722 163696 199748
rect 163696 199722 163700 199748
rect 163636 199684 163700 199722
rect 162532 199548 162596 199612
rect 163268 199548 163332 199612
rect 161244 199412 161308 199476
rect 163636 199472 163700 199476
rect 164924 199820 164988 199884
rect 165844 199820 165908 199884
rect 166028 199858 166032 199884
rect 166032 199858 166088 199884
rect 166088 199858 166092 199884
rect 166028 199820 166092 199858
rect 166580 199820 166644 199884
rect 167500 199820 167564 199884
rect 167684 199820 167748 199884
rect 164740 199684 164804 199748
rect 165292 199684 165356 199748
rect 168604 199820 168668 199884
rect 168788 199820 168852 199884
rect 169524 199956 169588 200020
rect 170812 199956 170876 200020
rect 163636 199416 163686 199472
rect 163686 199416 163700 199472
rect 163636 199412 163700 199416
rect 166396 199412 166460 199476
rect 168420 199608 168484 199612
rect 168420 199552 168470 199608
rect 168470 199552 168484 199608
rect 168420 199548 168484 199552
rect 169156 199608 169220 199612
rect 169892 199858 169896 199884
rect 169896 199858 169952 199884
rect 169952 199858 169956 199884
rect 169892 199820 169956 199858
rect 169156 199552 169170 199608
rect 169170 199552 169220 199608
rect 169156 199548 169220 199552
rect 170076 199684 170140 199748
rect 135484 199140 135548 199204
rect 136404 199200 136468 199204
rect 136404 199144 136418 199200
rect 136418 199144 136468 199200
rect 136404 199140 136468 199144
rect 136588 199140 136652 199204
rect 141924 198792 141988 198796
rect 141924 198736 141938 198792
rect 141938 198736 141988 198792
rect 141924 198732 141988 198736
rect 142660 198732 142724 198796
rect 143028 198792 143092 198796
rect 169340 199412 169404 199476
rect 169708 199412 169772 199476
rect 170628 199858 170632 199884
rect 170632 199858 170688 199884
rect 170688 199858 170692 199884
rect 170628 199820 170692 199858
rect 172836 199956 172900 200020
rect 174124 199956 174188 200020
rect 171364 199820 171428 199884
rect 171548 199820 171612 199884
rect 172468 199820 172532 199884
rect 172652 199858 172656 199884
rect 172656 199858 172712 199884
rect 172712 199858 172716 199884
rect 172652 199820 172716 199858
rect 173388 199820 173452 199884
rect 171732 199684 171796 199748
rect 171916 199684 171980 199748
rect 172468 199684 172532 199748
rect 172974 199684 173038 199748
rect 174860 199820 174924 199884
rect 175412 199820 175476 199884
rect 175964 199820 176028 199884
rect 176516 199820 176580 199884
rect 173572 199684 173636 199748
rect 174308 199684 174372 199748
rect 171732 199412 171796 199476
rect 168972 199276 169036 199340
rect 174860 199276 174924 199340
rect 200804 199140 200868 199204
rect 200620 199004 200684 199068
rect 174124 198928 174188 198932
rect 174124 198872 174174 198928
rect 174174 198872 174188 198928
rect 174124 198868 174188 198872
rect 174492 198868 174556 198932
rect 200988 198868 201052 198932
rect 143028 198736 143078 198792
rect 143078 198736 143092 198792
rect 143028 198732 143092 198736
rect 163268 198732 163332 198796
rect 189028 198732 189092 198796
rect 133644 198596 133708 198660
rect 134380 198596 134444 198660
rect 169156 198596 169220 198660
rect 171548 198596 171612 198660
rect 187924 198596 187988 198660
rect 138428 198460 138492 198524
rect 155172 198460 155236 198524
rect 175596 198460 175660 198524
rect 107516 198324 107580 198388
rect 161244 198324 161308 198388
rect 168604 198324 168668 198388
rect 201172 198324 201236 198388
rect 143580 198188 143644 198252
rect 148916 198188 148980 198252
rect 106964 198052 107028 198116
rect 141004 198112 141068 198116
rect 141004 198056 141018 198112
rect 141018 198056 141068 198112
rect 141004 198052 141068 198056
rect 148180 198052 148244 198116
rect 153516 198112 153580 198116
rect 153516 198056 153530 198112
rect 153530 198056 153580 198112
rect 153516 198052 153580 198056
rect 102916 197916 102980 197980
rect 153148 197916 153212 197980
rect 154436 197916 154500 197980
rect 165292 197916 165356 197980
rect 172284 197916 172348 197980
rect 157748 197780 157812 197844
rect 187004 197780 187068 197844
rect 176332 197644 176396 197708
rect 164924 197508 164988 197572
rect 188108 197508 188172 197572
rect 164740 197372 164804 197436
rect 173756 197372 173820 197436
rect 175964 197372 176028 197436
rect 136588 197236 136652 197300
rect 139716 197296 139780 197300
rect 139716 197240 139766 197296
rect 139766 197240 139780 197296
rect 139716 197236 139780 197240
rect 162348 197236 162412 197300
rect 136956 197100 137020 197164
rect 136772 196888 136836 196892
rect 136772 196832 136822 196888
rect 136822 196832 136836 196888
rect 136772 196828 136836 196832
rect 137508 196888 137572 196892
rect 137508 196832 137522 196888
rect 137522 196832 137572 196888
rect 137508 196828 137572 196832
rect 138060 196828 138124 196892
rect 142476 196828 142540 196892
rect 146708 196828 146772 196892
rect 147076 196828 147140 196892
rect 157196 196888 157260 196892
rect 157196 196832 157210 196888
rect 157210 196832 157260 196888
rect 157196 196828 157260 196832
rect 162532 196828 162596 196892
rect 163452 196828 163516 196892
rect 197308 196828 197372 196892
rect 157196 196692 157260 196756
rect 113036 196556 113100 196620
rect 148180 196556 148244 196620
rect 157564 196556 157628 196620
rect 142292 196420 142356 196484
rect 161060 196420 161124 196484
rect 163084 196420 163148 196484
rect 164924 196480 164988 196484
rect 164924 196424 164974 196480
rect 164974 196424 164988 196480
rect 164924 196420 164988 196424
rect 167684 196420 167748 196484
rect 169156 196480 169220 196484
rect 169156 196424 169170 196480
rect 169170 196424 169220 196480
rect 169156 196420 169220 196424
rect 170812 196420 170876 196484
rect 171364 196480 171428 196484
rect 171364 196424 171378 196480
rect 171378 196424 171428 196480
rect 171364 196420 171428 196424
rect 193260 196420 193324 196484
rect 134012 196284 134076 196348
rect 163820 196284 163884 196348
rect 166028 196344 166092 196348
rect 166028 196288 166078 196344
rect 166078 196288 166092 196344
rect 166028 196284 166092 196288
rect 168788 196284 168852 196348
rect 170076 196284 170140 196348
rect 172468 196344 172532 196348
rect 172468 196288 172518 196344
rect 172518 196288 172532 196344
rect 172468 196284 172532 196288
rect 173388 196284 173452 196348
rect 135300 196208 135364 196212
rect 135300 196152 135314 196208
rect 135314 196152 135364 196208
rect 135300 196148 135364 196152
rect 167500 196148 167564 196212
rect 169524 196148 169588 196212
rect 170628 196148 170692 196212
rect 171916 196148 171980 196212
rect 135300 196012 135364 196076
rect 158116 196012 158180 196076
rect 161428 196012 161492 196076
rect 165844 196012 165908 196076
rect 169892 196012 169956 196076
rect 135668 195876 135732 195940
rect 142844 195876 142908 195940
rect 184060 195876 184124 195940
rect 130332 195740 130396 195804
rect 139532 195740 139596 195804
rect 161796 195740 161860 195804
rect 166580 195740 166644 195804
rect 104020 195604 104084 195668
rect 146892 195604 146956 195668
rect 153884 195604 153948 195668
rect 160140 195332 160204 195396
rect 194548 195332 194612 195396
rect 119844 195196 119908 195260
rect 199332 195060 199396 195124
rect 175412 194788 175476 194852
rect 201724 194516 201788 194580
rect 102732 194380 102796 194444
rect 147260 194380 147324 194444
rect 173020 194380 173084 194444
rect 142292 194304 142356 194308
rect 142292 194248 142306 194304
rect 142306 194248 142356 194304
rect 142292 194244 142356 194248
rect 172652 194108 172716 194172
rect 173572 194032 173636 194036
rect 173572 193976 173622 194032
rect 173622 193976 173636 194032
rect 173572 193972 173636 193976
rect 175596 193972 175660 194036
rect 210004 193972 210068 194036
rect 100340 193836 100404 193900
rect 209820 193836 209884 193900
rect 201908 193156 201972 193220
rect 198780 193020 198844 193084
rect 201540 192884 201604 192948
rect 186084 192612 186148 192676
rect 103100 192476 103164 192540
rect 134012 191660 134076 191724
rect 135484 191388 135548 191452
rect 134196 191252 134260 191316
rect 139716 191116 139780 191180
rect 185348 191116 185412 191180
rect 135668 190980 135732 191044
rect 164924 190980 164988 191044
rect 138428 190028 138492 190092
rect 172284 190028 172348 190092
rect 100524 189892 100588 189956
rect 104204 189756 104268 189820
rect 136956 189756 137020 189820
rect 138244 189620 138308 189684
rect 158116 189620 158180 189684
rect 108436 187172 108500 187236
rect 108252 187036 108316 187100
rect 157012 187036 157076 187100
rect 139532 186900 139596 186964
rect 152964 186900 153028 186964
rect 169156 155620 169220 155684
rect 169340 155484 169404 155548
rect 176332 155348 176396 155412
rect 161244 155212 161308 155276
rect 148916 152356 148980 152420
rect 124076 151676 124140 151740
rect 108804 151404 108868 151468
rect 190500 151404 190564 151468
rect 136772 151268 136836 151332
rect 187740 151268 187804 151332
rect 138060 151132 138124 151196
rect 154436 151132 154500 151196
rect 136588 150996 136652 151060
rect 162348 150996 162412 151060
rect 191972 150452 192036 150516
rect 202092 150316 202156 150380
rect 207612 150316 207676 150380
rect 176516 150180 176580 150244
rect 203012 150044 203076 150108
rect 173756 149908 173820 149972
rect 202828 149908 202892 149972
rect 113404 149772 113468 149836
rect 205772 149772 205836 149836
rect 135300 149636 135364 149700
rect 205588 149636 205652 149700
rect 187740 149500 187804 149564
rect 203380 149092 203444 149156
rect 104388 148820 104452 148884
rect 120764 148684 120828 148748
rect 115428 148548 115492 148612
rect 117820 148412 117884 148476
rect 113588 148276 113652 148340
rect 122236 148140 122300 148204
rect 142292 148004 142356 148068
rect 122052 147732 122116 147796
rect 139348 147596 139412 147660
rect 192156 147596 192220 147660
rect 112300 147460 112364 147524
rect 194732 147460 194796 147524
rect 196572 147460 196636 147524
rect 110828 147324 110892 147388
rect 193812 147324 193876 147388
rect 115060 147188 115124 147252
rect 196204 147188 196268 147252
rect 112668 147052 112732 147116
rect 143580 147052 143644 147116
rect 197860 147052 197924 147116
rect 142476 146916 142540 146980
rect 157196 146916 157260 146980
rect 113956 146780 114020 146844
rect 197676 146780 197740 146844
rect 199516 146780 199580 146844
rect 122788 146704 122852 146708
rect 122788 146648 122802 146704
rect 122802 146648 122852 146704
rect 122788 146644 122852 146648
rect 109356 146236 109420 146300
rect 199332 146236 199396 146300
rect 109540 146100 109604 146164
rect 197676 146100 197740 146164
rect 116164 145964 116228 146028
rect 147076 145964 147140 146028
rect 196020 145964 196084 146028
rect 115796 145828 115860 145892
rect 199148 145828 199212 145892
rect 119660 145692 119724 145756
rect 112852 145556 112916 145620
rect 111196 145420 111260 145484
rect 193996 144740 194060 144804
rect 114140 144604 114204 144668
rect 189580 144604 189644 144668
rect 198964 144468 199028 144532
rect 111564 144332 111628 144396
rect 193444 144332 193508 144396
rect 116348 144196 116412 144260
rect 148180 144196 148244 144260
rect 189212 144196 189276 144260
rect 193628 144060 193692 144124
rect 116716 143924 116780 143988
rect 187188 143380 187252 143444
rect 111380 143244 111444 143308
rect 121316 143108 121380 143172
rect 121132 142972 121196 143036
rect 115612 142836 115676 142900
rect 130332 142836 130396 142900
rect 118372 142700 118436 142764
rect 121316 142564 121380 142628
rect 111012 142428 111076 142492
rect 116900 141884 116964 141948
rect 112852 141612 112916 141676
rect 121132 141476 121196 141540
rect 185900 141476 185964 141540
rect 118188 141340 118252 141404
rect 118740 140720 118804 140724
rect 118740 140664 118790 140720
rect 118790 140664 118804 140720
rect 118740 140660 118804 140664
rect 120948 140660 121012 140724
rect 119476 140388 119540 140452
rect 129044 140448 129108 140452
rect 129044 140392 129094 140448
rect 129094 140392 129108 140448
rect 129044 140388 129108 140392
rect 191604 140388 191668 140452
rect 124812 140312 124876 140316
rect 124812 140256 124862 140312
rect 124862 140256 124876 140312
rect 124812 140252 124876 140256
rect 126836 140252 126900 140316
rect 190868 140252 190932 140316
rect 146524 140116 146588 140180
rect 186268 140116 186332 140180
rect 146892 139980 146956 140044
rect 189396 139980 189460 140044
rect 116532 139708 116596 139772
rect 197492 139708 197556 139772
rect 124444 139632 124508 139636
rect 124444 139576 124494 139632
rect 124494 139576 124508 139632
rect 124444 139572 124508 139576
rect 125364 139572 125428 139636
rect 127388 139572 127452 139636
rect 188292 139572 188356 139636
rect 111196 139300 111260 139364
rect 115060 139300 115124 139364
rect 122972 139300 123036 139364
rect 124076 139300 124140 139364
rect 124260 139300 124324 139364
rect 118004 139164 118068 139228
rect 124444 139028 124508 139092
rect 124260 138892 124324 138956
rect 109540 138756 109604 138820
rect 125364 138756 125428 138820
rect 129044 138620 129108 138684
rect 191788 139436 191852 139500
rect 121316 138484 121380 138548
rect 124812 138348 124876 138412
rect 127388 138212 127452 138276
rect 185348 138212 185412 138276
rect 186636 138212 186700 138276
rect 122788 138076 122852 138140
rect 185900 138076 185964 138140
rect 186452 138076 186516 138140
rect 187188 138076 187252 138140
rect 188292 138076 188356 138140
rect 113772 137940 113836 138004
rect 123892 137940 123956 138004
rect 184060 137940 184124 138004
rect 126836 137804 126900 137868
rect 185348 137804 185412 137868
rect 199332 137260 199396 137324
rect 203564 136580 203628 136644
rect 186452 136036 186516 136100
rect 186636 135900 186700 135964
rect 122788 132500 122852 132564
rect 122788 132364 122852 132428
rect 122788 122844 122852 122908
rect 122788 122708 122852 122772
rect 122788 113188 122852 113252
rect 122788 113052 122852 113116
rect 122788 103532 122852 103596
rect 122788 103396 122852 103460
rect 118740 96596 118804 96660
rect 122788 93876 122852 93940
rect 186084 93740 186148 93804
rect 122788 92380 122852 92444
rect 186084 90340 186148 90404
rect 186084 84628 186148 84692
rect 186820 84628 186884 84692
rect 186452 82044 186516 82108
rect 125548 81908 125612 81972
rect 185716 81772 185780 81836
rect 186268 81772 186332 81836
rect 184060 81636 184124 81700
rect 181300 81500 181364 81564
rect 186268 81500 186332 81564
rect 185348 81364 185412 81428
rect 186820 81364 186884 81428
rect 201172 81424 201236 81428
rect 201172 81368 201222 81424
rect 201222 81368 201236 81424
rect 201172 81364 201236 81368
rect 176332 81228 176396 81292
rect 197676 81228 197740 81292
rect 129228 81092 129292 81156
rect 170444 81092 170508 81156
rect 192156 81092 192220 81156
rect 146892 80956 146956 81020
rect 174676 80956 174740 81020
rect 199148 80956 199212 81020
rect 149836 80820 149900 80884
rect 121132 80684 121196 80748
rect 129228 80548 129292 80612
rect 170628 80684 170692 80748
rect 196204 80820 196268 80884
rect 134012 79868 134076 79932
rect 133828 79596 133892 79660
rect 135484 79868 135548 79932
rect 133460 79460 133524 79524
rect 137692 79868 137756 79932
rect 138060 79868 138124 79932
rect 138980 79906 138984 79932
rect 138984 79906 139040 79932
rect 139040 79906 139044 79932
rect 138980 79868 139044 79906
rect 138612 79792 138676 79796
rect 138612 79736 138626 79792
rect 138626 79736 138676 79792
rect 138612 79732 138676 79736
rect 139716 79906 139720 79932
rect 139720 79906 139776 79932
rect 139776 79906 139780 79932
rect 139716 79868 139780 79906
rect 140084 79868 140148 79932
rect 141004 79868 141068 79932
rect 139900 79732 139964 79796
rect 143396 80004 143460 80068
rect 142660 79928 142724 79932
rect 142660 79872 142664 79928
rect 142664 79872 142720 79928
rect 142720 79872 142724 79928
rect 142660 79868 142724 79872
rect 143580 79928 143644 79932
rect 143580 79872 143584 79928
rect 143584 79872 143640 79928
rect 143640 79872 143644 79928
rect 143580 79868 143644 79872
rect 151308 80140 151372 80204
rect 173204 80276 173268 80340
rect 189028 80276 189092 80340
rect 138244 79596 138308 79660
rect 144316 79656 144380 79660
rect 144316 79600 144330 79656
rect 144330 79600 144380 79656
rect 144316 79596 144380 79600
rect 145604 79868 145668 79932
rect 145420 79460 145484 79524
rect 147076 79868 147140 79932
rect 147812 79906 147816 79932
rect 147816 79906 147872 79932
rect 147872 79906 147876 79932
rect 147812 79868 147876 79906
rect 148180 79906 148184 79932
rect 148184 79906 148240 79932
rect 148240 79906 148244 79932
rect 148180 79868 148244 79906
rect 146524 79732 146588 79796
rect 146892 79596 146956 79660
rect 149836 79868 149900 79932
rect 153884 79868 153948 79932
rect 152780 79732 152844 79796
rect 154988 79906 154992 79932
rect 154992 79906 155048 79932
rect 155048 79906 155052 79932
rect 154988 79868 155052 79906
rect 155540 79732 155604 79796
rect 155908 79906 155912 79932
rect 155912 79906 155968 79932
rect 155968 79906 155972 79932
rect 155908 79868 155972 79906
rect 157932 79868 157996 79932
rect 158484 79732 158548 79796
rect 147812 79384 147876 79388
rect 147812 79328 147862 79384
rect 147862 79328 147876 79384
rect 147812 79324 147876 79328
rect 148180 79384 148244 79388
rect 148180 79328 148194 79384
rect 148194 79328 148244 79384
rect 148180 79324 148244 79328
rect 154436 79324 154500 79388
rect 119660 79188 119724 79252
rect 156644 79188 156708 79252
rect 158116 79188 158180 79252
rect 159956 79928 160020 79932
rect 159956 79872 159960 79928
rect 159960 79872 160016 79928
rect 160016 79872 160020 79928
rect 159956 79868 160020 79872
rect 187740 80140 187804 80204
rect 188292 80140 188356 80204
rect 170444 80004 170508 80068
rect 161060 79868 161124 79932
rect 161244 79732 161308 79796
rect 162164 79868 162228 79932
rect 163268 79868 163332 79932
rect 163452 79868 163516 79932
rect 164556 79928 164620 79932
rect 164556 79872 164560 79928
rect 164560 79872 164616 79928
rect 164616 79872 164620 79928
rect 164556 79868 164620 79872
rect 165292 79868 165356 79932
rect 162532 79792 162596 79796
rect 162532 79736 162536 79792
rect 162536 79736 162592 79792
rect 162592 79736 162596 79792
rect 162532 79732 162596 79736
rect 163636 79596 163700 79660
rect 165108 79732 165172 79796
rect 166028 79906 166032 79932
rect 166032 79906 166088 79932
rect 166088 79906 166092 79932
rect 166028 79868 166092 79906
rect 166580 79868 166644 79932
rect 167868 79928 167932 79932
rect 167868 79872 167872 79928
rect 167872 79872 167928 79928
rect 167928 79872 167932 79928
rect 167868 79868 167932 79872
rect 166764 79732 166828 79796
rect 167684 79792 167748 79796
rect 167684 79736 167688 79792
rect 167688 79736 167744 79792
rect 167744 79736 167748 79792
rect 167684 79732 167748 79736
rect 168052 79792 168116 79796
rect 168052 79736 168056 79792
rect 168056 79736 168112 79792
rect 168112 79736 168116 79792
rect 168052 79732 168116 79736
rect 166396 79596 166460 79660
rect 170076 79868 170140 79932
rect 170996 79868 171060 79932
rect 171916 79868 171980 79932
rect 172100 79868 172164 79932
rect 173572 79868 173636 79932
rect 174676 79868 174740 79932
rect 176516 80004 176580 80068
rect 205772 80004 205836 80068
rect 170076 79732 170140 79796
rect 175964 79868 176028 79932
rect 171180 79732 171244 79796
rect 174492 79732 174556 79796
rect 169524 79460 169588 79524
rect 170628 79520 170692 79524
rect 170628 79464 170678 79520
rect 170678 79464 170692 79520
rect 170628 79460 170692 79464
rect 173756 79596 173820 79660
rect 175044 79596 175108 79660
rect 176332 79596 176396 79660
rect 186268 79520 186332 79524
rect 186268 79464 186282 79520
rect 186282 79464 186332 79520
rect 186268 79460 186332 79464
rect 189396 79324 189460 79388
rect 190868 79188 190932 79252
rect 120948 79052 121012 79116
rect 155908 79052 155972 79116
rect 143580 78976 143644 78980
rect 143580 78920 143594 78976
rect 143594 78920 143644 78976
rect 143580 78916 143644 78920
rect 158852 78780 158916 78844
rect 194732 79052 194796 79116
rect 173204 78916 173268 78980
rect 203012 78916 203076 78980
rect 158300 78644 158364 78708
rect 159956 78644 160020 78708
rect 134196 78568 134260 78572
rect 134196 78512 134210 78568
rect 134210 78512 134260 78568
rect 134196 78508 134260 78512
rect 138428 78508 138492 78572
rect 139348 78508 139412 78572
rect 148364 78508 148428 78572
rect 149468 78508 149532 78572
rect 170812 78508 170876 78572
rect 170996 78568 171060 78572
rect 170996 78512 171046 78568
rect 171046 78512 171060 78568
rect 170996 78508 171060 78512
rect 176332 78508 176396 78572
rect 134012 78372 134076 78436
rect 107516 77828 107580 77892
rect 122972 78236 123036 78300
rect 134012 78236 134076 78300
rect 137508 78236 137572 78300
rect 140820 78236 140884 78300
rect 157012 78236 157076 78300
rect 190500 78236 190564 78300
rect 149836 78100 149900 78164
rect 154988 78100 155052 78164
rect 138980 78024 139044 78028
rect 138980 77968 138994 78024
rect 138994 77968 139044 78024
rect 138980 77964 139044 77968
rect 143764 77964 143828 78028
rect 155724 77964 155788 78028
rect 141004 77828 141068 77892
rect 142660 77828 142724 77892
rect 143948 77828 144012 77892
rect 133276 77752 133340 77756
rect 133276 77696 133326 77752
rect 133326 77696 133340 77752
rect 133276 77692 133340 77696
rect 176148 77692 176212 77756
rect 188108 77692 188172 77756
rect 135300 77556 135364 77620
rect 147996 77556 148060 77620
rect 146892 77420 146956 77484
rect 148548 77480 148612 77484
rect 148548 77424 148598 77480
rect 148598 77424 148612 77480
rect 148548 77420 148612 77424
rect 150020 77420 150084 77484
rect 151676 77420 151740 77484
rect 152596 77420 152660 77484
rect 134380 77284 134444 77348
rect 135668 77284 135732 77348
rect 147444 77284 147508 77348
rect 147812 77284 147876 77348
rect 149652 77344 149716 77348
rect 149652 77288 149666 77344
rect 149666 77288 149716 77344
rect 149652 77284 149716 77288
rect 149836 77284 149900 77348
rect 164924 77284 164988 77348
rect 119660 77148 119724 77212
rect 174676 77148 174740 77212
rect 210004 77148 210068 77212
rect 160692 76876 160756 76940
rect 164556 76876 164620 76940
rect 167868 76876 167932 76940
rect 199516 76876 199580 76940
rect 111196 76604 111260 76668
rect 133092 76604 133156 76668
rect 152412 76740 152476 76804
rect 160876 76740 160940 76804
rect 162348 76800 162412 76804
rect 162348 76744 162362 76800
rect 162362 76744 162412 76800
rect 162348 76740 162412 76744
rect 165476 76740 165540 76804
rect 166028 76740 166092 76804
rect 167868 76800 167932 76804
rect 167868 76744 167882 76800
rect 167882 76744 167932 76800
rect 167868 76740 167932 76744
rect 169340 76800 169404 76804
rect 169340 76744 169354 76800
rect 169354 76744 169404 76800
rect 169340 76740 169404 76744
rect 170444 76740 170508 76804
rect 193812 76740 193876 76804
rect 191972 76604 192036 76668
rect 154252 76332 154316 76396
rect 191604 76332 191668 76396
rect 174860 76196 174924 76260
rect 187924 76196 187988 76260
rect 153884 76060 153948 76124
rect 170628 75924 170692 75988
rect 119660 75788 119724 75852
rect 113036 75652 113100 75716
rect 147444 75652 147508 75716
rect 156828 75712 156892 75716
rect 156828 75656 156842 75712
rect 156842 75656 156892 75712
rect 156828 75652 156892 75656
rect 122420 75516 122484 75580
rect 145604 75380 145668 75444
rect 202092 75380 202156 75444
rect 112668 75244 112732 75308
rect 157196 75244 157260 75308
rect 159036 75244 159100 75308
rect 185900 75244 185964 75308
rect 119660 75108 119724 75172
rect 187004 75108 187068 75172
rect 125548 74972 125612 75036
rect 170076 74972 170140 75036
rect 122788 74564 122852 74628
rect 117084 74428 117148 74492
rect 185900 74428 185964 74492
rect 113588 74292 113652 74356
rect 148548 74292 148612 74356
rect 134380 74156 134444 74220
rect 106780 74020 106844 74084
rect 122604 74020 122668 74084
rect 149468 74156 149532 74220
rect 118556 73884 118620 73948
rect 197860 73884 197924 73948
rect 196020 73612 196084 73676
rect 151676 73340 151740 73404
rect 145420 73068 145484 73132
rect 146524 72932 146588 72996
rect 147076 72796 147140 72860
rect 148364 72660 148428 72724
rect 205772 72660 205836 72724
rect 188292 72388 188356 72452
rect 116164 71708 116228 71772
rect 115428 71572 115492 71636
rect 122052 71436 122116 71500
rect 146892 71300 146956 71364
rect 184060 71300 184124 71364
rect 200988 71300 201052 71364
rect 122604 71164 122668 71228
rect 106964 71028 107028 71092
rect 117820 70212 117884 70276
rect 113956 70076 114020 70140
rect 120764 69940 120828 70004
rect 122236 69804 122300 69868
rect 147812 69668 147876 69732
rect 148364 69668 148428 69732
rect 103100 68912 103164 68916
rect 103100 68856 103114 68912
rect 103114 68856 103164 68912
rect 103100 68852 103164 68856
rect 118004 68852 118068 68916
rect 118188 68716 118252 68780
rect 187924 68852 187988 68916
rect 189580 68852 189644 68916
rect 200804 68912 200868 68916
rect 200804 68856 200818 68912
rect 200818 68856 200868 68912
rect 200804 68852 200868 68856
rect 181300 68716 181364 68780
rect 116348 68580 116412 68644
rect 144132 68444 144196 68508
rect 149652 68444 149716 68508
rect 147444 68308 147508 68372
rect 102916 68172 102980 68236
rect 146524 68172 146588 68236
rect 145604 67628 145668 67692
rect 144316 67492 144380 67556
rect 149836 67492 149900 67556
rect 113404 67356 113468 67420
rect 114140 67356 114204 67420
rect 115612 67356 115676 67420
rect 147996 67356 148060 67420
rect 170628 67356 170692 67420
rect 140820 67220 140884 67284
rect 108436 66948 108500 67012
rect 104020 66812 104084 66876
rect 108252 66132 108316 66196
rect 124076 66132 124140 66196
rect 170812 66132 170876 66196
rect 109540 65996 109604 66060
rect 203564 66056 203628 66060
rect 203564 66000 203614 66056
rect 203614 66000 203628 66056
rect 203564 65996 203628 66000
rect 110828 65860 110892 65924
rect 139900 65860 139964 65924
rect 108804 65724 108868 65788
rect 112852 65588 112916 65652
rect 135668 64772 135732 64836
rect 143580 64772 143644 64836
rect 144316 64772 144380 64836
rect 104204 64696 104268 64700
rect 104204 64640 104254 64696
rect 104254 64640 104268 64696
rect 104204 64636 104268 64640
rect 143764 64636 143828 64700
rect 144500 64636 144564 64700
rect 174492 64636 174556 64700
rect 200620 64636 200684 64700
rect 201356 64636 201420 64700
rect 143580 64500 143644 64564
rect 186084 64500 186148 64564
rect 187188 64560 187252 64564
rect 187188 64504 187202 64560
rect 187202 64504 187252 64560
rect 187188 64500 187252 64504
rect 156644 64364 156708 64428
rect 201356 64092 201420 64156
rect 138612 63412 138676 63476
rect 160692 63412 160756 63476
rect 100340 63276 100404 63340
rect 133460 63276 133524 63340
rect 174676 63276 174740 63340
rect 138428 63140 138492 63204
rect 100340 62732 100404 62796
rect 148548 62732 148612 62796
rect 102732 62112 102796 62116
rect 102732 62056 102746 62112
rect 102746 62056 102796 62112
rect 102732 62052 102796 62056
rect 139716 62052 139780 62116
rect 173572 62052 173636 62116
rect 199332 61916 199396 61980
rect 112300 60616 112364 60620
rect 112300 60560 112314 60616
rect 112314 60560 112364 60616
rect 112300 60556 112364 60560
rect 163268 60556 163332 60620
rect 150020 60420 150084 60484
rect 164924 60284 164988 60348
rect 191788 59876 191852 59940
rect 104388 59196 104452 59260
rect 172100 59196 172164 59260
rect 138244 57836 138308 57900
rect 152596 57836 152660 57900
rect 134196 57700 134260 57764
rect 175964 57700 176028 57764
rect 169340 57564 169404 57628
rect 165108 57428 165172 57492
rect 196572 57292 196636 57356
rect 147076 57156 147140 57220
rect 99420 56476 99484 56540
rect 100524 56476 100588 56540
rect 133276 56476 133340 56540
rect 157932 56476 157996 56540
rect 162348 56340 162412 56404
rect 154252 56204 154316 56268
rect 113772 55932 113836 55996
rect 99420 55796 99484 55860
rect 171916 55796 171980 55860
rect 139532 55116 139596 55180
rect 166396 55116 166460 55180
rect 139348 54980 139412 55044
rect 160876 54980 160940 55044
rect 203380 54768 203444 54772
rect 203380 54712 203394 54768
rect 203394 54712 203444 54768
rect 203380 54708 203444 54712
rect 137508 53756 137572 53820
rect 161060 53756 161124 53820
rect 194548 53756 194612 53820
rect 158116 53620 158180 53684
rect 146892 53076 146956 53140
rect 194548 53076 194612 53140
rect 114140 52532 114204 52596
rect 133092 52396 133156 52460
rect 193260 52456 193324 52460
rect 193260 52400 193274 52456
rect 193274 52400 193324 52456
rect 193260 52396 193324 52400
rect 201908 52456 201972 52460
rect 201908 52400 201958 52456
rect 201958 52400 201972 52456
rect 201908 52396 201972 52400
rect 156828 52260 156892 52324
rect 174860 52124 174924 52188
rect 152780 51988 152844 52052
rect 138060 50900 138124 50964
rect 207060 50900 207124 50964
rect 134012 50764 134076 50828
rect 158300 50764 158364 50828
rect 161244 50492 161308 50556
rect 193996 50492 194060 50556
rect 165292 50356 165356 50420
rect 176148 50220 176212 50284
rect 209820 50220 209884 50284
rect 133828 49540 133892 49604
rect 162532 49540 162596 49604
rect 176332 49404 176396 49468
rect 135484 48180 135548 48244
rect 170996 48180 171060 48244
rect 163452 48044 163516 48108
rect 169524 47908 169588 47972
rect 135300 46820 135364 46884
rect 152412 46820 152476 46884
rect 167684 46684 167748 46748
rect 167868 46548 167932 46612
rect 207612 46684 207676 46748
rect 201724 46140 201788 46204
rect 207612 45596 207676 45660
rect 175044 45460 175108 45524
rect 148364 45324 148428 45388
rect 162164 45188 162228 45252
rect 166580 45052 166644 45116
rect 198780 45052 198844 45116
rect 173756 44916 173820 44980
rect 203012 44916 203076 44980
rect 116532 44236 116596 44300
rect 137692 44100 137756 44164
rect 154436 44100 154500 44164
rect 166764 43964 166828 44028
rect 163636 43828 163700 43892
rect 197308 43828 197372 43892
rect 168052 43420 168116 43484
rect 201540 43420 201604 43484
rect 155540 38524 155604 38588
rect 176516 37164 176580 37228
rect 157012 37028 157076 37092
rect 157196 35804 157260 35868
rect 144500 35124 144564 35188
rect 151308 34444 151372 34508
rect 148180 30908 148244 30972
rect 165476 26148 165540 26212
rect 145420 22612 145484 22676
rect 158484 21932 158548 21996
rect 158852 21796 158916 21860
rect 159036 21660 159100 21724
rect 155724 17852 155788 17916
rect 111012 10236 111076 10300
rect 144316 8876 144380 8940
rect 144132 6156 144196 6220
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 682954 -8106 711002
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 -8106 682954
rect -8726 682634 -8106 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 -8106 682634
rect -8726 646954 -8106 682398
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 -8106 646954
rect -8726 646634 -8106 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 -8106 646634
rect -8726 610954 -8106 646398
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 -8106 610954
rect -8726 610634 -8106 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 -8106 610634
rect -8726 574954 -8106 610398
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 -8106 574954
rect -8726 574634 -8106 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 -8106 574634
rect -8726 538954 -8106 574398
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 -8106 538954
rect -8726 538634 -8106 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 -8106 538634
rect -8726 502954 -8106 538398
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 -8106 502954
rect -8726 502634 -8106 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 -8106 502634
rect -8726 466954 -8106 502398
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 -8106 466954
rect -8726 466634 -8106 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 -8106 466634
rect -8726 430954 -8106 466398
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 -8106 430954
rect -8726 430634 -8106 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 -8106 430634
rect -8726 394954 -8106 430398
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 -8106 394954
rect -8726 394634 -8106 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 -8106 394634
rect -8726 358954 -8106 394398
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 -8106 358954
rect -8726 358634 -8106 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 -8106 358634
rect -8726 322954 -8106 358398
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 -8106 322954
rect -8726 322634 -8106 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 -8106 322634
rect -8726 286954 -8106 322398
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 -8106 286954
rect -8726 286634 -8106 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 -8106 286634
rect -8726 250954 -8106 286398
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 -8106 250954
rect -8726 250634 -8106 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 -8106 250634
rect -8726 214954 -8106 250398
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 -8106 214954
rect -8726 214634 -8106 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 -8106 214634
rect -8726 178954 -8106 214398
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 -8106 178954
rect -8726 178634 -8106 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 -8106 178634
rect -8726 142954 -8106 178398
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 -8106 142954
rect -8726 142634 -8106 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 -8106 142634
rect -8726 106954 -8106 142398
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 -8106 106954
rect -8726 106634 -8106 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 -8106 106634
rect -8726 70954 -8106 106398
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 -8106 70954
rect -8726 70634 -8106 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 -8106 70634
rect -8726 34954 -8106 70398
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 -8106 34954
rect -8726 34634 -8106 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 -8106 34634
rect -8726 -7066 -8106 34398
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 678454 -7146 710042
rect -7766 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 -7146 678454
rect -7766 678134 -7146 678218
rect -7766 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 -7146 678134
rect -7766 642454 -7146 677898
rect -7766 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 -7146 642454
rect -7766 642134 -7146 642218
rect -7766 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 -7146 642134
rect -7766 606454 -7146 641898
rect -7766 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 -7146 606454
rect -7766 606134 -7146 606218
rect -7766 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 -7146 606134
rect -7766 570454 -7146 605898
rect -7766 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 -7146 570454
rect -7766 570134 -7146 570218
rect -7766 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 -7146 570134
rect -7766 534454 -7146 569898
rect -7766 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 -7146 534454
rect -7766 534134 -7146 534218
rect -7766 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 -7146 534134
rect -7766 498454 -7146 533898
rect -7766 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 -7146 498454
rect -7766 498134 -7146 498218
rect -7766 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 -7146 498134
rect -7766 462454 -7146 497898
rect -7766 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 -7146 462454
rect -7766 462134 -7146 462218
rect -7766 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 -7146 462134
rect -7766 426454 -7146 461898
rect -7766 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 -7146 426454
rect -7766 426134 -7146 426218
rect -7766 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 -7146 426134
rect -7766 390454 -7146 425898
rect -7766 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 -7146 390454
rect -7766 390134 -7146 390218
rect -7766 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 -7146 390134
rect -7766 354454 -7146 389898
rect -7766 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 -7146 354454
rect -7766 354134 -7146 354218
rect -7766 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 -7146 354134
rect -7766 318454 -7146 353898
rect -7766 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 -7146 318454
rect -7766 318134 -7146 318218
rect -7766 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 -7146 318134
rect -7766 282454 -7146 317898
rect -7766 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 -7146 282454
rect -7766 282134 -7146 282218
rect -7766 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 -7146 282134
rect -7766 246454 -7146 281898
rect -7766 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 -7146 246454
rect -7766 246134 -7146 246218
rect -7766 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 -7146 246134
rect -7766 210454 -7146 245898
rect -7766 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 -7146 210454
rect -7766 210134 -7146 210218
rect -7766 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 -7146 210134
rect -7766 174454 -7146 209898
rect -7766 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 -7146 174454
rect -7766 174134 -7146 174218
rect -7766 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 -7146 174134
rect -7766 138454 -7146 173898
rect -7766 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 -7146 138454
rect -7766 138134 -7146 138218
rect -7766 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 -7146 138134
rect -7766 102454 -7146 137898
rect -7766 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 -7146 102454
rect -7766 102134 -7146 102218
rect -7766 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 -7146 102134
rect -7766 66454 -7146 101898
rect -7766 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 -7146 66454
rect -7766 66134 -7146 66218
rect -7766 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 -7146 66134
rect -7766 30454 -7146 65898
rect -7766 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 -7146 30454
rect -7766 30134 -7146 30218
rect -7766 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 -7146 30134
rect -7766 -6106 -7146 29898
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 673954 -6186 709082
rect -6806 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 -6186 673954
rect -6806 673634 -6186 673718
rect -6806 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 -6186 673634
rect -6806 637954 -6186 673398
rect -6806 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 -6186 637954
rect -6806 637634 -6186 637718
rect -6806 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 -6186 637634
rect -6806 601954 -6186 637398
rect -6806 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 -6186 601954
rect -6806 601634 -6186 601718
rect -6806 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 -6186 601634
rect -6806 565954 -6186 601398
rect -6806 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 -6186 565954
rect -6806 565634 -6186 565718
rect -6806 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 -6186 565634
rect -6806 529954 -6186 565398
rect -6806 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 -6186 529954
rect -6806 529634 -6186 529718
rect -6806 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 -6186 529634
rect -6806 493954 -6186 529398
rect -6806 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 -6186 493954
rect -6806 493634 -6186 493718
rect -6806 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 -6186 493634
rect -6806 457954 -6186 493398
rect -6806 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 -6186 457954
rect -6806 457634 -6186 457718
rect -6806 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 -6186 457634
rect -6806 421954 -6186 457398
rect -6806 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 -6186 421954
rect -6806 421634 -6186 421718
rect -6806 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 -6186 421634
rect -6806 385954 -6186 421398
rect -6806 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 -6186 385954
rect -6806 385634 -6186 385718
rect -6806 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 -6186 385634
rect -6806 349954 -6186 385398
rect -6806 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 -6186 349954
rect -6806 349634 -6186 349718
rect -6806 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 -6186 349634
rect -6806 313954 -6186 349398
rect -6806 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 -6186 313954
rect -6806 313634 -6186 313718
rect -6806 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 -6186 313634
rect -6806 277954 -6186 313398
rect -6806 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 -6186 277954
rect -6806 277634 -6186 277718
rect -6806 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 -6186 277634
rect -6806 241954 -6186 277398
rect -6806 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 -6186 241954
rect -6806 241634 -6186 241718
rect -6806 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 -6186 241634
rect -6806 205954 -6186 241398
rect -6806 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 -6186 205954
rect -6806 205634 -6186 205718
rect -6806 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 -6186 205634
rect -6806 169954 -6186 205398
rect -6806 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 -6186 169954
rect -6806 169634 -6186 169718
rect -6806 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 -6186 169634
rect -6806 133954 -6186 169398
rect -6806 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 -6186 133954
rect -6806 133634 -6186 133718
rect -6806 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 -6186 133634
rect -6806 97954 -6186 133398
rect -6806 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 -6186 97954
rect -6806 97634 -6186 97718
rect -6806 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 -6186 97634
rect -6806 61954 -6186 97398
rect -6806 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 -6186 61954
rect -6806 61634 -6186 61718
rect -6806 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 -6186 61634
rect -6806 25954 -6186 61398
rect -6806 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 -6186 25954
rect -6806 25634 -6186 25718
rect -6806 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 -6186 25634
rect -6806 -5146 -6186 25398
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 669454 -5226 708122
rect -5846 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 -5226 669454
rect -5846 669134 -5226 669218
rect -5846 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 -5226 669134
rect -5846 633454 -5226 668898
rect -5846 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 -5226 633454
rect -5846 633134 -5226 633218
rect -5846 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 -5226 633134
rect -5846 597454 -5226 632898
rect -5846 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 -5226 597454
rect -5846 597134 -5226 597218
rect -5846 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 -5226 597134
rect -5846 561454 -5226 596898
rect -5846 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 -5226 561454
rect -5846 561134 -5226 561218
rect -5846 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 -5226 561134
rect -5846 525454 -5226 560898
rect -5846 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 -5226 525454
rect -5846 525134 -5226 525218
rect -5846 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 -5226 525134
rect -5846 489454 -5226 524898
rect -5846 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 -5226 489454
rect -5846 489134 -5226 489218
rect -5846 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 -5226 489134
rect -5846 453454 -5226 488898
rect -5846 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 -5226 453454
rect -5846 453134 -5226 453218
rect -5846 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 -5226 453134
rect -5846 417454 -5226 452898
rect -5846 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 -5226 417454
rect -5846 417134 -5226 417218
rect -5846 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 -5226 417134
rect -5846 381454 -5226 416898
rect -5846 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 -5226 381454
rect -5846 381134 -5226 381218
rect -5846 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 -5226 381134
rect -5846 345454 -5226 380898
rect -5846 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 -5226 345454
rect -5846 345134 -5226 345218
rect -5846 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 -5226 345134
rect -5846 309454 -5226 344898
rect -5846 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 -5226 309454
rect -5846 309134 -5226 309218
rect -5846 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 -5226 309134
rect -5846 273454 -5226 308898
rect -5846 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 -5226 273454
rect -5846 273134 -5226 273218
rect -5846 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 -5226 273134
rect -5846 237454 -5226 272898
rect -5846 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 -5226 237454
rect -5846 237134 -5226 237218
rect -5846 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 -5226 237134
rect -5846 201454 -5226 236898
rect -5846 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 -5226 201454
rect -5846 201134 -5226 201218
rect -5846 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 -5226 201134
rect -5846 165454 -5226 200898
rect -5846 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 -5226 165454
rect -5846 165134 -5226 165218
rect -5846 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 -5226 165134
rect -5846 129454 -5226 164898
rect -5846 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 -5226 129454
rect -5846 129134 -5226 129218
rect -5846 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 -5226 129134
rect -5846 93454 -5226 128898
rect -5846 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 -5226 93454
rect -5846 93134 -5226 93218
rect -5846 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 -5226 93134
rect -5846 57454 -5226 92898
rect -5846 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 -5226 57454
rect -5846 57134 -5226 57218
rect -5846 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 -5226 57134
rect -5846 21454 -5226 56898
rect -5846 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 -5226 21454
rect -5846 21134 -5226 21218
rect -5846 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 -5226 21134
rect -5846 -4186 -5226 20898
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 700954 -4266 707162
rect -4886 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 -4266 700954
rect -4886 700634 -4266 700718
rect -4886 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 -4266 700634
rect -4886 664954 -4266 700398
rect -4886 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 -4266 664954
rect -4886 664634 -4266 664718
rect -4886 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 -4266 664634
rect -4886 628954 -4266 664398
rect -4886 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 -4266 628954
rect -4886 628634 -4266 628718
rect -4886 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 -4266 628634
rect -4886 592954 -4266 628398
rect -4886 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 -4266 592954
rect -4886 592634 -4266 592718
rect -4886 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 -4266 592634
rect -4886 556954 -4266 592398
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 -4266 556954
rect -4886 556634 -4266 556718
rect -4886 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 -4266 556634
rect -4886 520954 -4266 556398
rect -4886 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 -4266 520954
rect -4886 520634 -4266 520718
rect -4886 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 -4266 520634
rect -4886 484954 -4266 520398
rect -4886 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 -4266 484954
rect -4886 484634 -4266 484718
rect -4886 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 -4266 484634
rect -4886 448954 -4266 484398
rect -4886 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 -4266 448954
rect -4886 448634 -4266 448718
rect -4886 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 -4266 448634
rect -4886 412954 -4266 448398
rect -4886 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 -4266 412954
rect -4886 412634 -4266 412718
rect -4886 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 -4266 412634
rect -4886 376954 -4266 412398
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 -4266 376954
rect -4886 376634 -4266 376718
rect -4886 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 -4266 376634
rect -4886 340954 -4266 376398
rect -4886 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 -4266 340954
rect -4886 340634 -4266 340718
rect -4886 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 -4266 340634
rect -4886 304954 -4266 340398
rect -4886 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 -4266 304954
rect -4886 304634 -4266 304718
rect -4886 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 -4266 304634
rect -4886 268954 -4266 304398
rect -4886 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 -4266 268954
rect -4886 268634 -4266 268718
rect -4886 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 -4266 268634
rect -4886 232954 -4266 268398
rect -4886 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 -4266 232954
rect -4886 232634 -4266 232718
rect -4886 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 -4266 232634
rect -4886 196954 -4266 232398
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 -4266 196954
rect -4886 196634 -4266 196718
rect -4886 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 -4266 196634
rect -4886 160954 -4266 196398
rect -4886 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 -4266 160954
rect -4886 160634 -4266 160718
rect -4886 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 -4266 160634
rect -4886 124954 -4266 160398
rect -4886 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 -4266 124954
rect -4886 124634 -4266 124718
rect -4886 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 -4266 124634
rect -4886 88954 -4266 124398
rect -4886 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 -4266 88954
rect -4886 88634 -4266 88718
rect -4886 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 -4266 88634
rect -4886 52954 -4266 88398
rect -4886 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 -4266 52954
rect -4886 52634 -4266 52718
rect -4886 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 -4266 52634
rect -4886 16954 -4266 52398
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 -4266 16954
rect -4886 16634 -4266 16718
rect -4886 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 -4266 16634
rect -4886 -3226 -4266 16398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 696454 -3306 706202
rect -3926 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 -3306 696454
rect -3926 696134 -3306 696218
rect -3926 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 -3306 696134
rect -3926 660454 -3306 695898
rect -3926 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 -3306 660454
rect -3926 660134 -3306 660218
rect -3926 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 -3306 660134
rect -3926 624454 -3306 659898
rect -3926 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 -3306 624454
rect -3926 624134 -3306 624218
rect -3926 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 -3306 624134
rect -3926 588454 -3306 623898
rect -3926 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 -3306 588454
rect -3926 588134 -3306 588218
rect -3926 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 -3306 588134
rect -3926 552454 -3306 587898
rect -3926 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 -3306 552454
rect -3926 552134 -3306 552218
rect -3926 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 -3306 552134
rect -3926 516454 -3306 551898
rect -3926 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 -3306 516454
rect -3926 516134 -3306 516218
rect -3926 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 -3306 516134
rect -3926 480454 -3306 515898
rect -3926 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 -3306 480454
rect -3926 480134 -3306 480218
rect -3926 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 -3306 480134
rect -3926 444454 -3306 479898
rect -3926 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 -3306 444454
rect -3926 444134 -3306 444218
rect -3926 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 -3306 444134
rect -3926 408454 -3306 443898
rect -3926 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 -3306 408454
rect -3926 408134 -3306 408218
rect -3926 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 -3306 408134
rect -3926 372454 -3306 407898
rect -3926 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 -3306 372454
rect -3926 372134 -3306 372218
rect -3926 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 -3306 372134
rect -3926 336454 -3306 371898
rect -3926 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 -3306 336454
rect -3926 336134 -3306 336218
rect -3926 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 -3306 336134
rect -3926 300454 -3306 335898
rect -3926 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 -3306 300454
rect -3926 300134 -3306 300218
rect -3926 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 -3306 300134
rect -3926 264454 -3306 299898
rect -3926 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 -3306 264454
rect -3926 264134 -3306 264218
rect -3926 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 -3306 264134
rect -3926 228454 -3306 263898
rect -3926 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 -3306 228454
rect -3926 228134 -3306 228218
rect -3926 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 -3306 228134
rect -3926 192454 -3306 227898
rect -3926 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 -3306 192454
rect -3926 192134 -3306 192218
rect -3926 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 -3306 192134
rect -3926 156454 -3306 191898
rect -3926 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 -3306 156454
rect -3926 156134 -3306 156218
rect -3926 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 -3306 156134
rect -3926 120454 -3306 155898
rect -3926 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 -3306 120454
rect -3926 120134 -3306 120218
rect -3926 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 -3306 120134
rect -3926 84454 -3306 119898
rect -3926 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 -3306 84454
rect -3926 84134 -3306 84218
rect -3926 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 -3306 84134
rect -3926 48454 -3306 83898
rect -3926 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 -3306 48454
rect -3926 48134 -3306 48218
rect -3926 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 -3306 48134
rect -3926 12454 -3306 47898
rect -3926 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 -3306 12454
rect -3926 12134 -3306 12218
rect -3926 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 -3306 12134
rect -3926 -2266 -3306 11898
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691954 -2346 705242
rect -2966 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 -2346 691954
rect -2966 691634 -2346 691718
rect -2966 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 -2346 691634
rect -2966 655954 -2346 691398
rect -2966 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 -2346 655954
rect -2966 655634 -2346 655718
rect -2966 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 -2346 655634
rect -2966 619954 -2346 655398
rect -2966 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 -2346 619954
rect -2966 619634 -2346 619718
rect -2966 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 -2346 619634
rect -2966 583954 -2346 619398
rect -2966 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 -2346 583954
rect -2966 583634 -2346 583718
rect -2966 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 -2346 583634
rect -2966 547954 -2346 583398
rect -2966 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 -2346 547954
rect -2966 547634 -2346 547718
rect -2966 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 -2346 547634
rect -2966 511954 -2346 547398
rect -2966 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 -2346 511954
rect -2966 511634 -2346 511718
rect -2966 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 -2346 511634
rect -2966 475954 -2346 511398
rect -2966 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 -2346 475954
rect -2966 475634 -2346 475718
rect -2966 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 -2346 475634
rect -2966 439954 -2346 475398
rect -2966 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 -2346 439954
rect -2966 439634 -2346 439718
rect -2966 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 -2346 439634
rect -2966 403954 -2346 439398
rect -2966 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 -2346 403954
rect -2966 403634 -2346 403718
rect -2966 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 -2346 403634
rect -2966 367954 -2346 403398
rect -2966 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 -2346 367954
rect -2966 367634 -2346 367718
rect -2966 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 -2346 367634
rect -2966 331954 -2346 367398
rect -2966 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 -2346 331954
rect -2966 331634 -2346 331718
rect -2966 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 -2346 331634
rect -2966 295954 -2346 331398
rect -2966 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 -2346 295954
rect -2966 295634 -2346 295718
rect -2966 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 -2346 295634
rect -2966 259954 -2346 295398
rect -2966 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 -2346 259954
rect -2966 259634 -2346 259718
rect -2966 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 -2346 259634
rect -2966 223954 -2346 259398
rect -2966 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 -2346 223954
rect -2966 223634 -2346 223718
rect -2966 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 -2346 223634
rect -2966 187954 -2346 223398
rect -2966 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 -2346 187954
rect -2966 187634 -2346 187718
rect -2966 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 -2346 187634
rect -2966 151954 -2346 187398
rect -2966 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 -2346 151954
rect -2966 151634 -2346 151718
rect -2966 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 -2346 151634
rect -2966 115954 -2346 151398
rect -2966 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 -2346 115954
rect -2966 115634 -2346 115718
rect -2966 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 -2346 115634
rect -2966 79954 -2346 115398
rect -2966 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 -2346 79954
rect -2966 79634 -2346 79718
rect -2966 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 -2346 79634
rect -2966 43954 -2346 79398
rect -2966 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 -2346 43954
rect -2966 43634 -2346 43718
rect -2966 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 -2346 43634
rect -2966 7954 -2346 43398
rect -2966 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 -2346 7954
rect -2966 7634 -2346 7718
rect -2966 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 -2346 7634
rect -2966 -1306 -2346 7398
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 6294 705798 6914 711590
rect 6294 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 6914 705798
rect 6294 705478 6914 705562
rect 6294 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 6914 705478
rect 6294 691954 6914 705242
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1306 6914 7398
rect 6294 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 6914 -1306
rect 6294 -1626 6914 -1542
rect 6294 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 6914 -1626
rect 6294 -7654 6914 -1862
rect 10794 706758 11414 711590
rect 10794 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 11414 706758
rect 10794 706438 11414 706522
rect 10794 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 11414 706438
rect 10794 696454 11414 706202
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2266 11414 11898
rect 10794 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 11414 -2266
rect 10794 -2586 11414 -2502
rect 10794 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 11414 -2586
rect 10794 -7654 11414 -2822
rect 15294 707718 15914 711590
rect 15294 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 15914 707718
rect 15294 707398 15914 707482
rect 15294 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 15914 707398
rect 15294 700954 15914 707162
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3226 15914 16398
rect 15294 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 15914 -3226
rect 15294 -3546 15914 -3462
rect 15294 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 15914 -3546
rect 15294 -7654 15914 -3782
rect 19794 708678 20414 711590
rect 19794 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 20414 708678
rect 19794 708358 20414 708442
rect 19794 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 20414 708358
rect 19794 669454 20414 708122
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4186 20414 20898
rect 19794 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 20414 -4186
rect 19794 -4506 20414 -4422
rect 19794 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 20414 -4506
rect 19794 -7654 20414 -4742
rect 24294 709638 24914 711590
rect 24294 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 24914 709638
rect 24294 709318 24914 709402
rect 24294 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 24914 709318
rect 24294 673954 24914 709082
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 133954 24914 169398
rect 24294 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 24914 133954
rect 24294 133634 24914 133718
rect 24294 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 24914 133634
rect 24294 97954 24914 133398
rect 24294 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 24914 97954
rect 24294 97634 24914 97718
rect 24294 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 24914 97634
rect 24294 61954 24914 97398
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5146 24914 25398
rect 24294 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 24914 -5146
rect 24294 -5466 24914 -5382
rect 24294 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 24914 -5466
rect 24294 -7654 24914 -5702
rect 28794 710598 29414 711590
rect 28794 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 29414 710598
rect 28794 710278 29414 710362
rect 28794 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 29414 710278
rect 28794 678454 29414 710042
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 138454 29414 173898
rect 28794 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 29414 138454
rect 28794 138134 29414 138218
rect 28794 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 29414 138134
rect 28794 102454 29414 137898
rect 28794 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 29414 102454
rect 28794 102134 29414 102218
rect 28794 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 29414 102134
rect 28794 66454 29414 101898
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6106 29414 29898
rect 28794 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 29414 -6106
rect 28794 -6426 29414 -6342
rect 28794 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 29414 -6426
rect 28794 -7654 29414 -6662
rect 33294 711558 33914 711590
rect 33294 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 33914 711558
rect 33294 711238 33914 711322
rect 33294 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 33914 711238
rect 33294 682954 33914 711002
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 646954 33914 682398
rect 33294 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 33914 646954
rect 33294 646634 33914 646718
rect 33294 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 33914 646634
rect 33294 610954 33914 646398
rect 33294 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 33914 610954
rect 33294 610634 33914 610718
rect 33294 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 33914 610634
rect 33294 574954 33914 610398
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 33294 502954 33914 538398
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 33294 466954 33914 502398
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 33294 394954 33914 430398
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 142954 33914 178398
rect 33294 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 33914 142954
rect 33294 142634 33914 142718
rect 33294 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 33914 142634
rect 33294 106954 33914 142398
rect 33294 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 33914 106954
rect 33294 106634 33914 106718
rect 33294 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 33914 106634
rect 33294 70954 33914 106398
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7066 33914 34398
rect 33294 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 33914 -7066
rect 33294 -7386 33914 -7302
rect 33294 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 33914 -7386
rect 33294 -7654 33914 -7622
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 42294 705798 42914 711590
rect 42294 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 42914 705798
rect 42294 705478 42914 705562
rect 42294 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 42914 705478
rect 42294 691954 42914 705242
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 655954 42914 691398
rect 42294 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 42914 655954
rect 42294 655634 42914 655718
rect 42294 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 42914 655634
rect 42294 619954 42914 655398
rect 42294 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 42914 619954
rect 42294 619634 42914 619718
rect 42294 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 42914 619634
rect 42294 583954 42914 619398
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 511954 42914 547398
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 42294 475954 42914 511398
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42294 439954 42914 475398
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42294 151954 42914 187398
rect 42294 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 42914 151954
rect 42294 151634 42914 151718
rect 42294 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 42914 151634
rect 42294 115954 42914 151398
rect 42294 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 42914 115954
rect 42294 115634 42914 115718
rect 42294 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 42914 115634
rect 42294 79954 42914 115398
rect 42294 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 42914 79954
rect 42294 79634 42914 79718
rect 42294 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 42914 79634
rect 42294 43954 42914 79398
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1306 42914 7398
rect 42294 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 42914 -1306
rect 42294 -1626 42914 -1542
rect 42294 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 42914 -1626
rect 42294 -7654 42914 -1862
rect 46794 706758 47414 711590
rect 46794 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 47414 706758
rect 46794 706438 47414 706522
rect 46794 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 47414 706438
rect 46794 696454 47414 706202
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 660454 47414 695898
rect 46794 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 47414 660454
rect 46794 660134 47414 660218
rect 46794 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 47414 660134
rect 46794 624454 47414 659898
rect 46794 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 47414 624454
rect 46794 624134 47414 624218
rect 46794 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 47414 624134
rect 46794 588454 47414 623898
rect 46794 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 47414 588454
rect 46794 588134 47414 588218
rect 46794 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 47414 588134
rect 46794 552454 47414 587898
rect 46794 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 47414 552454
rect 46794 552134 47414 552218
rect 46794 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 47414 552134
rect 46794 516454 47414 551898
rect 46794 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 47414 516454
rect 46794 516134 47414 516218
rect 46794 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 47414 516134
rect 46794 480454 47414 515898
rect 46794 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 47414 480454
rect 46794 480134 47414 480218
rect 46794 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 47414 480134
rect 46794 444454 47414 479898
rect 46794 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 47414 444454
rect 46794 444134 47414 444218
rect 46794 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 47414 444134
rect 46794 408454 47414 443898
rect 46794 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 47414 408454
rect 46794 408134 47414 408218
rect 46794 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 47414 408134
rect 46794 372454 47414 407898
rect 46794 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 47414 372454
rect 46794 372134 47414 372218
rect 46794 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 47414 372134
rect 46794 336454 47414 371898
rect 46794 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 47414 336454
rect 46794 336134 47414 336218
rect 46794 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 47414 336134
rect 46794 300454 47414 335898
rect 46794 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 47414 300454
rect 46794 300134 47414 300218
rect 46794 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 47414 300134
rect 46794 264454 47414 299898
rect 46794 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 47414 264454
rect 46794 264134 47414 264218
rect 46794 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 47414 264134
rect 46794 228454 47414 263898
rect 46794 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 47414 228454
rect 46794 228134 47414 228218
rect 46794 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 47414 228134
rect 46794 192454 47414 227898
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46794 120454 47414 155898
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 84454 47414 119898
rect 46794 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 47414 84454
rect 46794 84134 47414 84218
rect 46794 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 47414 84134
rect 46794 48454 47414 83898
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2266 47414 11898
rect 46794 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 47414 -2266
rect 46794 -2586 47414 -2502
rect 46794 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 47414 -2586
rect 46794 -7654 47414 -2822
rect 51294 707718 51914 711590
rect 51294 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 51914 707718
rect 51294 707398 51914 707482
rect 51294 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 51914 707398
rect 51294 700954 51914 707162
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 664954 51914 700398
rect 51294 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 51914 664954
rect 51294 664634 51914 664718
rect 51294 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 51914 664634
rect 51294 628954 51914 664398
rect 51294 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 51914 628954
rect 51294 628634 51914 628718
rect 51294 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 51914 628634
rect 51294 592954 51914 628398
rect 51294 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 51914 592954
rect 51294 592634 51914 592718
rect 51294 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 51914 592634
rect 51294 556954 51914 592398
rect 51294 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 51914 556954
rect 51294 556634 51914 556718
rect 51294 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 51914 556634
rect 51294 520954 51914 556398
rect 51294 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 51914 520954
rect 51294 520634 51914 520718
rect 51294 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 51914 520634
rect 51294 484954 51914 520398
rect 51294 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 51914 484954
rect 51294 484634 51914 484718
rect 51294 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 51914 484634
rect 51294 448954 51914 484398
rect 51294 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 51914 448954
rect 51294 448634 51914 448718
rect 51294 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 51914 448634
rect 51294 412954 51914 448398
rect 51294 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 51914 412954
rect 51294 412634 51914 412718
rect 51294 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 51914 412634
rect 51294 376954 51914 412398
rect 51294 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 51914 376954
rect 51294 376634 51914 376718
rect 51294 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 51914 376634
rect 51294 340954 51914 376398
rect 51294 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 51914 340954
rect 51294 340634 51914 340718
rect 51294 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 51914 340634
rect 51294 304954 51914 340398
rect 51294 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 51914 304954
rect 51294 304634 51914 304718
rect 51294 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 51914 304634
rect 51294 268954 51914 304398
rect 51294 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 51914 268954
rect 51294 268634 51914 268718
rect 51294 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 51914 268634
rect 51294 232954 51914 268398
rect 51294 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 51914 232954
rect 51294 232634 51914 232718
rect 51294 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 51914 232634
rect 51294 196954 51914 232398
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 51294 160954 51914 196398
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 124954 51914 160398
rect 51294 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 51914 124954
rect 51294 124634 51914 124718
rect 51294 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 51914 124634
rect 51294 88954 51914 124398
rect 51294 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 51914 88954
rect 51294 88634 51914 88718
rect 51294 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 51914 88634
rect 51294 52954 51914 88398
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3226 51914 16398
rect 51294 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 51914 -3226
rect 51294 -3546 51914 -3462
rect 51294 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 51914 -3546
rect 51294 -7654 51914 -3782
rect 55794 708678 56414 711590
rect 55794 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 56414 708678
rect 55794 708358 56414 708442
rect 55794 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 56414 708358
rect 55794 669454 56414 708122
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4186 56414 20898
rect 55794 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 56414 -4186
rect 55794 -4506 56414 -4422
rect 55794 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 56414 -4506
rect 55794 -7654 56414 -4742
rect 60294 709638 60914 711590
rect 60294 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 60914 709638
rect 60294 709318 60914 709402
rect 60294 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 60914 709318
rect 60294 673954 60914 709082
rect 60294 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 60914 673954
rect 60294 673634 60914 673718
rect 60294 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 60914 673634
rect 60294 637954 60914 673398
rect 60294 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 60914 637954
rect 60294 637634 60914 637718
rect 60294 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 60914 637634
rect 60294 601954 60914 637398
rect 60294 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 60914 601954
rect 60294 601634 60914 601718
rect 60294 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 60914 601634
rect 60294 565954 60914 601398
rect 60294 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 60914 565954
rect 60294 565634 60914 565718
rect 60294 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 60914 565634
rect 60294 529954 60914 565398
rect 60294 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 60914 529954
rect 60294 529634 60914 529718
rect 60294 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 60914 529634
rect 60294 493954 60914 529398
rect 60294 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 60914 493954
rect 60294 493634 60914 493718
rect 60294 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 60914 493634
rect 60294 457954 60914 493398
rect 60294 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 60914 457954
rect 60294 457634 60914 457718
rect 60294 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 60914 457634
rect 60294 421954 60914 457398
rect 60294 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 60914 421954
rect 60294 421634 60914 421718
rect 60294 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 60914 421634
rect 60294 385954 60914 421398
rect 60294 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 60914 385954
rect 60294 385634 60914 385718
rect 60294 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 60914 385634
rect 60294 349954 60914 385398
rect 60294 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 60914 349954
rect 60294 349634 60914 349718
rect 60294 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 60914 349634
rect 60294 313954 60914 349398
rect 60294 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 60914 313954
rect 60294 313634 60914 313718
rect 60294 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 60914 313634
rect 60294 277954 60914 313398
rect 60294 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 60914 277954
rect 60294 277634 60914 277718
rect 60294 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 60914 277634
rect 60294 241954 60914 277398
rect 60294 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 60914 241954
rect 60294 241634 60914 241718
rect 60294 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 60914 241634
rect 60294 205954 60914 241398
rect 60294 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 60914 205954
rect 60294 205634 60914 205718
rect 60294 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 60914 205634
rect 60294 169954 60914 205398
rect 60294 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 60914 169954
rect 60294 169634 60914 169718
rect 60294 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 60914 169634
rect 60294 133954 60914 169398
rect 60294 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 60914 133954
rect 60294 133634 60914 133718
rect 60294 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 60914 133634
rect 60294 97954 60914 133398
rect 60294 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 60914 97954
rect 60294 97634 60914 97718
rect 60294 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 60914 97634
rect 60294 61954 60914 97398
rect 60294 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 60914 61954
rect 60294 61634 60914 61718
rect 60294 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 60914 61634
rect 60294 25954 60914 61398
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 60294 -5146 60914 25398
rect 60294 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 60914 -5146
rect 60294 -5466 60914 -5382
rect 60294 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 60914 -5466
rect 60294 -7654 60914 -5702
rect 64794 710598 65414 711590
rect 64794 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 65414 710598
rect 64794 710278 65414 710362
rect 64794 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 65414 710278
rect 64794 678454 65414 710042
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 642454 65414 677898
rect 64794 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 65414 642454
rect 64794 642134 65414 642218
rect 64794 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 65414 642134
rect 64794 606454 65414 641898
rect 64794 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 65414 606454
rect 64794 606134 65414 606218
rect 64794 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 65414 606134
rect 64794 570454 65414 605898
rect 64794 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 65414 570454
rect 64794 570134 65414 570218
rect 64794 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 65414 570134
rect 64794 534454 65414 569898
rect 64794 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 65414 534454
rect 64794 534134 65414 534218
rect 64794 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 65414 534134
rect 64794 498454 65414 533898
rect 64794 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 65414 498454
rect 64794 498134 65414 498218
rect 64794 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 65414 498134
rect 64794 462454 65414 497898
rect 64794 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 65414 462454
rect 64794 462134 65414 462218
rect 64794 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 65414 462134
rect 64794 426454 65414 461898
rect 64794 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 65414 426454
rect 64794 426134 65414 426218
rect 64794 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 65414 426134
rect 64794 390454 65414 425898
rect 64794 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 65414 390454
rect 64794 390134 65414 390218
rect 64794 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 65414 390134
rect 64794 354454 65414 389898
rect 64794 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 65414 354454
rect 64794 354134 65414 354218
rect 64794 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 65414 354134
rect 64794 318454 65414 353898
rect 64794 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 65414 318454
rect 64794 318134 65414 318218
rect 64794 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 65414 318134
rect 64794 282454 65414 317898
rect 64794 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 65414 282454
rect 64794 282134 65414 282218
rect 64794 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 65414 282134
rect 64794 246454 65414 281898
rect 64794 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 65414 246454
rect 64794 246134 65414 246218
rect 64794 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 65414 246134
rect 64794 210454 65414 245898
rect 64794 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 65414 210454
rect 64794 210134 65414 210218
rect 64794 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 65414 210134
rect 64794 174454 65414 209898
rect 64794 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 65414 174454
rect 64794 174134 65414 174218
rect 64794 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 65414 174134
rect 64794 138454 65414 173898
rect 64794 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 65414 138454
rect 64794 138134 65414 138218
rect 64794 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 65414 138134
rect 64794 102454 65414 137898
rect 64794 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 65414 102454
rect 64794 102134 65414 102218
rect 64794 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 65414 102134
rect 64794 66454 65414 101898
rect 64794 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 65414 66454
rect 64794 66134 65414 66218
rect 64794 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 65414 66134
rect 64794 30454 65414 65898
rect 64794 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 65414 30454
rect 64794 30134 65414 30218
rect 64794 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 65414 30134
rect 64794 -6106 65414 29898
rect 64794 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 65414 -6106
rect 64794 -6426 65414 -6342
rect 64794 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 65414 -6426
rect 64794 -7654 65414 -6662
rect 69294 711558 69914 711590
rect 69294 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 69914 711558
rect 69294 711238 69914 711322
rect 69294 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 69914 711238
rect 69294 682954 69914 711002
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 646954 69914 682398
rect 69294 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 69914 646954
rect 69294 646634 69914 646718
rect 69294 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 69914 646634
rect 69294 610954 69914 646398
rect 69294 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 69914 610954
rect 69294 610634 69914 610718
rect 69294 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 69914 610634
rect 69294 574954 69914 610398
rect 69294 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 69914 574954
rect 69294 574634 69914 574718
rect 69294 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 69914 574634
rect 69294 538954 69914 574398
rect 69294 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 69914 538954
rect 69294 538634 69914 538718
rect 69294 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 69914 538634
rect 69294 502954 69914 538398
rect 69294 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 69914 502954
rect 69294 502634 69914 502718
rect 69294 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 69914 502634
rect 69294 466954 69914 502398
rect 69294 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 69914 466954
rect 69294 466634 69914 466718
rect 69294 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 69914 466634
rect 69294 430954 69914 466398
rect 69294 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 69914 430954
rect 69294 430634 69914 430718
rect 69294 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 69914 430634
rect 69294 394954 69914 430398
rect 69294 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 69914 394954
rect 69294 394634 69914 394718
rect 69294 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 69914 394634
rect 69294 358954 69914 394398
rect 69294 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 69914 358954
rect 69294 358634 69914 358718
rect 69294 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 69914 358634
rect 69294 322954 69914 358398
rect 69294 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 69914 322954
rect 69294 322634 69914 322718
rect 69294 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 69914 322634
rect 69294 286954 69914 322398
rect 69294 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 69914 286954
rect 69294 286634 69914 286718
rect 69294 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 69914 286634
rect 69294 250954 69914 286398
rect 69294 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 69914 250954
rect 69294 250634 69914 250718
rect 69294 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 69914 250634
rect 69294 214954 69914 250398
rect 69294 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 69914 214954
rect 69294 214634 69914 214718
rect 69294 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 69914 214634
rect 69294 178954 69914 214398
rect 69294 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 69914 178954
rect 69294 178634 69914 178718
rect 69294 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 69914 178634
rect 69294 142954 69914 178398
rect 69294 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 69914 142954
rect 69294 142634 69914 142718
rect 69294 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 69914 142634
rect 69294 106954 69914 142398
rect 69294 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 69914 106954
rect 69294 106634 69914 106718
rect 69294 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 69914 106634
rect 69294 70954 69914 106398
rect 69294 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 69914 70954
rect 69294 70634 69914 70718
rect 69294 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 69914 70634
rect 69294 34954 69914 70398
rect 69294 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 69914 34954
rect 69294 34634 69914 34718
rect 69294 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 69914 34634
rect 69294 -7066 69914 34398
rect 69294 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 69914 -7066
rect 69294 -7386 69914 -7302
rect 69294 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 69914 -7386
rect 69294 -7654 69914 -7622
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 78294 705798 78914 711590
rect 78294 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 78914 705798
rect 78294 705478 78914 705562
rect 78294 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 78914 705478
rect 78294 691954 78914 705242
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 655954 78914 691398
rect 78294 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 78914 655954
rect 78294 655634 78914 655718
rect 78294 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 78914 655634
rect 78294 619954 78914 655398
rect 78294 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 78914 619954
rect 78294 619634 78914 619718
rect 78294 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 78914 619634
rect 78294 583954 78914 619398
rect 78294 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 78914 583954
rect 78294 583634 78914 583718
rect 78294 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 78914 583634
rect 78294 547954 78914 583398
rect 78294 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 78914 547954
rect 78294 547634 78914 547718
rect 78294 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 78914 547634
rect 78294 511954 78914 547398
rect 78294 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 78914 511954
rect 78294 511634 78914 511718
rect 78294 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 78914 511634
rect 78294 475954 78914 511398
rect 78294 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 78914 475954
rect 78294 475634 78914 475718
rect 78294 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 78914 475634
rect 78294 439954 78914 475398
rect 78294 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 78914 439954
rect 78294 439634 78914 439718
rect 78294 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 78914 439634
rect 78294 403954 78914 439398
rect 78294 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 78914 403954
rect 78294 403634 78914 403718
rect 78294 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 78914 403634
rect 78294 367954 78914 403398
rect 78294 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 78914 367954
rect 78294 367634 78914 367718
rect 78294 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 78914 367634
rect 78294 331954 78914 367398
rect 78294 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 78914 331954
rect 78294 331634 78914 331718
rect 78294 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 78914 331634
rect 78294 295954 78914 331398
rect 78294 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 78914 295954
rect 78294 295634 78914 295718
rect 78294 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 78914 295634
rect 78294 259954 78914 295398
rect 78294 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 78914 259954
rect 78294 259634 78914 259718
rect 78294 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 78914 259634
rect 78294 223954 78914 259398
rect 78294 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 78914 223954
rect 78294 223634 78914 223718
rect 78294 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 78914 223634
rect 78294 187954 78914 223398
rect 78294 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 78914 187954
rect 78294 187634 78914 187718
rect 78294 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 78914 187634
rect 78294 151954 78914 187398
rect 78294 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 78914 151954
rect 78294 151634 78914 151718
rect 78294 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 78914 151634
rect 78294 115954 78914 151398
rect 78294 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 78914 115954
rect 78294 115634 78914 115718
rect 78294 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 78914 115634
rect 78294 79954 78914 115398
rect 78294 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 78914 79954
rect 78294 79634 78914 79718
rect 78294 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 78914 79634
rect 78294 43954 78914 79398
rect 78294 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 78914 43954
rect 78294 43634 78914 43718
rect 78294 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 78914 43634
rect 78294 7954 78914 43398
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1306 78914 7398
rect 78294 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 78914 -1306
rect 78294 -1626 78914 -1542
rect 78294 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 78914 -1626
rect 78294 -7654 78914 -1862
rect 82794 706758 83414 711590
rect 82794 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 83414 706758
rect 82794 706438 83414 706522
rect 82794 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 83414 706438
rect 82794 696454 83414 706202
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 660454 83414 695898
rect 82794 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 83414 660454
rect 82794 660134 83414 660218
rect 82794 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 83414 660134
rect 82794 624454 83414 659898
rect 82794 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 83414 624454
rect 82794 624134 83414 624218
rect 82794 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 83414 624134
rect 82794 588454 83414 623898
rect 82794 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 83414 588454
rect 82794 588134 83414 588218
rect 82794 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 83414 588134
rect 82794 552454 83414 587898
rect 82794 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 83414 552454
rect 82794 552134 83414 552218
rect 82794 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 83414 552134
rect 82794 516454 83414 551898
rect 82794 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 83414 516454
rect 82794 516134 83414 516218
rect 82794 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 83414 516134
rect 82794 480454 83414 515898
rect 82794 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 83414 480454
rect 82794 480134 83414 480218
rect 82794 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 83414 480134
rect 82794 444454 83414 479898
rect 82794 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 83414 444454
rect 82794 444134 83414 444218
rect 82794 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 83414 444134
rect 82794 408454 83414 443898
rect 82794 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 83414 408454
rect 82794 408134 83414 408218
rect 82794 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 83414 408134
rect 82794 372454 83414 407898
rect 82794 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 83414 372454
rect 82794 372134 83414 372218
rect 82794 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 83414 372134
rect 82794 336454 83414 371898
rect 82794 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 83414 336454
rect 82794 336134 83414 336218
rect 82794 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 83414 336134
rect 82794 300454 83414 335898
rect 82794 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 83414 300454
rect 82794 300134 83414 300218
rect 82794 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 83414 300134
rect 82794 264454 83414 299898
rect 82794 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 83414 264454
rect 82794 264134 83414 264218
rect 82794 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 83414 264134
rect 82794 228454 83414 263898
rect 82794 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 83414 228454
rect 82794 228134 83414 228218
rect 82794 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 83414 228134
rect 82794 192454 83414 227898
rect 82794 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 83414 192454
rect 82794 192134 83414 192218
rect 82794 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 83414 192134
rect 82794 156454 83414 191898
rect 82794 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 83414 156454
rect 82794 156134 83414 156218
rect 82794 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 83414 156134
rect 82794 120454 83414 155898
rect 82794 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 83414 120454
rect 82794 120134 83414 120218
rect 82794 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 83414 120134
rect 82794 84454 83414 119898
rect 82794 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 83414 84454
rect 82794 84134 83414 84218
rect 82794 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 83414 84134
rect 82794 48454 83414 83898
rect 82794 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 83414 48454
rect 82794 48134 83414 48218
rect 82794 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 83414 48134
rect 82794 12454 83414 47898
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2266 83414 11898
rect 82794 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 83414 -2266
rect 82794 -2586 83414 -2502
rect 82794 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 83414 -2586
rect 82794 -7654 83414 -2822
rect 87294 707718 87914 711590
rect 87294 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 87914 707718
rect 87294 707398 87914 707482
rect 87294 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 87914 707398
rect 87294 700954 87914 707162
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 664954 87914 700398
rect 87294 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 87914 664954
rect 87294 664634 87914 664718
rect 87294 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 87914 664634
rect 87294 628954 87914 664398
rect 87294 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 87914 628954
rect 87294 628634 87914 628718
rect 87294 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 87914 628634
rect 87294 592954 87914 628398
rect 87294 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 87914 592954
rect 87294 592634 87914 592718
rect 87294 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 87914 592634
rect 87294 556954 87914 592398
rect 87294 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 87914 556954
rect 87294 556634 87914 556718
rect 87294 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 87914 556634
rect 87294 520954 87914 556398
rect 87294 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 87914 520954
rect 87294 520634 87914 520718
rect 87294 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 87914 520634
rect 87294 484954 87914 520398
rect 87294 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 87914 484954
rect 87294 484634 87914 484718
rect 87294 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 87914 484634
rect 87294 448954 87914 484398
rect 87294 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 87914 448954
rect 87294 448634 87914 448718
rect 87294 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 87914 448634
rect 87294 412954 87914 448398
rect 87294 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 87914 412954
rect 87294 412634 87914 412718
rect 87294 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 87914 412634
rect 87294 376954 87914 412398
rect 87294 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 87914 376954
rect 87294 376634 87914 376718
rect 87294 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 87914 376634
rect 87294 340954 87914 376398
rect 87294 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 87914 340954
rect 87294 340634 87914 340718
rect 87294 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 87914 340634
rect 87294 304954 87914 340398
rect 87294 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 87914 304954
rect 87294 304634 87914 304718
rect 87294 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 87914 304634
rect 87294 268954 87914 304398
rect 87294 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 87914 268954
rect 87294 268634 87914 268718
rect 87294 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 87914 268634
rect 87294 232954 87914 268398
rect 87294 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 87914 232954
rect 87294 232634 87914 232718
rect 87294 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 87914 232634
rect 87294 196954 87914 232398
rect 87294 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 87914 196954
rect 87294 196634 87914 196718
rect 87294 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 87914 196634
rect 87294 160954 87914 196398
rect 87294 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 87914 160954
rect 87294 160634 87914 160718
rect 87294 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 87914 160634
rect 87294 124954 87914 160398
rect 87294 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 87914 124954
rect 87294 124634 87914 124718
rect 87294 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 87914 124634
rect 87294 88954 87914 124398
rect 87294 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 87914 88954
rect 87294 88634 87914 88718
rect 87294 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 87914 88634
rect 87294 52954 87914 88398
rect 87294 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 87914 52954
rect 87294 52634 87914 52718
rect 87294 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 87914 52634
rect 87294 16954 87914 52398
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3226 87914 16398
rect 87294 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 87914 -3226
rect 87294 -3546 87914 -3462
rect 87294 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 87914 -3546
rect 87294 -7654 87914 -3782
rect 91794 708678 92414 711590
rect 91794 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 92414 708678
rect 91794 708358 92414 708442
rect 91794 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 92414 708358
rect 91794 669454 92414 708122
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4186 92414 20898
rect 91794 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 92414 -4186
rect 91794 -4506 92414 -4422
rect 91794 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 92414 -4506
rect 91794 -7654 92414 -4742
rect 96294 709638 96914 711590
rect 96294 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 96914 709638
rect 96294 709318 96914 709402
rect 96294 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 96914 709318
rect 96294 673954 96914 709082
rect 96294 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 96914 673954
rect 96294 673634 96914 673718
rect 96294 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 96914 673634
rect 96294 637954 96914 673398
rect 96294 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 96914 637954
rect 96294 637634 96914 637718
rect 96294 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 96914 637634
rect 96294 601954 96914 637398
rect 96294 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 96914 601954
rect 96294 601634 96914 601718
rect 96294 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 96914 601634
rect 96294 565954 96914 601398
rect 96294 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 96914 565954
rect 96294 565634 96914 565718
rect 96294 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 96914 565634
rect 96294 529954 96914 565398
rect 96294 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 96914 529954
rect 96294 529634 96914 529718
rect 96294 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 96914 529634
rect 96294 493954 96914 529398
rect 96294 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 96914 493954
rect 96294 493634 96914 493718
rect 96294 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 96914 493634
rect 96294 457954 96914 493398
rect 96294 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 96914 457954
rect 96294 457634 96914 457718
rect 96294 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 96914 457634
rect 96294 421954 96914 457398
rect 96294 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 96914 421954
rect 96294 421634 96914 421718
rect 96294 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 96914 421634
rect 96294 385954 96914 421398
rect 96294 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 96914 385954
rect 96294 385634 96914 385718
rect 96294 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 96914 385634
rect 96294 349954 96914 385398
rect 96294 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 96914 349954
rect 96294 349634 96914 349718
rect 96294 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 96914 349634
rect 96294 313954 96914 349398
rect 96294 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 96914 313954
rect 96294 313634 96914 313718
rect 96294 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 96914 313634
rect 96294 277954 96914 313398
rect 96294 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 96914 277954
rect 96294 277634 96914 277718
rect 96294 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 96914 277634
rect 96294 241954 96914 277398
rect 96294 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 96914 241954
rect 96294 241634 96914 241718
rect 96294 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 96914 241634
rect 96294 205954 96914 241398
rect 96294 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 96914 205954
rect 96294 205634 96914 205718
rect 96294 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 96914 205634
rect 96294 169954 96914 205398
rect 100794 710598 101414 711590
rect 100794 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 101414 710598
rect 100794 710278 101414 710362
rect 100794 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 101414 710278
rect 100794 678454 101414 710042
rect 100794 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 101414 678454
rect 100794 678134 101414 678218
rect 100794 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 101414 678134
rect 100794 642454 101414 677898
rect 100794 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 101414 642454
rect 100794 642134 101414 642218
rect 100794 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 101414 642134
rect 100794 606454 101414 641898
rect 100794 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 101414 606454
rect 100794 606134 101414 606218
rect 100794 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 101414 606134
rect 100794 570454 101414 605898
rect 100794 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 101414 570454
rect 100794 570134 101414 570218
rect 100794 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 101414 570134
rect 100794 534454 101414 569898
rect 100794 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 101414 534454
rect 100794 534134 101414 534218
rect 100794 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 101414 534134
rect 100794 498454 101414 533898
rect 100794 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 101414 498454
rect 100794 498134 101414 498218
rect 100794 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 101414 498134
rect 100794 462454 101414 497898
rect 100794 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 101414 462454
rect 100794 462134 101414 462218
rect 100794 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 101414 462134
rect 100794 426454 101414 461898
rect 100794 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 101414 426454
rect 100794 426134 101414 426218
rect 100794 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 101414 426134
rect 100794 390454 101414 425898
rect 100794 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 101414 390454
rect 100794 390134 101414 390218
rect 100794 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 101414 390134
rect 100794 354454 101414 389898
rect 100794 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 101414 354454
rect 100794 354134 101414 354218
rect 100794 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 101414 354134
rect 100794 318454 101414 353898
rect 100794 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 101414 318454
rect 100794 318134 101414 318218
rect 100794 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 101414 318134
rect 100794 282454 101414 317898
rect 100794 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 101414 282454
rect 100794 282134 101414 282218
rect 100794 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 101414 282134
rect 100794 246454 101414 281898
rect 100794 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 101414 246454
rect 100794 246134 101414 246218
rect 100794 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 101414 246134
rect 100794 210454 101414 245898
rect 100794 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 101414 210454
rect 100794 210134 101414 210218
rect 100794 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 101414 210134
rect 100339 193900 100405 193901
rect 100339 193836 100340 193900
rect 100404 193836 100405 193900
rect 100339 193835 100405 193836
rect 96294 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 96914 169954
rect 96294 169634 96914 169718
rect 96294 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 96914 169634
rect 96294 133954 96914 169398
rect 96294 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 96914 133954
rect 96294 133634 96914 133718
rect 96294 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 96914 133634
rect 96294 97954 96914 133398
rect 96294 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 96914 97954
rect 96294 97634 96914 97718
rect 96294 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 96914 97634
rect 96294 61954 96914 97398
rect 100342 63341 100402 193835
rect 100523 189956 100589 189957
rect 100523 189892 100524 189956
rect 100588 189892 100589 189956
rect 100523 189891 100589 189892
rect 100339 63340 100405 63341
rect 100339 63276 100340 63340
rect 100404 63276 100405 63340
rect 100339 63275 100405 63276
rect 100342 62797 100402 63275
rect 100339 62796 100405 62797
rect 100339 62732 100340 62796
rect 100404 62732 100405 62796
rect 100339 62731 100405 62732
rect 96294 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 96914 61954
rect 96294 61634 96914 61718
rect 96294 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 96914 61634
rect 96294 25954 96914 61398
rect 100526 56541 100586 189891
rect 100794 174454 101414 209898
rect 105294 711558 105914 711590
rect 105294 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 105914 711558
rect 105294 711238 105914 711322
rect 105294 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 105914 711238
rect 105294 682954 105914 711002
rect 105294 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 105914 682954
rect 105294 682634 105914 682718
rect 105294 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 105914 682634
rect 105294 646954 105914 682398
rect 105294 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 105914 646954
rect 105294 646634 105914 646718
rect 105294 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 105914 646634
rect 105294 610954 105914 646398
rect 105294 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 105914 610954
rect 105294 610634 105914 610718
rect 105294 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 105914 610634
rect 105294 574954 105914 610398
rect 105294 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 105914 574954
rect 105294 574634 105914 574718
rect 105294 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 105914 574634
rect 105294 538954 105914 574398
rect 105294 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 105914 538954
rect 105294 538634 105914 538718
rect 105294 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 105914 538634
rect 105294 502954 105914 538398
rect 105294 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 105914 502954
rect 105294 502634 105914 502718
rect 105294 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 105914 502634
rect 105294 466954 105914 502398
rect 105294 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 105914 466954
rect 105294 466634 105914 466718
rect 105294 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 105914 466634
rect 105294 430954 105914 466398
rect 105294 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 105914 430954
rect 105294 430634 105914 430718
rect 105294 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 105914 430634
rect 105294 394954 105914 430398
rect 105294 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 105914 394954
rect 105294 394634 105914 394718
rect 105294 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 105914 394634
rect 105294 358954 105914 394398
rect 105294 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 105914 358954
rect 105294 358634 105914 358718
rect 105294 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 105914 358634
rect 105294 322954 105914 358398
rect 105294 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 105914 322954
rect 105294 322634 105914 322718
rect 105294 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 105914 322634
rect 105294 286954 105914 322398
rect 105294 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 105914 286954
rect 105294 286634 105914 286718
rect 105294 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 105914 286634
rect 105294 250954 105914 286398
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109539 265300 109605 265301
rect 109539 265236 109540 265300
rect 109604 265236 109605 265300
rect 109539 265235 109605 265236
rect 109355 261084 109421 261085
rect 109355 261020 109356 261084
rect 109420 261020 109421 261084
rect 109355 261019 109421 261020
rect 105294 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 105914 250954
rect 105294 250634 105914 250718
rect 105294 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 105914 250634
rect 105294 214954 105914 250398
rect 105294 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 105914 214954
rect 105294 214634 105914 214718
rect 105294 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 105914 214634
rect 102915 197980 102981 197981
rect 102915 197916 102916 197980
rect 102980 197916 102981 197980
rect 102915 197915 102981 197916
rect 102731 194444 102797 194445
rect 102731 194380 102732 194444
rect 102796 194380 102797 194444
rect 102731 194379 102797 194380
rect 100794 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 101414 174454
rect 100794 174134 101414 174218
rect 100794 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 101414 174134
rect 100794 138454 101414 173898
rect 100794 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 101414 138454
rect 100794 138134 101414 138218
rect 100794 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 101414 138134
rect 100794 102454 101414 137898
rect 100794 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 101414 102454
rect 100794 102134 101414 102218
rect 100794 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 101414 102134
rect 100794 66454 101414 101898
rect 100794 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 101414 66454
rect 100794 66134 101414 66218
rect 100794 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 101414 66134
rect 99419 56540 99485 56541
rect 99419 56476 99420 56540
rect 99484 56476 99485 56540
rect 99419 56475 99485 56476
rect 100523 56540 100589 56541
rect 100523 56476 100524 56540
rect 100588 56476 100589 56540
rect 100523 56475 100589 56476
rect 99422 55861 99482 56475
rect 99419 55860 99485 55861
rect 99419 55796 99420 55860
rect 99484 55796 99485 55860
rect 99419 55795 99485 55796
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96294 -5146 96914 25398
rect 96294 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 96914 -5146
rect 96294 -5466 96914 -5382
rect 96294 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 96914 -5466
rect 96294 -7654 96914 -5702
rect 100794 30454 101414 65898
rect 102734 62117 102794 194379
rect 102918 68237 102978 197915
rect 104019 195668 104085 195669
rect 104019 195604 104020 195668
rect 104084 195604 104085 195668
rect 104019 195603 104085 195604
rect 103099 192540 103165 192541
rect 103099 192476 103100 192540
rect 103164 192476 103165 192540
rect 103099 192475 103165 192476
rect 103102 68917 103162 192475
rect 103099 68916 103165 68917
rect 103099 68852 103100 68916
rect 103164 68852 103165 68916
rect 103099 68851 103165 68852
rect 102915 68236 102981 68237
rect 102915 68172 102916 68236
rect 102980 68172 102981 68236
rect 102915 68171 102981 68172
rect 104022 66877 104082 195603
rect 104203 189820 104269 189821
rect 104203 189756 104204 189820
rect 104268 189756 104269 189820
rect 104203 189755 104269 189756
rect 104019 66876 104085 66877
rect 104019 66812 104020 66876
rect 104084 66812 104085 66876
rect 104019 66811 104085 66812
rect 104206 64701 104266 189755
rect 105294 178954 105914 214398
rect 106779 200564 106845 200565
rect 106779 200500 106780 200564
rect 106844 200500 106845 200564
rect 106779 200499 106845 200500
rect 105294 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 105914 178954
rect 105294 178634 105914 178718
rect 105294 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 105914 178634
rect 104387 148884 104453 148885
rect 104387 148820 104388 148884
rect 104452 148820 104453 148884
rect 104387 148819 104453 148820
rect 104203 64700 104269 64701
rect 104203 64636 104204 64700
rect 104268 64636 104269 64700
rect 104203 64635 104269 64636
rect 102731 62116 102797 62117
rect 102731 62052 102732 62116
rect 102796 62052 102797 62116
rect 102731 62051 102797 62052
rect 104390 59261 104450 148819
rect 105294 142954 105914 178398
rect 105294 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 105914 142954
rect 105294 142634 105914 142718
rect 105294 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 105914 142634
rect 105294 106954 105914 142398
rect 105294 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 105914 106954
rect 105294 106634 105914 106718
rect 105294 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 105914 106634
rect 105294 70954 105914 106398
rect 106782 74085 106842 200499
rect 107515 198388 107581 198389
rect 107515 198324 107516 198388
rect 107580 198324 107581 198388
rect 107515 198323 107581 198324
rect 106963 198116 107029 198117
rect 106963 198052 106964 198116
rect 107028 198052 107029 198116
rect 106963 198051 107029 198052
rect 106779 74084 106845 74085
rect 106779 74020 106780 74084
rect 106844 74020 106845 74084
rect 106779 74019 106845 74020
rect 106966 71093 107026 198051
rect 107518 77893 107578 198323
rect 108435 187236 108501 187237
rect 108435 187172 108436 187236
rect 108500 187172 108501 187236
rect 108435 187171 108501 187172
rect 108251 187100 108317 187101
rect 108251 187036 108252 187100
rect 108316 187036 108317 187100
rect 108251 187035 108317 187036
rect 107515 77892 107581 77893
rect 107515 77828 107516 77892
rect 107580 77828 107581 77892
rect 107515 77827 107581 77828
rect 106963 71092 107029 71093
rect 106963 71028 106964 71092
rect 107028 71028 107029 71092
rect 106963 71027 107029 71028
rect 105294 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 105914 70954
rect 105294 70634 105914 70718
rect 105294 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 105914 70634
rect 104387 59260 104453 59261
rect 104387 59196 104388 59260
rect 104452 59196 104453 59260
rect 104387 59195 104453 59196
rect 100794 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 101414 30454
rect 100794 30134 101414 30218
rect 100794 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 101414 30134
rect 100794 -6106 101414 29898
rect 100794 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 101414 -6106
rect 100794 -6426 101414 -6342
rect 100794 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 101414 -6426
rect 100794 -7654 101414 -6662
rect 105294 34954 105914 70398
rect 108254 66197 108314 187035
rect 108438 67013 108498 187171
rect 108803 151468 108869 151469
rect 108803 151404 108804 151468
rect 108868 151404 108869 151468
rect 108803 151403 108869 151404
rect 108435 67012 108501 67013
rect 108435 66948 108436 67012
rect 108500 66948 108501 67012
rect 108435 66947 108501 66948
rect 108251 66196 108317 66197
rect 108251 66132 108252 66196
rect 108316 66132 108317 66196
rect 108251 66131 108317 66132
rect 108806 65789 108866 151403
rect 109358 146301 109418 261019
rect 109355 146300 109421 146301
rect 109355 146236 109356 146300
rect 109420 146236 109421 146300
rect 109355 146235 109421 146236
rect 109542 146165 109602 265235
rect 109794 255454 110414 290898
rect 114294 705798 114914 711590
rect 114294 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 114914 705798
rect 114294 705478 114914 705562
rect 114294 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 114914 705478
rect 114294 691954 114914 705242
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 655954 114914 691398
rect 114294 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 114914 655954
rect 114294 655634 114914 655718
rect 114294 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 114914 655634
rect 114294 619954 114914 655398
rect 114294 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 114914 619954
rect 114294 619634 114914 619718
rect 114294 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 114914 619634
rect 114294 583954 114914 619398
rect 114294 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 114914 583954
rect 114294 583634 114914 583718
rect 114294 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 114914 583634
rect 114294 547954 114914 583398
rect 114294 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 114914 547954
rect 114294 547634 114914 547718
rect 114294 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 114914 547634
rect 114294 511954 114914 547398
rect 114294 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 114914 511954
rect 114294 511634 114914 511718
rect 114294 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 114914 511634
rect 114294 475954 114914 511398
rect 114294 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 114914 475954
rect 114294 475634 114914 475718
rect 114294 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 114914 475634
rect 114294 439954 114914 475398
rect 114294 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 114914 439954
rect 114294 439634 114914 439718
rect 114294 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 114914 439634
rect 114294 403954 114914 439398
rect 114294 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 114914 403954
rect 114294 403634 114914 403718
rect 114294 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 114914 403634
rect 114294 367954 114914 403398
rect 114294 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 114914 367954
rect 114294 367634 114914 367718
rect 114294 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 114914 367634
rect 114294 331954 114914 367398
rect 114294 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 114914 331954
rect 114294 331634 114914 331718
rect 114294 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 114914 331634
rect 114294 295954 114914 331398
rect 114294 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 114914 295954
rect 114294 295634 114914 295718
rect 114294 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 114914 295634
rect 112851 265028 112917 265029
rect 112851 264964 112852 265028
rect 112916 264964 112917 265028
rect 112851 264963 112917 264964
rect 111563 262580 111629 262581
rect 111563 262516 111564 262580
rect 111628 262516 111629 262580
rect 111563 262515 111629 262516
rect 111379 261220 111445 261221
rect 111379 261156 111380 261220
rect 111444 261156 111445 261220
rect 111379 261155 111445 261156
rect 111195 260948 111261 260949
rect 111195 260884 111196 260948
rect 111260 260884 111261 260948
rect 111195 260883 111261 260884
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 110827 147388 110893 147389
rect 110827 147324 110828 147388
rect 110892 147324 110893 147388
rect 110827 147323 110893 147324
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109539 146164 109605 146165
rect 109539 146100 109540 146164
rect 109604 146100 109605 146164
rect 109539 146099 109605 146100
rect 109539 138820 109605 138821
rect 109539 138756 109540 138820
rect 109604 138756 109605 138820
rect 109539 138755 109605 138756
rect 109542 66061 109602 138755
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109539 66060 109605 66061
rect 109539 65996 109540 66060
rect 109604 65996 109605 66060
rect 109539 65995 109605 65996
rect 108803 65788 108869 65789
rect 108803 65724 108804 65788
rect 108868 65724 108869 65788
rect 108803 65723 108869 65724
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 105294 -7066 105914 34398
rect 105294 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 105914 -7066
rect 105294 -7386 105914 -7302
rect 105294 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 105914 -7386
rect 105294 -7654 105914 -7622
rect 109794 39454 110414 74898
rect 110830 65925 110890 147323
rect 111198 145485 111258 260883
rect 111195 145484 111261 145485
rect 111195 145420 111196 145484
rect 111260 145420 111261 145484
rect 111195 145419 111261 145420
rect 111382 143309 111442 261155
rect 111566 144397 111626 262515
rect 112299 147524 112365 147525
rect 112299 147460 112300 147524
rect 112364 147460 112365 147524
rect 112299 147459 112365 147460
rect 111563 144396 111629 144397
rect 111563 144332 111564 144396
rect 111628 144332 111629 144396
rect 111563 144331 111629 144332
rect 111379 143308 111445 143309
rect 111379 143244 111380 143308
rect 111444 143244 111445 143308
rect 111379 143243 111445 143244
rect 111011 142492 111077 142493
rect 111011 142428 111012 142492
rect 111076 142428 111077 142492
rect 111011 142427 111077 142428
rect 110827 65924 110893 65925
rect 110827 65860 110828 65924
rect 110892 65860 110893 65924
rect 110827 65859 110893 65860
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 111014 10301 111074 142427
rect 111195 139364 111261 139365
rect 111195 139300 111196 139364
rect 111260 139300 111261 139364
rect 111195 139299 111261 139300
rect 111198 76669 111258 139299
rect 111195 76668 111261 76669
rect 111195 76604 111196 76668
rect 111260 76604 111261 76668
rect 111195 76603 111261 76604
rect 112302 60621 112362 147459
rect 112667 147116 112733 147117
rect 112667 147052 112668 147116
rect 112732 147052 112733 147116
rect 112667 147051 112733 147052
rect 112670 75309 112730 147051
rect 112854 145621 112914 264963
rect 114139 262852 114205 262853
rect 114139 262788 114140 262852
rect 114204 262788 114205 262852
rect 114139 262787 114205 262788
rect 113035 196620 113101 196621
rect 113035 196556 113036 196620
rect 113100 196556 113101 196620
rect 113035 196555 113101 196556
rect 112851 145620 112917 145621
rect 112851 145556 112852 145620
rect 112916 145556 112917 145620
rect 112851 145555 112917 145556
rect 112851 141676 112917 141677
rect 112851 141612 112852 141676
rect 112916 141612 112917 141676
rect 112851 141611 112917 141612
rect 112667 75308 112733 75309
rect 112667 75244 112668 75308
rect 112732 75244 112733 75308
rect 112667 75243 112733 75244
rect 112854 65653 112914 141611
rect 113038 75717 113098 196555
rect 113403 149836 113469 149837
rect 113403 149772 113404 149836
rect 113468 149772 113469 149836
rect 113403 149771 113469 149772
rect 113035 75716 113101 75717
rect 113035 75652 113036 75716
rect 113100 75652 113101 75716
rect 113035 75651 113101 75652
rect 113406 67421 113466 149771
rect 113587 148340 113653 148341
rect 113587 148276 113588 148340
rect 113652 148276 113653 148340
rect 113587 148275 113653 148276
rect 113590 74357 113650 148275
rect 113955 146844 114021 146845
rect 113955 146780 113956 146844
rect 114020 146780 114021 146844
rect 113955 146779 114021 146780
rect 113771 138004 113837 138005
rect 113771 137940 113772 138004
rect 113836 137940 113837 138004
rect 113771 137939 113837 137940
rect 113587 74356 113653 74357
rect 113587 74292 113588 74356
rect 113652 74292 113653 74356
rect 113587 74291 113653 74292
rect 113403 67420 113469 67421
rect 113403 67356 113404 67420
rect 113468 67356 113469 67420
rect 113403 67355 113469 67356
rect 112851 65652 112917 65653
rect 112851 65588 112852 65652
rect 112916 65588 112917 65652
rect 112851 65587 112917 65588
rect 112299 60620 112365 60621
rect 112299 60556 112300 60620
rect 112364 60556 112365 60620
rect 112299 60555 112365 60556
rect 113774 55997 113834 137939
rect 113958 70141 114018 146779
rect 114142 144669 114202 262787
rect 114294 259954 114914 295398
rect 118794 706758 119414 711590
rect 118794 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 119414 706758
rect 118794 706438 119414 706522
rect 118794 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 119414 706438
rect 118794 696454 119414 706202
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 660454 119414 695898
rect 118794 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 119414 660454
rect 118794 660134 119414 660218
rect 118794 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 119414 660134
rect 118794 624454 119414 659898
rect 118794 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 119414 624454
rect 118794 624134 119414 624218
rect 118794 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 119414 624134
rect 118794 588454 119414 623898
rect 118794 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 119414 588454
rect 118794 588134 119414 588218
rect 118794 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 119414 588134
rect 118794 552454 119414 587898
rect 118794 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 119414 552454
rect 118794 552134 119414 552218
rect 118794 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 119414 552134
rect 118794 516454 119414 551898
rect 118794 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 119414 516454
rect 118794 516134 119414 516218
rect 118794 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 119414 516134
rect 118794 480454 119414 515898
rect 118794 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 119414 480454
rect 118794 480134 119414 480218
rect 118794 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 119414 480134
rect 118794 444454 119414 479898
rect 118794 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 119414 444454
rect 118794 444134 119414 444218
rect 118794 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 119414 444134
rect 118794 408454 119414 443898
rect 118794 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 119414 408454
rect 118794 408134 119414 408218
rect 118794 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 119414 408134
rect 118794 372454 119414 407898
rect 118794 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 119414 372454
rect 118794 372134 119414 372218
rect 118794 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 119414 372134
rect 118794 336454 119414 371898
rect 118794 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 119414 336454
rect 118794 336134 119414 336218
rect 118794 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 119414 336134
rect 118794 300454 119414 335898
rect 118794 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 119414 300454
rect 118794 300134 119414 300218
rect 118794 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 119414 300134
rect 115795 265164 115861 265165
rect 115795 265100 115796 265164
rect 115860 265100 115861 265164
rect 115795 265099 115861 265100
rect 114294 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 114914 259954
rect 114294 259634 114914 259718
rect 114294 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 114914 259634
rect 114294 223954 114914 259398
rect 114294 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 114914 223954
rect 114294 223634 114914 223718
rect 114294 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 114914 223634
rect 114294 187954 114914 223398
rect 114294 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 114914 187954
rect 114294 187634 114914 187718
rect 114294 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 114914 187634
rect 114294 151954 114914 187398
rect 114294 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 114914 151954
rect 114294 151634 114914 151718
rect 114294 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 114914 151634
rect 114139 144668 114205 144669
rect 114139 144604 114140 144668
rect 114204 144604 114205 144668
rect 114139 144603 114205 144604
rect 114294 115954 114914 151398
rect 115427 148612 115493 148613
rect 115427 148548 115428 148612
rect 115492 148548 115493 148612
rect 115427 148547 115493 148548
rect 115059 147252 115125 147253
rect 115059 147188 115060 147252
rect 115124 147188 115125 147252
rect 115059 147187 115125 147188
rect 115062 139365 115122 147187
rect 115059 139364 115125 139365
rect 115059 139300 115060 139364
rect 115124 139300 115125 139364
rect 115059 139299 115125 139300
rect 114294 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 114914 115954
rect 114294 115634 114914 115718
rect 114294 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 114914 115634
rect 114294 79954 114914 115398
rect 114294 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 114914 79954
rect 114294 79634 114914 79718
rect 114294 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 114914 79634
rect 113955 70140 114021 70141
rect 113955 70076 113956 70140
rect 114020 70076 114021 70140
rect 113955 70075 114021 70076
rect 114139 67420 114205 67421
rect 114139 67356 114140 67420
rect 114204 67356 114205 67420
rect 114139 67355 114205 67356
rect 113771 55996 113837 55997
rect 113771 55932 113772 55996
rect 113836 55932 113837 55996
rect 113771 55931 113837 55932
rect 114142 52597 114202 67355
rect 114139 52596 114205 52597
rect 114139 52532 114140 52596
rect 114204 52532 114205 52596
rect 114139 52531 114205 52532
rect 114294 43954 114914 79398
rect 115430 71637 115490 148547
rect 115798 145893 115858 265099
rect 118794 264454 119414 299898
rect 118794 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 119414 264454
rect 118794 264134 119414 264218
rect 118794 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 119414 264134
rect 123294 707718 123914 711590
rect 123294 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 123914 707718
rect 123294 707398 123914 707482
rect 123294 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 123914 707398
rect 123294 700954 123914 707162
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 664954 123914 700398
rect 123294 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 123914 664954
rect 123294 664634 123914 664718
rect 123294 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 123914 664634
rect 123294 628954 123914 664398
rect 123294 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 123914 628954
rect 123294 628634 123914 628718
rect 123294 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 123914 628634
rect 123294 592954 123914 628398
rect 123294 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 123914 592954
rect 123294 592634 123914 592718
rect 123294 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 123914 592634
rect 123294 556954 123914 592398
rect 123294 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 123914 556954
rect 123294 556634 123914 556718
rect 123294 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 123914 556634
rect 123294 520954 123914 556398
rect 123294 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 123914 520954
rect 123294 520634 123914 520718
rect 123294 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 123914 520634
rect 123294 484954 123914 520398
rect 123294 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 123914 484954
rect 123294 484634 123914 484718
rect 123294 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 123914 484634
rect 123294 448954 123914 484398
rect 123294 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 123914 448954
rect 123294 448634 123914 448718
rect 123294 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 123914 448634
rect 123294 412954 123914 448398
rect 123294 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 123914 412954
rect 123294 412634 123914 412718
rect 123294 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 123914 412634
rect 123294 376954 123914 412398
rect 123294 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 123914 376954
rect 123294 376634 123914 376718
rect 123294 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 123914 376634
rect 123294 340954 123914 376398
rect 123294 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 123914 340954
rect 123294 340634 123914 340718
rect 123294 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 123914 340634
rect 123294 304954 123914 340398
rect 123294 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 123914 304954
rect 123294 304634 123914 304718
rect 123294 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 123914 304634
rect 123294 268954 123914 304398
rect 123294 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 123914 268954
rect 123294 268634 123914 268718
rect 123294 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 123914 268634
rect 118371 263668 118437 263669
rect 118371 263604 118372 263668
rect 118436 263604 118437 263668
rect 118371 263603 118437 263604
rect 116899 259996 116965 259997
rect 116899 259932 116900 259996
rect 116964 259932 116965 259996
rect 116899 259931 116965 259932
rect 116715 259588 116781 259589
rect 116715 259524 116716 259588
rect 116780 259524 116781 259588
rect 116715 259523 116781 259524
rect 116163 146028 116229 146029
rect 116163 145964 116164 146028
rect 116228 145964 116229 146028
rect 116163 145963 116229 145964
rect 115795 145892 115861 145893
rect 115795 145828 115796 145892
rect 115860 145828 115861 145892
rect 115795 145827 115861 145828
rect 115611 142900 115677 142901
rect 115611 142836 115612 142900
rect 115676 142836 115677 142900
rect 115611 142835 115677 142836
rect 115427 71636 115493 71637
rect 115427 71572 115428 71636
rect 115492 71572 115493 71636
rect 115427 71571 115493 71572
rect 115614 67421 115674 142835
rect 116166 71773 116226 145963
rect 116347 144260 116413 144261
rect 116347 144196 116348 144260
rect 116412 144196 116413 144260
rect 116347 144195 116413 144196
rect 116163 71772 116229 71773
rect 116163 71708 116164 71772
rect 116228 71708 116229 71772
rect 116163 71707 116229 71708
rect 116350 68645 116410 144195
rect 116718 143989 116778 259523
rect 116715 143988 116781 143989
rect 116715 143924 116716 143988
rect 116780 143924 116781 143988
rect 116715 143923 116781 143924
rect 116902 141949 116962 259931
rect 117083 200836 117149 200837
rect 117083 200772 117084 200836
rect 117148 200772 117149 200836
rect 117083 200771 117149 200772
rect 116899 141948 116965 141949
rect 116899 141884 116900 141948
rect 116964 141884 116965 141948
rect 116899 141883 116965 141884
rect 116531 139772 116597 139773
rect 116531 139708 116532 139772
rect 116596 139708 116597 139772
rect 116531 139707 116597 139708
rect 116347 68644 116413 68645
rect 116347 68580 116348 68644
rect 116412 68580 116413 68644
rect 116347 68579 116413 68580
rect 115611 67420 115677 67421
rect 115611 67356 115612 67420
rect 115676 67356 115677 67420
rect 115611 67355 115677 67356
rect 116534 44301 116594 139707
rect 117086 74493 117146 200771
rect 117819 148476 117885 148477
rect 117819 148412 117820 148476
rect 117884 148412 117885 148476
rect 117819 148411 117885 148412
rect 117083 74492 117149 74493
rect 117083 74428 117084 74492
rect 117148 74428 117149 74492
rect 117083 74427 117149 74428
rect 117822 70277 117882 148411
rect 118374 142765 118434 263603
rect 118794 262000 119414 263898
rect 121131 263940 121197 263941
rect 121131 263876 121132 263940
rect 121196 263876 121197 263940
rect 121131 263875 121197 263876
rect 118555 199340 118621 199341
rect 118555 199276 118556 199340
rect 118620 199276 118621 199340
rect 118555 199275 118621 199276
rect 118371 142764 118437 142765
rect 118371 142700 118372 142764
rect 118436 142700 118437 142764
rect 118371 142699 118437 142700
rect 118187 141404 118253 141405
rect 118187 141340 118188 141404
rect 118252 141340 118253 141404
rect 118187 141339 118253 141340
rect 118003 139228 118069 139229
rect 118003 139164 118004 139228
rect 118068 139164 118069 139228
rect 118003 139163 118069 139164
rect 117819 70276 117885 70277
rect 117819 70212 117820 70276
rect 117884 70212 117885 70276
rect 117819 70211 117885 70212
rect 118006 68917 118066 139163
rect 118003 68916 118069 68917
rect 118003 68852 118004 68916
rect 118068 68852 118069 68916
rect 118003 68851 118069 68852
rect 118190 68781 118250 141339
rect 118558 73949 118618 199275
rect 118794 192454 119414 198000
rect 119843 195260 119909 195261
rect 119843 195196 119844 195260
rect 119908 195196 119909 195260
rect 119843 195195 119909 195196
rect 118794 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 119414 192454
rect 118794 192134 119414 192218
rect 118794 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 119414 192134
rect 118794 156454 119414 191898
rect 118794 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 119414 156454
rect 118794 156134 119414 156218
rect 118794 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 119414 156134
rect 118794 142000 119414 155898
rect 119659 145756 119725 145757
rect 119659 145692 119660 145756
rect 119724 145692 119725 145756
rect 119659 145691 119725 145692
rect 118739 140724 118805 140725
rect 118739 140660 118740 140724
rect 118804 140660 118805 140724
rect 118739 140659 118805 140660
rect 118742 96661 118802 140659
rect 119475 140452 119541 140453
rect 119475 140388 119476 140452
rect 119540 140388 119541 140452
rect 119475 140387 119541 140388
rect 118739 96660 118805 96661
rect 118739 96596 118740 96660
rect 118804 96596 118805 96660
rect 118739 96595 118805 96596
rect 119478 78570 119538 140387
rect 119662 79253 119722 145691
rect 119659 79252 119725 79253
rect 119659 79188 119660 79252
rect 119724 79188 119725 79252
rect 119659 79187 119725 79188
rect 119478 78510 119722 78570
rect 118555 73948 118621 73949
rect 118555 73884 118556 73948
rect 118620 73884 118621 73948
rect 118555 73883 118621 73884
rect 118187 68780 118253 68781
rect 118187 68716 118188 68780
rect 118252 68716 118253 68780
rect 118187 68715 118253 68716
rect 118794 48454 119414 78000
rect 119662 77213 119722 78510
rect 119659 77212 119725 77213
rect 119659 77148 119660 77212
rect 119724 77148 119725 77212
rect 119659 77147 119725 77148
rect 119659 75852 119725 75853
rect 119659 75788 119660 75852
rect 119724 75850 119725 75852
rect 119846 75850 119906 195195
rect 120763 148748 120829 148749
rect 120763 148684 120764 148748
rect 120828 148684 120829 148748
rect 120763 148683 120829 148684
rect 119724 75790 119906 75850
rect 119724 75788 119725 75790
rect 119659 75787 119725 75788
rect 119662 75173 119722 75787
rect 119659 75172 119725 75173
rect 119659 75108 119660 75172
rect 119724 75108 119725 75172
rect 119659 75107 119725 75108
rect 120766 70005 120826 148683
rect 121134 143037 121194 263875
rect 121315 263804 121381 263805
rect 121315 263740 121316 263804
rect 121380 263740 121381 263804
rect 121315 263739 121381 263740
rect 121318 143173 121378 263739
rect 123294 262000 123914 268398
rect 127794 708678 128414 711590
rect 127794 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 128414 708678
rect 127794 708358 128414 708442
rect 127794 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 128414 708358
rect 127794 669454 128414 708122
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 262000 128414 272898
rect 132294 709638 132914 711590
rect 132294 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 132914 709638
rect 132294 709318 132914 709402
rect 132294 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 132914 709318
rect 132294 673954 132914 709082
rect 132294 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 132914 673954
rect 132294 673634 132914 673718
rect 132294 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 132914 673634
rect 132294 637954 132914 673398
rect 132294 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 132914 637954
rect 132294 637634 132914 637718
rect 132294 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 132914 637634
rect 132294 601954 132914 637398
rect 132294 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 132914 601954
rect 132294 601634 132914 601718
rect 132294 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 132914 601634
rect 132294 565954 132914 601398
rect 132294 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 132914 565954
rect 132294 565634 132914 565718
rect 132294 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 132914 565634
rect 132294 529954 132914 565398
rect 132294 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 132914 529954
rect 132294 529634 132914 529718
rect 132294 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 132914 529634
rect 132294 493954 132914 529398
rect 132294 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 132914 493954
rect 132294 493634 132914 493718
rect 132294 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 132914 493634
rect 132294 457954 132914 493398
rect 132294 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 132914 457954
rect 132294 457634 132914 457718
rect 132294 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 132914 457634
rect 132294 421954 132914 457398
rect 132294 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 132914 421954
rect 132294 421634 132914 421718
rect 132294 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 132914 421634
rect 132294 385954 132914 421398
rect 132294 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 132914 385954
rect 132294 385634 132914 385718
rect 132294 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 132914 385634
rect 132294 349954 132914 385398
rect 132294 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 132914 349954
rect 132294 349634 132914 349718
rect 132294 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 132914 349634
rect 132294 313954 132914 349398
rect 132294 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 132914 313954
rect 132294 313634 132914 313718
rect 132294 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 132914 313634
rect 132294 277954 132914 313398
rect 132294 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 132914 277954
rect 132294 277634 132914 277718
rect 132294 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 132914 277634
rect 132294 262000 132914 277398
rect 136794 710598 137414 711590
rect 136794 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 137414 710598
rect 136794 710278 137414 710362
rect 136794 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 137414 710278
rect 136794 678454 137414 710042
rect 136794 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 137414 678454
rect 136794 678134 137414 678218
rect 136794 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 137414 678134
rect 136794 642454 137414 677898
rect 136794 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 137414 642454
rect 136794 642134 137414 642218
rect 136794 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 137414 642134
rect 136794 606454 137414 641898
rect 136794 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 137414 606454
rect 136794 606134 137414 606218
rect 136794 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 137414 606134
rect 136794 570454 137414 605898
rect 136794 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 137414 570454
rect 136794 570134 137414 570218
rect 136794 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 137414 570134
rect 136794 534454 137414 569898
rect 136794 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 137414 534454
rect 136794 534134 137414 534218
rect 136794 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 137414 534134
rect 136794 498454 137414 533898
rect 136794 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 137414 498454
rect 136794 498134 137414 498218
rect 136794 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 137414 498134
rect 136794 462454 137414 497898
rect 136794 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 137414 462454
rect 136794 462134 137414 462218
rect 136794 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 137414 462134
rect 136794 426454 137414 461898
rect 136794 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 137414 426454
rect 136794 426134 137414 426218
rect 136794 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 137414 426134
rect 136794 390454 137414 425898
rect 136794 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 137414 390454
rect 136794 390134 137414 390218
rect 136794 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 137414 390134
rect 136794 354454 137414 389898
rect 136794 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 137414 354454
rect 136794 354134 137414 354218
rect 136794 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 137414 354134
rect 136794 318454 137414 353898
rect 136794 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 137414 318454
rect 136794 318134 137414 318218
rect 136794 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 137414 318134
rect 136794 282454 137414 317898
rect 136794 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 137414 282454
rect 136794 282134 137414 282218
rect 136794 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 137414 282134
rect 136794 262000 137414 281898
rect 141294 711558 141914 711590
rect 141294 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 141914 711558
rect 141294 711238 141914 711322
rect 141294 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 141914 711238
rect 141294 682954 141914 711002
rect 141294 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 141914 682954
rect 141294 682634 141914 682718
rect 141294 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 141914 682634
rect 141294 646954 141914 682398
rect 141294 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 141914 646954
rect 141294 646634 141914 646718
rect 141294 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 141914 646634
rect 141294 610954 141914 646398
rect 141294 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 141914 610954
rect 141294 610634 141914 610718
rect 141294 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 141914 610634
rect 141294 574954 141914 610398
rect 141294 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 141914 574954
rect 141294 574634 141914 574718
rect 141294 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 141914 574634
rect 141294 538954 141914 574398
rect 141294 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 141914 538954
rect 141294 538634 141914 538718
rect 141294 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 141914 538634
rect 141294 502954 141914 538398
rect 141294 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 141914 502954
rect 141294 502634 141914 502718
rect 141294 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 141914 502634
rect 141294 466954 141914 502398
rect 141294 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 141914 466954
rect 141294 466634 141914 466718
rect 141294 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 141914 466634
rect 141294 430954 141914 466398
rect 141294 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 141914 430954
rect 141294 430634 141914 430718
rect 141294 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 141914 430634
rect 141294 394954 141914 430398
rect 141294 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 141914 394954
rect 141294 394634 141914 394718
rect 141294 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 141914 394634
rect 141294 358954 141914 394398
rect 141294 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 141914 358954
rect 141294 358634 141914 358718
rect 141294 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 141914 358634
rect 141294 322954 141914 358398
rect 141294 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 141914 322954
rect 141294 322634 141914 322718
rect 141294 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 141914 322634
rect 141294 286954 141914 322398
rect 141294 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 141914 286954
rect 141294 286634 141914 286718
rect 141294 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 141914 286634
rect 141294 262000 141914 286398
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 262000 146414 290898
rect 150294 705798 150914 711590
rect 150294 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 150914 705798
rect 150294 705478 150914 705562
rect 150294 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 150914 705478
rect 150294 691954 150914 705242
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 655954 150914 691398
rect 150294 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 150914 655954
rect 150294 655634 150914 655718
rect 150294 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 150914 655634
rect 150294 619954 150914 655398
rect 150294 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 150914 619954
rect 150294 619634 150914 619718
rect 150294 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 150914 619634
rect 150294 583954 150914 619398
rect 150294 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 150914 583954
rect 150294 583634 150914 583718
rect 150294 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 150914 583634
rect 150294 547954 150914 583398
rect 150294 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 150914 547954
rect 150294 547634 150914 547718
rect 150294 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 150914 547634
rect 150294 511954 150914 547398
rect 150294 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 150914 511954
rect 150294 511634 150914 511718
rect 150294 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 150914 511634
rect 150294 475954 150914 511398
rect 150294 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 150914 475954
rect 150294 475634 150914 475718
rect 150294 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 150914 475634
rect 150294 439954 150914 475398
rect 150294 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 150914 439954
rect 150294 439634 150914 439718
rect 150294 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 150914 439634
rect 150294 403954 150914 439398
rect 150294 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 150914 403954
rect 150294 403634 150914 403718
rect 150294 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 150914 403634
rect 150294 367954 150914 403398
rect 150294 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 150914 367954
rect 150294 367634 150914 367718
rect 150294 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 150914 367634
rect 150294 331954 150914 367398
rect 150294 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 150914 331954
rect 150294 331634 150914 331718
rect 150294 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 150914 331634
rect 150294 295954 150914 331398
rect 150294 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 150914 295954
rect 150294 295634 150914 295718
rect 150294 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 150914 295634
rect 150294 262000 150914 295398
rect 154794 706758 155414 711590
rect 154794 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 155414 706758
rect 154794 706438 155414 706522
rect 154794 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 155414 706438
rect 154794 696454 155414 706202
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 660454 155414 695898
rect 154794 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 155414 660454
rect 154794 660134 155414 660218
rect 154794 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 155414 660134
rect 154794 624454 155414 659898
rect 154794 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 155414 624454
rect 154794 624134 155414 624218
rect 154794 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 155414 624134
rect 154794 588454 155414 623898
rect 154794 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 155414 588454
rect 154794 588134 155414 588218
rect 154794 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 155414 588134
rect 154794 552454 155414 587898
rect 154794 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 155414 552454
rect 154794 552134 155414 552218
rect 154794 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 155414 552134
rect 154794 516454 155414 551898
rect 154794 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 155414 516454
rect 154794 516134 155414 516218
rect 154794 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 155414 516134
rect 154794 480454 155414 515898
rect 154794 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 155414 480454
rect 154794 480134 155414 480218
rect 154794 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 155414 480134
rect 154794 444454 155414 479898
rect 154794 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 155414 444454
rect 154794 444134 155414 444218
rect 154794 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 155414 444134
rect 154794 408454 155414 443898
rect 154794 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 155414 408454
rect 154794 408134 155414 408218
rect 154794 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 155414 408134
rect 154794 372454 155414 407898
rect 154794 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 155414 372454
rect 154794 372134 155414 372218
rect 154794 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 155414 372134
rect 154794 336454 155414 371898
rect 154794 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 155414 336454
rect 154794 336134 155414 336218
rect 154794 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 155414 336134
rect 154794 300454 155414 335898
rect 154794 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 155414 300454
rect 154794 300134 155414 300218
rect 154794 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 155414 300134
rect 154794 264454 155414 299898
rect 154794 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 155414 264454
rect 154794 264134 155414 264218
rect 154794 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 155414 264134
rect 154794 262000 155414 263898
rect 159294 707718 159914 711590
rect 159294 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 159914 707718
rect 159294 707398 159914 707482
rect 159294 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 159914 707398
rect 159294 700954 159914 707162
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 664954 159914 700398
rect 159294 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 159914 664954
rect 159294 664634 159914 664718
rect 159294 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 159914 664634
rect 159294 628954 159914 664398
rect 159294 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 159914 628954
rect 159294 628634 159914 628718
rect 159294 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 159914 628634
rect 159294 592954 159914 628398
rect 159294 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 159914 592954
rect 159294 592634 159914 592718
rect 159294 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 159914 592634
rect 159294 556954 159914 592398
rect 159294 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 159914 556954
rect 159294 556634 159914 556718
rect 159294 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 159914 556634
rect 159294 520954 159914 556398
rect 159294 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 159914 520954
rect 159294 520634 159914 520718
rect 159294 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 159914 520634
rect 159294 484954 159914 520398
rect 159294 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 159914 484954
rect 159294 484634 159914 484718
rect 159294 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 159914 484634
rect 159294 448954 159914 484398
rect 159294 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 159914 448954
rect 159294 448634 159914 448718
rect 159294 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 159914 448634
rect 159294 412954 159914 448398
rect 159294 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 159914 412954
rect 159294 412634 159914 412718
rect 159294 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 159914 412634
rect 159294 376954 159914 412398
rect 159294 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 159914 376954
rect 159294 376634 159914 376718
rect 159294 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 159914 376634
rect 159294 340954 159914 376398
rect 159294 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 159914 340954
rect 159294 340634 159914 340718
rect 159294 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 159914 340634
rect 159294 304954 159914 340398
rect 159294 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 159914 304954
rect 159294 304634 159914 304718
rect 159294 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 159914 304634
rect 159294 268954 159914 304398
rect 159294 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 159914 268954
rect 159294 268634 159914 268718
rect 159294 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 159914 268634
rect 159294 262000 159914 268398
rect 163794 708678 164414 711590
rect 163794 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 164414 708678
rect 163794 708358 164414 708442
rect 163794 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 164414 708358
rect 163794 669454 164414 708122
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 262000 164414 272898
rect 168294 709638 168914 711590
rect 168294 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 168914 709638
rect 168294 709318 168914 709402
rect 168294 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 168914 709318
rect 168294 673954 168914 709082
rect 168294 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 168914 673954
rect 168294 673634 168914 673718
rect 168294 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 168914 673634
rect 168294 637954 168914 673398
rect 168294 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 168914 637954
rect 168294 637634 168914 637718
rect 168294 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 168914 637634
rect 168294 601954 168914 637398
rect 168294 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 168914 601954
rect 168294 601634 168914 601718
rect 168294 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 168914 601634
rect 168294 565954 168914 601398
rect 168294 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 168914 565954
rect 168294 565634 168914 565718
rect 168294 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 168914 565634
rect 168294 529954 168914 565398
rect 168294 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 168914 529954
rect 168294 529634 168914 529718
rect 168294 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 168914 529634
rect 168294 493954 168914 529398
rect 168294 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 168914 493954
rect 168294 493634 168914 493718
rect 168294 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 168914 493634
rect 168294 457954 168914 493398
rect 168294 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 168914 457954
rect 168294 457634 168914 457718
rect 168294 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 168914 457634
rect 168294 421954 168914 457398
rect 168294 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 168914 421954
rect 168294 421634 168914 421718
rect 168294 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 168914 421634
rect 168294 385954 168914 421398
rect 168294 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 168914 385954
rect 168294 385634 168914 385718
rect 168294 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 168914 385634
rect 168294 349954 168914 385398
rect 168294 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 168914 349954
rect 168294 349634 168914 349718
rect 168294 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 168914 349634
rect 168294 313954 168914 349398
rect 168294 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 168914 313954
rect 168294 313634 168914 313718
rect 168294 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 168914 313634
rect 168294 277954 168914 313398
rect 168294 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 168914 277954
rect 168294 277634 168914 277718
rect 168294 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 168914 277634
rect 168294 262000 168914 277398
rect 172794 710598 173414 711590
rect 172794 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 173414 710598
rect 172794 710278 173414 710362
rect 172794 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 173414 710278
rect 172794 678454 173414 710042
rect 172794 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 173414 678454
rect 172794 678134 173414 678218
rect 172794 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 173414 678134
rect 172794 642454 173414 677898
rect 172794 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 173414 642454
rect 172794 642134 173414 642218
rect 172794 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 173414 642134
rect 172794 606454 173414 641898
rect 172794 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 173414 606454
rect 172794 606134 173414 606218
rect 172794 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 173414 606134
rect 172794 570454 173414 605898
rect 172794 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 173414 570454
rect 172794 570134 173414 570218
rect 172794 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 173414 570134
rect 172794 534454 173414 569898
rect 172794 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 173414 534454
rect 172794 534134 173414 534218
rect 172794 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 173414 534134
rect 172794 498454 173414 533898
rect 172794 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 173414 498454
rect 172794 498134 173414 498218
rect 172794 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 173414 498134
rect 172794 462454 173414 497898
rect 172794 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 173414 462454
rect 172794 462134 173414 462218
rect 172794 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 173414 462134
rect 172794 426454 173414 461898
rect 172794 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 173414 426454
rect 172794 426134 173414 426218
rect 172794 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 173414 426134
rect 172794 390454 173414 425898
rect 172794 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 173414 390454
rect 172794 390134 173414 390218
rect 172794 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 173414 390134
rect 172794 354454 173414 389898
rect 172794 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 173414 354454
rect 172794 354134 173414 354218
rect 172794 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 173414 354134
rect 172794 318454 173414 353898
rect 172794 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 173414 318454
rect 172794 318134 173414 318218
rect 172794 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 173414 318134
rect 172794 282454 173414 317898
rect 172794 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 173414 282454
rect 172794 282134 173414 282218
rect 172794 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 173414 282134
rect 172794 262000 173414 281898
rect 177294 711558 177914 711590
rect 177294 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 177914 711558
rect 177294 711238 177914 711322
rect 177294 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 177914 711238
rect 177294 682954 177914 711002
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 177294 646954 177914 682398
rect 177294 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 177914 646954
rect 177294 646634 177914 646718
rect 177294 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 177914 646634
rect 177294 610954 177914 646398
rect 177294 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 177914 610954
rect 177294 610634 177914 610718
rect 177294 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 177914 610634
rect 177294 574954 177914 610398
rect 177294 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 177914 574954
rect 177294 574634 177914 574718
rect 177294 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 177914 574634
rect 177294 538954 177914 574398
rect 177294 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 177914 538954
rect 177294 538634 177914 538718
rect 177294 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 177914 538634
rect 177294 502954 177914 538398
rect 177294 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 177914 502954
rect 177294 502634 177914 502718
rect 177294 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 177914 502634
rect 177294 466954 177914 502398
rect 177294 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 177914 466954
rect 177294 466634 177914 466718
rect 177294 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 177914 466634
rect 177294 430954 177914 466398
rect 177294 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 177914 430954
rect 177294 430634 177914 430718
rect 177294 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 177914 430634
rect 177294 394954 177914 430398
rect 177294 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 177914 394954
rect 177294 394634 177914 394718
rect 177294 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 177914 394634
rect 177294 358954 177914 394398
rect 177294 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 177914 358954
rect 177294 358634 177914 358718
rect 177294 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 177914 358634
rect 177294 322954 177914 358398
rect 177294 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 177914 322954
rect 177294 322634 177914 322718
rect 177294 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 177914 322634
rect 177294 286954 177914 322398
rect 177294 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 177914 286954
rect 177294 286634 177914 286718
rect 177294 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 177914 286634
rect 177294 262000 177914 286398
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 262000 182414 290898
rect 186294 705798 186914 711590
rect 186294 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 186914 705798
rect 186294 705478 186914 705562
rect 186294 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 186914 705478
rect 186294 691954 186914 705242
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 655954 186914 691398
rect 186294 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 186914 655954
rect 186294 655634 186914 655718
rect 186294 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 186914 655634
rect 186294 619954 186914 655398
rect 186294 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 186914 619954
rect 186294 619634 186914 619718
rect 186294 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 186914 619634
rect 186294 583954 186914 619398
rect 186294 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 186914 583954
rect 186294 583634 186914 583718
rect 186294 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 186914 583634
rect 186294 547954 186914 583398
rect 186294 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 186914 547954
rect 186294 547634 186914 547718
rect 186294 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 186914 547634
rect 186294 511954 186914 547398
rect 186294 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 186914 511954
rect 186294 511634 186914 511718
rect 186294 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 186914 511634
rect 186294 475954 186914 511398
rect 186294 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 186914 475954
rect 186294 475634 186914 475718
rect 186294 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 186914 475634
rect 186294 439954 186914 475398
rect 186294 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 186914 439954
rect 186294 439634 186914 439718
rect 186294 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 186914 439634
rect 186294 403954 186914 439398
rect 186294 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 186914 403954
rect 186294 403634 186914 403718
rect 186294 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 186914 403634
rect 186294 367954 186914 403398
rect 186294 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 186914 367954
rect 186294 367634 186914 367718
rect 186294 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 186914 367634
rect 186294 331954 186914 367398
rect 186294 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 186914 331954
rect 186294 331634 186914 331718
rect 186294 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 186914 331634
rect 186294 295954 186914 331398
rect 186294 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 186914 295954
rect 186294 295634 186914 295718
rect 186294 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 186914 295634
rect 186294 262000 186914 295398
rect 190794 706758 191414 711590
rect 190794 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 191414 706758
rect 190794 706438 191414 706522
rect 190794 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 191414 706438
rect 190794 696454 191414 706202
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 660454 191414 695898
rect 190794 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 191414 660454
rect 190794 660134 191414 660218
rect 190794 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 191414 660134
rect 190794 624454 191414 659898
rect 190794 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 191414 624454
rect 190794 624134 191414 624218
rect 190794 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 191414 624134
rect 190794 588454 191414 623898
rect 190794 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 191414 588454
rect 190794 588134 191414 588218
rect 190794 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 191414 588134
rect 190794 552454 191414 587898
rect 190794 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 191414 552454
rect 190794 552134 191414 552218
rect 190794 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 191414 552134
rect 190794 516454 191414 551898
rect 190794 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 191414 516454
rect 190794 516134 191414 516218
rect 190794 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 191414 516134
rect 190794 480454 191414 515898
rect 190794 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 191414 480454
rect 190794 480134 191414 480218
rect 190794 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 191414 480134
rect 190794 444454 191414 479898
rect 190794 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 191414 444454
rect 190794 444134 191414 444218
rect 190794 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 191414 444134
rect 190794 408454 191414 443898
rect 190794 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 191414 408454
rect 190794 408134 191414 408218
rect 190794 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 191414 408134
rect 190794 372454 191414 407898
rect 190794 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 191414 372454
rect 190794 372134 191414 372218
rect 190794 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 191414 372134
rect 190794 336454 191414 371898
rect 190794 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 191414 336454
rect 190794 336134 191414 336218
rect 190794 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 191414 336134
rect 190794 300454 191414 335898
rect 190794 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 191414 300454
rect 190794 300134 191414 300218
rect 190794 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 191414 300134
rect 187739 274684 187805 274685
rect 187739 274620 187740 274684
rect 187804 274620 187805 274684
rect 187739 274619 187805 274620
rect 186083 259588 186149 259589
rect 186083 259524 186084 259588
rect 186148 259524 186149 259588
rect 186083 259523 186149 259524
rect 124208 255454 124528 255486
rect 124208 255218 124250 255454
rect 124486 255218 124528 255454
rect 124208 255134 124528 255218
rect 124208 254898 124250 255134
rect 124486 254898 124528 255134
rect 124208 254866 124528 254898
rect 154928 255454 155248 255486
rect 154928 255218 154970 255454
rect 155206 255218 155248 255454
rect 154928 255134 155248 255218
rect 154928 254898 154970 255134
rect 155206 254898 155248 255134
rect 154928 254866 155248 254898
rect 185648 255454 185968 255486
rect 185648 255218 185690 255454
rect 185926 255218 185968 255454
rect 185648 255134 185968 255218
rect 185648 254898 185690 255134
rect 185926 254898 185968 255134
rect 185648 254866 185968 254898
rect 139568 223954 139888 223986
rect 139568 223718 139610 223954
rect 139846 223718 139888 223954
rect 139568 223634 139888 223718
rect 139568 223398 139610 223634
rect 139846 223398 139888 223634
rect 139568 223366 139888 223398
rect 170288 223954 170608 223986
rect 170288 223718 170330 223954
rect 170566 223718 170608 223954
rect 170288 223634 170608 223718
rect 170288 223398 170330 223634
rect 170566 223398 170608 223634
rect 170288 223366 170608 223398
rect 124208 219454 124528 219486
rect 124208 219218 124250 219454
rect 124486 219218 124528 219454
rect 124208 219134 124528 219218
rect 124208 218898 124250 219134
rect 124486 218898 124528 219134
rect 124208 218866 124528 218898
rect 154928 219454 155248 219486
rect 154928 219218 154970 219454
rect 155206 219218 155248 219454
rect 154928 219134 155248 219218
rect 154928 218898 154970 219134
rect 155206 218898 155248 219134
rect 154928 218866 155248 218898
rect 185648 219454 185968 219486
rect 185648 219218 185690 219454
rect 185926 219218 185968 219454
rect 185648 219134 185968 219218
rect 185648 218898 185690 219134
rect 185926 218898 185968 219134
rect 185648 218866 185968 218898
rect 186086 212533 186146 259523
rect 186083 212532 186149 212533
rect 186083 212468 186084 212532
rect 186148 212468 186149 212532
rect 186083 212467 186149 212468
rect 187187 212532 187253 212533
rect 187187 212468 187188 212532
rect 187252 212468 187253 212532
rect 187187 212467 187253 212468
rect 132171 201244 132237 201245
rect 132171 201180 132172 201244
rect 132236 201180 132237 201244
rect 132171 201179 132237 201180
rect 139899 201244 139965 201245
rect 139899 201180 139900 201244
rect 139964 201180 139965 201244
rect 139899 201179 139965 201180
rect 131619 201108 131685 201109
rect 131619 201044 131620 201108
rect 131684 201044 131685 201108
rect 131619 201043 131685 201044
rect 122419 200428 122485 200429
rect 122419 200364 122420 200428
rect 122484 200364 122485 200428
rect 122419 200363 122485 200364
rect 122235 148204 122301 148205
rect 122235 148140 122236 148204
rect 122300 148140 122301 148204
rect 122235 148139 122301 148140
rect 122051 147796 122117 147797
rect 122051 147732 122052 147796
rect 122116 147732 122117 147796
rect 122051 147731 122117 147732
rect 121315 143172 121381 143173
rect 121315 143108 121316 143172
rect 121380 143108 121381 143172
rect 121315 143107 121381 143108
rect 121131 143036 121197 143037
rect 121131 142972 121132 143036
rect 121196 142972 121197 143036
rect 121131 142971 121197 142972
rect 121315 142628 121381 142629
rect 121315 142564 121316 142628
rect 121380 142564 121381 142628
rect 121315 142563 121381 142564
rect 121131 141540 121197 141541
rect 121131 141476 121132 141540
rect 121196 141476 121197 141540
rect 121131 141475 121197 141476
rect 120947 140724 121013 140725
rect 120947 140660 120948 140724
rect 121012 140660 121013 140724
rect 120947 140659 121013 140660
rect 120950 79117 121010 140659
rect 121134 80749 121194 141475
rect 121318 138549 121378 142563
rect 121315 138548 121381 138549
rect 121315 138484 121316 138548
rect 121380 138484 121381 138548
rect 121315 138483 121381 138484
rect 121131 80748 121197 80749
rect 121131 80684 121132 80748
rect 121196 80684 121197 80748
rect 121131 80683 121197 80684
rect 120947 79116 121013 79117
rect 120947 79052 120948 79116
rect 121012 79052 121013 79116
rect 120947 79051 121013 79052
rect 122054 71501 122114 147731
rect 122051 71500 122117 71501
rect 122051 71436 122052 71500
rect 122116 71436 122117 71500
rect 122051 71435 122117 71436
rect 120763 70004 120829 70005
rect 120763 69940 120764 70004
rect 120828 69940 120829 70004
rect 120763 69939 120829 69940
rect 122238 69869 122298 148139
rect 122422 75581 122482 200363
rect 122603 200292 122669 200293
rect 122603 200228 122604 200292
rect 122668 200228 122669 200292
rect 122603 200227 122669 200228
rect 122419 75580 122485 75581
rect 122419 75516 122420 75580
rect 122484 75516 122485 75580
rect 122419 75515 122485 75516
rect 122606 74085 122666 200227
rect 131622 199477 131682 201043
rect 131803 200836 131869 200837
rect 131803 200772 131804 200836
rect 131868 200772 131869 200836
rect 131803 200771 131869 200772
rect 131806 199613 131866 200771
rect 131803 199612 131869 199613
rect 131803 199548 131804 199612
rect 131868 199548 131869 199612
rect 131803 199547 131869 199548
rect 132174 199477 132234 201179
rect 138795 201108 138861 201109
rect 138795 201044 138796 201108
rect 138860 201044 138861 201108
rect 138795 201043 138861 201044
rect 136587 200836 136653 200837
rect 136587 200772 136588 200836
rect 136652 200772 136653 200836
rect 136587 200771 136653 200772
rect 133459 200020 133525 200021
rect 133459 199956 133460 200020
rect 133524 200018 133525 200020
rect 133524 199958 134442 200018
rect 133524 199956 133525 199958
rect 133459 199955 133525 199956
rect 133643 199884 133709 199885
rect 133643 199820 133644 199884
rect 133708 199820 133709 199884
rect 133643 199819 133709 199820
rect 134195 199884 134261 199885
rect 134195 199820 134196 199884
rect 134260 199820 134261 199884
rect 134195 199819 134261 199820
rect 131619 199476 131685 199477
rect 131619 199412 131620 199476
rect 131684 199412 131685 199476
rect 131619 199411 131685 199412
rect 132171 199476 132237 199477
rect 132171 199412 132172 199476
rect 132236 199412 132237 199476
rect 132171 199411 132237 199412
rect 133646 198661 133706 199819
rect 133643 198660 133709 198661
rect 133643 198596 133644 198660
rect 133708 198596 133709 198660
rect 133643 198595 133709 198596
rect 123294 196954 123914 198000
rect 123294 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 123914 196954
rect 123294 196634 123914 196718
rect 123294 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 123914 196634
rect 123294 160954 123914 196398
rect 134011 196348 134077 196349
rect 134011 196284 134012 196348
rect 134076 196284 134077 196348
rect 134011 196283 134077 196284
rect 130331 195804 130397 195805
rect 130331 195740 130332 195804
rect 130396 195740 130397 195804
rect 130331 195739 130397 195740
rect 123294 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 123914 160954
rect 123294 160634 123914 160718
rect 123294 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 123914 160634
rect 122787 146708 122853 146709
rect 122787 146644 122788 146708
rect 122852 146644 122853 146708
rect 122787 146643 122853 146644
rect 122790 138141 122850 146643
rect 123294 142000 123914 160398
rect 124075 151740 124141 151741
rect 124075 151676 124076 151740
rect 124140 151676 124141 151740
rect 124075 151675 124141 151676
rect 124078 141810 124138 151675
rect 130334 142901 130394 195739
rect 134014 191725 134074 196283
rect 134011 191724 134077 191725
rect 134011 191660 134012 191724
rect 134076 191660 134077 191724
rect 134011 191659 134077 191660
rect 134198 191317 134258 199819
rect 134382 198661 134442 199958
rect 135299 199884 135365 199885
rect 135299 199820 135300 199884
rect 135364 199820 135365 199884
rect 135299 199819 135365 199820
rect 136403 199884 136469 199885
rect 136403 199820 136404 199884
rect 136468 199820 136469 199884
rect 136403 199819 136469 199820
rect 134379 198660 134445 198661
rect 134379 198596 134380 198660
rect 134444 198596 134445 198660
rect 134379 198595 134445 198596
rect 135302 196213 135362 199819
rect 136406 199205 136466 199819
rect 136590 199205 136650 200771
rect 138798 199885 138858 201043
rect 139902 199885 139962 201179
rect 151491 200972 151557 200973
rect 151491 200908 151492 200972
rect 151556 200908 151557 200972
rect 151491 200907 151557 200908
rect 140083 200564 140149 200565
rect 140083 200500 140084 200564
rect 140148 200500 140149 200564
rect 140083 200499 140149 200500
rect 140086 200157 140146 200499
rect 140083 200156 140149 200157
rect 140083 200092 140084 200156
rect 140148 200092 140149 200156
rect 140083 200091 140149 200092
rect 151494 199885 151554 200907
rect 153331 200700 153397 200701
rect 153331 200636 153332 200700
rect 153396 200636 153397 200700
rect 153331 200635 153397 200636
rect 151675 200428 151741 200429
rect 151675 200364 151676 200428
rect 151740 200364 151741 200428
rect 151675 200363 151741 200364
rect 137139 199884 137205 199885
rect 137139 199820 137140 199884
rect 137204 199820 137205 199884
rect 137139 199819 137205 199820
rect 137507 199884 137573 199885
rect 137507 199820 137508 199884
rect 137572 199820 137573 199884
rect 137507 199819 137573 199820
rect 138059 199884 138125 199885
rect 138059 199820 138060 199884
rect 138124 199882 138125 199884
rect 138795 199884 138861 199885
rect 138124 199822 138306 199882
rect 138124 199820 138125 199822
rect 138059 199819 138125 199820
rect 137142 199477 137202 199819
rect 137139 199476 137205 199477
rect 137139 199412 137140 199476
rect 137204 199412 137205 199476
rect 137139 199411 137205 199412
rect 135483 199204 135549 199205
rect 135483 199140 135484 199204
rect 135548 199140 135549 199204
rect 135483 199139 135549 199140
rect 136403 199204 136469 199205
rect 136403 199140 136404 199204
rect 136468 199140 136469 199204
rect 136403 199139 136469 199140
rect 136587 199204 136653 199205
rect 136587 199140 136588 199204
rect 136652 199140 136653 199204
rect 136587 199139 136653 199140
rect 135299 196212 135365 196213
rect 135299 196148 135300 196212
rect 135364 196148 135365 196212
rect 135299 196147 135365 196148
rect 135299 196076 135365 196077
rect 135299 196012 135300 196076
rect 135364 196012 135365 196076
rect 135299 196011 135365 196012
rect 134195 191316 134261 191317
rect 134195 191252 134196 191316
rect 134260 191252 134261 191316
rect 134195 191251 134261 191252
rect 135302 149701 135362 196011
rect 135486 191453 135546 199139
rect 136587 197300 136653 197301
rect 136587 197236 136588 197300
rect 136652 197236 136653 197300
rect 136587 197235 136653 197236
rect 135667 195940 135733 195941
rect 135667 195876 135668 195940
rect 135732 195876 135733 195940
rect 135667 195875 135733 195876
rect 135483 191452 135549 191453
rect 135483 191388 135484 191452
rect 135548 191388 135549 191452
rect 135483 191387 135549 191388
rect 135670 191045 135730 195875
rect 135667 191044 135733 191045
rect 135667 190980 135668 191044
rect 135732 190980 135733 191044
rect 135667 190979 135733 190980
rect 136590 151061 136650 197235
rect 136955 197164 137021 197165
rect 136955 197100 136956 197164
rect 137020 197100 137021 197164
rect 136955 197099 137021 197100
rect 136771 196892 136837 196893
rect 136771 196828 136772 196892
rect 136836 196828 136837 196892
rect 136771 196827 136837 196828
rect 136774 151333 136834 196827
rect 136958 189821 137018 197099
rect 137510 196893 137570 199819
rect 137507 196892 137573 196893
rect 137507 196828 137508 196892
rect 137572 196828 137573 196892
rect 137507 196827 137573 196828
rect 138059 196892 138125 196893
rect 138059 196828 138060 196892
rect 138124 196828 138125 196892
rect 138059 196827 138125 196828
rect 136955 189820 137021 189821
rect 136955 189756 136956 189820
rect 137020 189756 137021 189820
rect 136955 189755 137021 189756
rect 136771 151332 136837 151333
rect 136771 151268 136772 151332
rect 136836 151268 136837 151332
rect 136771 151267 136837 151268
rect 138062 151197 138122 196827
rect 138246 189685 138306 199822
rect 138795 199820 138796 199884
rect 138860 199820 138861 199884
rect 138795 199819 138861 199820
rect 139531 199884 139597 199885
rect 139531 199820 139532 199884
rect 139596 199820 139597 199884
rect 139531 199819 139597 199820
rect 139899 199884 139965 199885
rect 139899 199820 139900 199884
rect 139964 199820 139965 199884
rect 139899 199819 139965 199820
rect 141003 199884 141069 199885
rect 141003 199820 141004 199884
rect 141068 199820 141069 199884
rect 141003 199819 141069 199820
rect 142291 199884 142357 199885
rect 142291 199820 142292 199884
rect 142356 199820 142357 199884
rect 142291 199819 142357 199820
rect 143027 199884 143093 199885
rect 143027 199820 143028 199884
rect 143092 199820 143093 199884
rect 143027 199819 143093 199820
rect 146707 199884 146773 199885
rect 146707 199820 146708 199884
rect 146772 199820 146773 199884
rect 146707 199819 146773 199820
rect 147259 199884 147325 199885
rect 147259 199820 147260 199884
rect 147324 199820 147325 199884
rect 147259 199819 147325 199820
rect 148179 199884 148245 199885
rect 148179 199820 148180 199884
rect 148244 199820 148245 199884
rect 148179 199819 148245 199820
rect 151491 199884 151557 199885
rect 151491 199820 151492 199884
rect 151556 199820 151557 199884
rect 151491 199819 151557 199820
rect 139534 198750 139594 199819
rect 139350 198690 139594 198750
rect 138427 198524 138493 198525
rect 138427 198460 138428 198524
rect 138492 198460 138493 198524
rect 138427 198459 138493 198460
rect 138430 190093 138490 198459
rect 138427 190092 138493 190093
rect 138427 190028 138428 190092
rect 138492 190028 138493 190092
rect 138427 190027 138493 190028
rect 138243 189684 138309 189685
rect 138243 189620 138244 189684
rect 138308 189620 138309 189684
rect 138243 189619 138309 189620
rect 138059 151196 138125 151197
rect 138059 151132 138060 151196
rect 138124 151132 138125 151196
rect 138059 151131 138125 151132
rect 136587 151060 136653 151061
rect 136587 150996 136588 151060
rect 136652 150996 136653 151060
rect 136587 150995 136653 150996
rect 135299 149700 135365 149701
rect 135299 149636 135300 149700
rect 135364 149636 135365 149700
rect 135299 149635 135365 149636
rect 139350 147661 139410 198690
rect 141006 198117 141066 199819
rect 141555 199748 141621 199749
rect 141555 199746 141556 199748
rect 141190 199686 141556 199746
rect 141190 199613 141250 199686
rect 141555 199684 141556 199686
rect 141620 199684 141621 199748
rect 141555 199683 141621 199684
rect 141187 199612 141253 199613
rect 141187 199548 141188 199612
rect 141252 199548 141253 199612
rect 141187 199547 141253 199548
rect 141923 199612 141989 199613
rect 141923 199548 141924 199612
rect 141988 199548 141989 199612
rect 141923 199547 141989 199548
rect 141926 198797 141986 199547
rect 141923 198796 141989 198797
rect 141923 198732 141924 198796
rect 141988 198732 141989 198796
rect 141923 198731 141989 198732
rect 141003 198116 141069 198117
rect 141003 198052 141004 198116
rect 141068 198052 141069 198116
rect 141003 198051 141069 198052
rect 139715 197300 139781 197301
rect 139715 197236 139716 197300
rect 139780 197236 139781 197300
rect 139715 197235 139781 197236
rect 139531 195804 139597 195805
rect 139531 195740 139532 195804
rect 139596 195740 139597 195804
rect 139531 195739 139597 195740
rect 139534 186965 139594 195739
rect 139718 191181 139778 197235
rect 139715 191180 139781 191181
rect 139715 191116 139716 191180
rect 139780 191116 139781 191180
rect 139715 191115 139781 191116
rect 139531 186964 139597 186965
rect 139531 186900 139532 186964
rect 139596 186900 139597 186964
rect 139531 186899 139597 186900
rect 141294 178954 141914 198000
rect 142294 196485 142354 199819
rect 142843 199612 142909 199613
rect 142843 199610 142844 199612
rect 142662 199550 142844 199610
rect 142662 198797 142722 199550
rect 142843 199548 142844 199550
rect 142908 199548 142909 199612
rect 142843 199547 142909 199548
rect 142843 199476 142909 199477
rect 142843 199412 142844 199476
rect 142908 199412 142909 199476
rect 142843 199411 142909 199412
rect 142659 198796 142725 198797
rect 142659 198732 142660 198796
rect 142724 198732 142725 198796
rect 142659 198731 142725 198732
rect 142475 196892 142541 196893
rect 142475 196828 142476 196892
rect 142540 196828 142541 196892
rect 142475 196827 142541 196828
rect 142291 196484 142357 196485
rect 142291 196420 142292 196484
rect 142356 196420 142357 196484
rect 142291 196419 142357 196420
rect 142291 194308 142357 194309
rect 142291 194244 142292 194308
rect 142356 194244 142357 194308
rect 142291 194243 142357 194244
rect 141294 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 141914 178954
rect 141294 178634 141914 178718
rect 141294 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 141914 178634
rect 139347 147660 139413 147661
rect 139347 147596 139348 147660
rect 139412 147596 139413 147660
rect 139347 147595 139413 147596
rect 141294 142954 141914 178398
rect 142294 148069 142354 194243
rect 142291 148068 142357 148069
rect 142291 148004 142292 148068
rect 142356 148004 142357 148068
rect 142291 148003 142357 148004
rect 142478 146981 142538 196827
rect 142846 195941 142906 199411
rect 143030 198797 143090 199819
rect 146523 199612 146589 199613
rect 146523 199548 146524 199612
rect 146588 199548 146589 199612
rect 146523 199547 146589 199548
rect 143027 198796 143093 198797
rect 143027 198732 143028 198796
rect 143092 198732 143093 198796
rect 143027 198731 143093 198732
rect 143579 198252 143645 198253
rect 143579 198188 143580 198252
rect 143644 198188 143645 198252
rect 143579 198187 143645 198188
rect 142843 195940 142909 195941
rect 142843 195876 142844 195940
rect 142908 195876 142909 195940
rect 142843 195875 142909 195876
rect 143582 147117 143642 198187
rect 145794 183454 146414 198000
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 143579 147116 143645 147117
rect 143579 147052 143580 147116
rect 143644 147052 143645 147116
rect 143579 147051 143645 147052
rect 142475 146980 142541 146981
rect 142475 146916 142476 146980
rect 142540 146916 142541 146980
rect 142475 146915 142541 146916
rect 130331 142900 130397 142901
rect 130331 142836 130332 142900
rect 130396 142836 130397 142900
rect 130331 142835 130397 142836
rect 141294 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 141914 142954
rect 141294 142634 141914 142718
rect 141294 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 141914 142634
rect 141294 142000 141914 142398
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 142000 146414 146898
rect 123894 141750 124138 141810
rect 122971 139364 123037 139365
rect 122971 139300 122972 139364
rect 123036 139300 123037 139364
rect 122971 139299 123037 139300
rect 122787 138140 122853 138141
rect 122787 138076 122788 138140
rect 122852 138076 122853 138140
rect 122787 138075 122853 138076
rect 122787 132564 122853 132565
rect 122787 132500 122788 132564
rect 122852 132500 122853 132564
rect 122787 132499 122853 132500
rect 122790 132429 122850 132499
rect 122787 132428 122853 132429
rect 122787 132364 122788 132428
rect 122852 132364 122853 132428
rect 122787 132363 122853 132364
rect 122787 122908 122853 122909
rect 122787 122844 122788 122908
rect 122852 122844 122853 122908
rect 122787 122843 122853 122844
rect 122790 122773 122850 122843
rect 122787 122772 122853 122773
rect 122787 122708 122788 122772
rect 122852 122708 122853 122772
rect 122787 122707 122853 122708
rect 122787 113252 122853 113253
rect 122787 113188 122788 113252
rect 122852 113188 122853 113252
rect 122787 113187 122853 113188
rect 122790 113117 122850 113187
rect 122787 113116 122853 113117
rect 122787 113052 122788 113116
rect 122852 113052 122853 113116
rect 122787 113051 122853 113052
rect 122787 103596 122853 103597
rect 122787 103532 122788 103596
rect 122852 103532 122853 103596
rect 122787 103531 122853 103532
rect 122790 103461 122850 103531
rect 122787 103460 122853 103461
rect 122787 103396 122788 103460
rect 122852 103396 122853 103460
rect 122787 103395 122853 103396
rect 122787 93940 122853 93941
rect 122787 93876 122788 93940
rect 122852 93876 122853 93940
rect 122787 93875 122853 93876
rect 122790 92445 122850 93875
rect 122787 92444 122853 92445
rect 122787 92380 122788 92444
rect 122852 92380 122853 92444
rect 122787 92379 122853 92380
rect 122974 78301 123034 139299
rect 123894 138005 123954 141750
rect 129043 140452 129109 140453
rect 129043 140388 129044 140452
rect 129108 140388 129109 140452
rect 129043 140387 129109 140388
rect 124811 140316 124877 140317
rect 124811 140252 124812 140316
rect 124876 140252 124877 140316
rect 124811 140251 124877 140252
rect 126835 140316 126901 140317
rect 126835 140252 126836 140316
rect 126900 140252 126901 140316
rect 126835 140251 126901 140252
rect 124443 139636 124509 139637
rect 124443 139572 124444 139636
rect 124508 139572 124509 139636
rect 124443 139571 124509 139572
rect 124075 139364 124141 139365
rect 124075 139300 124076 139364
rect 124140 139300 124141 139364
rect 124075 139299 124141 139300
rect 124259 139364 124325 139365
rect 124259 139300 124260 139364
rect 124324 139300 124325 139364
rect 124259 139299 124325 139300
rect 123891 138004 123957 138005
rect 123891 137940 123892 138004
rect 123956 137940 123957 138004
rect 123891 137939 123957 137940
rect 122971 78300 123037 78301
rect 122971 78236 122972 78300
rect 123036 78236 123037 78300
rect 122971 78235 123037 78236
rect 122787 74628 122853 74629
rect 122787 74564 122788 74628
rect 122852 74564 122853 74628
rect 122787 74563 122853 74564
rect 122790 74490 122850 74563
rect 122790 74430 123034 74490
rect 122603 74084 122669 74085
rect 122603 74020 122604 74084
rect 122668 74020 122669 74084
rect 122603 74019 122669 74020
rect 122974 73810 123034 74430
rect 122606 73750 123034 73810
rect 122606 71229 122666 73750
rect 122603 71228 122669 71229
rect 122603 71164 122604 71228
rect 122668 71164 122669 71228
rect 122603 71163 122669 71164
rect 122235 69868 122301 69869
rect 122235 69804 122236 69868
rect 122300 69804 122301 69868
rect 122235 69803 122301 69804
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 116531 44300 116597 44301
rect 116531 44236 116532 44300
rect 116596 44236 116597 44300
rect 116531 44235 116597 44236
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 111011 10300 111077 10301
rect 111011 10236 111012 10300
rect 111076 10236 111077 10300
rect 111011 10235 111077 10236
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 114294 7954 114914 43398
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1306 114914 7398
rect 114294 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 114914 -1306
rect 114294 -1626 114914 -1542
rect 114294 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 114914 -1626
rect 114294 -7654 114914 -1862
rect 118794 12454 119414 47898
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2266 119414 11898
rect 118794 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 119414 -2266
rect 118794 -2586 119414 -2502
rect 118794 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 119414 -2586
rect 118794 -7654 119414 -2822
rect 123294 52954 123914 78000
rect 124078 66197 124138 139299
rect 124262 138957 124322 139299
rect 124446 139093 124506 139571
rect 124443 139092 124509 139093
rect 124443 139028 124444 139092
rect 124508 139028 124509 139092
rect 124443 139027 124509 139028
rect 124259 138956 124325 138957
rect 124259 138892 124260 138956
rect 124324 138892 124325 138956
rect 124259 138891 124325 138892
rect 124814 138413 124874 140251
rect 125363 139636 125429 139637
rect 125363 139572 125364 139636
rect 125428 139572 125429 139636
rect 125363 139571 125429 139572
rect 125366 138821 125426 139571
rect 125363 138820 125429 138821
rect 125363 138756 125364 138820
rect 125428 138756 125429 138820
rect 125363 138755 125429 138756
rect 124811 138412 124877 138413
rect 124811 138348 124812 138412
rect 124876 138348 124877 138412
rect 124811 138347 124877 138348
rect 126838 137869 126898 140251
rect 127387 139636 127453 139637
rect 127387 139572 127388 139636
rect 127452 139572 127453 139636
rect 127387 139571 127453 139572
rect 127390 138277 127450 139571
rect 129046 138685 129106 140387
rect 146526 140181 146586 199547
rect 146710 196893 146770 199819
rect 146707 196892 146773 196893
rect 146707 196828 146708 196892
rect 146772 196828 146773 196892
rect 146707 196827 146773 196828
rect 147075 196892 147141 196893
rect 147075 196828 147076 196892
rect 147140 196828 147141 196892
rect 147075 196827 147141 196828
rect 146891 195668 146957 195669
rect 146891 195604 146892 195668
rect 146956 195604 146957 195668
rect 146891 195603 146957 195604
rect 146523 140180 146589 140181
rect 146523 140116 146524 140180
rect 146588 140116 146589 140180
rect 146523 140115 146589 140116
rect 146894 140045 146954 195603
rect 147078 146029 147138 196827
rect 147262 194445 147322 199819
rect 148182 198117 148242 199819
rect 151678 199749 151738 200363
rect 152963 199884 153029 199885
rect 152963 199820 152964 199884
rect 153028 199820 153029 199884
rect 152963 199819 153029 199820
rect 153147 199884 153213 199885
rect 153147 199820 153148 199884
rect 153212 199820 153213 199884
rect 153147 199819 153213 199820
rect 151675 199748 151741 199749
rect 151675 199684 151676 199748
rect 151740 199684 151741 199748
rect 151675 199683 151741 199684
rect 148915 198252 148981 198253
rect 148915 198188 148916 198252
rect 148980 198188 148981 198252
rect 148915 198187 148981 198188
rect 148179 198116 148245 198117
rect 148179 198052 148180 198116
rect 148244 198052 148245 198116
rect 148179 198051 148245 198052
rect 148179 196620 148245 196621
rect 148179 196556 148180 196620
rect 148244 196556 148245 196620
rect 148179 196555 148245 196556
rect 147259 194444 147325 194445
rect 147259 194380 147260 194444
rect 147324 194380 147325 194444
rect 147259 194379 147325 194380
rect 147075 146028 147141 146029
rect 147075 145964 147076 146028
rect 147140 145964 147141 146028
rect 147075 145963 147141 145964
rect 148182 144261 148242 196555
rect 148918 152421 148978 198187
rect 150294 187954 150914 198000
rect 150294 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 150914 187954
rect 150294 187634 150914 187718
rect 150294 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 150914 187634
rect 148915 152420 148981 152421
rect 148915 152356 148916 152420
rect 148980 152356 148981 152420
rect 148915 152355 148981 152356
rect 150294 151954 150914 187398
rect 152966 186965 153026 199819
rect 153150 197981 153210 199819
rect 153334 199613 153394 200635
rect 168419 200292 168485 200293
rect 168419 200228 168420 200292
rect 168484 200228 168485 200292
rect 168419 200227 168485 200228
rect 154803 200156 154869 200157
rect 154803 200092 154804 200156
rect 154868 200092 154869 200156
rect 154803 200091 154869 200092
rect 166395 200156 166461 200157
rect 166395 200092 166396 200156
rect 166460 200092 166461 200156
rect 166395 200091 166461 200092
rect 153515 199884 153581 199885
rect 153515 199820 153516 199884
rect 153580 199820 153581 199884
rect 153515 199819 153581 199820
rect 153883 199884 153949 199885
rect 153883 199820 153884 199884
rect 153948 199820 153949 199884
rect 153883 199819 153949 199820
rect 153331 199612 153397 199613
rect 153331 199548 153332 199612
rect 153396 199548 153397 199612
rect 153331 199547 153397 199548
rect 153518 198117 153578 199819
rect 153515 198116 153581 198117
rect 153515 198052 153516 198116
rect 153580 198052 153581 198116
rect 153515 198051 153581 198052
rect 153147 197980 153213 197981
rect 153147 197916 153148 197980
rect 153212 197916 153213 197980
rect 153147 197915 153213 197916
rect 153886 195669 153946 199819
rect 154806 199610 154866 200091
rect 155171 199884 155237 199885
rect 155171 199820 155172 199884
rect 155236 199820 155237 199884
rect 155171 199819 155237 199820
rect 156643 199884 156709 199885
rect 156643 199820 156644 199884
rect 156708 199820 156709 199884
rect 156643 199819 156709 199820
rect 157747 199884 157813 199885
rect 157747 199820 157748 199884
rect 157812 199820 157813 199884
rect 157747 199819 157813 199820
rect 160139 199884 160205 199885
rect 160139 199820 160140 199884
rect 160204 199820 160205 199884
rect 160139 199819 160205 199820
rect 161059 199884 161125 199885
rect 161059 199820 161060 199884
rect 161124 199820 161125 199884
rect 161059 199819 161125 199820
rect 161795 199884 161861 199885
rect 161795 199820 161796 199884
rect 161860 199820 161861 199884
rect 161795 199819 161861 199820
rect 163083 199884 163149 199885
rect 163083 199820 163084 199884
rect 163148 199820 163149 199884
rect 163083 199819 163149 199820
rect 163819 199884 163885 199885
rect 163819 199820 163820 199884
rect 163884 199820 163885 199884
rect 163819 199819 163885 199820
rect 164923 199884 164989 199885
rect 164923 199820 164924 199884
rect 164988 199820 164989 199884
rect 164923 199819 164989 199820
rect 165843 199884 165909 199885
rect 165843 199820 165844 199884
rect 165908 199820 165909 199884
rect 165843 199819 165909 199820
rect 166027 199884 166093 199885
rect 166027 199820 166028 199884
rect 166092 199820 166093 199884
rect 166027 199819 166093 199820
rect 154622 199550 154866 199610
rect 154622 199477 154682 199550
rect 154619 199476 154685 199477
rect 154619 199412 154620 199476
rect 154684 199412 154685 199476
rect 154619 199411 154685 199412
rect 155174 198525 155234 199819
rect 155171 198524 155237 198525
rect 155171 198460 155172 198524
rect 155236 198460 155237 198524
rect 155171 198459 155237 198460
rect 154435 197980 154501 197981
rect 154435 197916 154436 197980
rect 154500 197916 154501 197980
rect 154435 197915 154501 197916
rect 153883 195668 153949 195669
rect 153883 195604 153884 195668
rect 153948 195604 153949 195668
rect 153883 195603 153949 195604
rect 152963 186964 153029 186965
rect 152963 186900 152964 186964
rect 153028 186900 153029 186964
rect 152963 186899 153029 186900
rect 150294 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 150914 151954
rect 150294 151634 150914 151718
rect 150294 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 150914 151634
rect 148179 144260 148245 144261
rect 148179 144196 148180 144260
rect 148244 144196 148245 144260
rect 148179 144195 148245 144196
rect 150294 142000 150914 151398
rect 154438 151197 154498 197915
rect 154794 192454 155414 198000
rect 156646 193230 156706 199819
rect 157195 199748 157261 199749
rect 157195 199684 157196 199748
rect 157260 199684 157261 199748
rect 157195 199683 157261 199684
rect 157563 199748 157629 199749
rect 157563 199684 157564 199748
rect 157628 199684 157629 199748
rect 157563 199683 157629 199684
rect 157198 196893 157258 199683
rect 157195 196892 157261 196893
rect 157195 196828 157196 196892
rect 157260 196828 157261 196892
rect 157195 196827 157261 196828
rect 157195 196756 157261 196757
rect 157195 196692 157196 196756
rect 157260 196692 157261 196756
rect 157195 196691 157261 196692
rect 156646 193170 157074 193230
rect 154794 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 155414 192454
rect 154794 192134 155414 192218
rect 154794 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 155414 192134
rect 154794 156454 155414 191898
rect 157014 187101 157074 193170
rect 157011 187100 157077 187101
rect 157011 187036 157012 187100
rect 157076 187036 157077 187100
rect 157011 187035 157077 187036
rect 154794 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 155414 156454
rect 154794 156134 155414 156218
rect 154794 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 155414 156134
rect 154435 151196 154501 151197
rect 154435 151132 154436 151196
rect 154500 151132 154501 151196
rect 154435 151131 154501 151132
rect 154794 142000 155414 155898
rect 157198 146981 157258 196691
rect 157566 196621 157626 199683
rect 157750 197845 157810 199819
rect 157747 197844 157813 197845
rect 157747 197780 157748 197844
rect 157812 197780 157813 197844
rect 157747 197779 157813 197780
rect 159294 196954 159914 198000
rect 159294 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 159914 196954
rect 159294 196634 159914 196718
rect 157563 196620 157629 196621
rect 157563 196556 157564 196620
rect 157628 196556 157629 196620
rect 157563 196555 157629 196556
rect 159294 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 159914 196634
rect 158115 196076 158181 196077
rect 158115 196012 158116 196076
rect 158180 196012 158181 196076
rect 158115 196011 158181 196012
rect 158118 189685 158178 196011
rect 158115 189684 158181 189685
rect 158115 189620 158116 189684
rect 158180 189620 158181 189684
rect 158115 189619 158181 189620
rect 159294 160954 159914 196398
rect 160142 195397 160202 199819
rect 161062 196485 161122 199819
rect 161243 199748 161309 199749
rect 161243 199684 161244 199748
rect 161308 199684 161309 199748
rect 161243 199683 161309 199684
rect 161427 199748 161493 199749
rect 161427 199684 161428 199748
rect 161492 199684 161493 199748
rect 161427 199683 161493 199684
rect 161246 199477 161306 199683
rect 161243 199476 161309 199477
rect 161243 199412 161244 199476
rect 161308 199412 161309 199476
rect 161243 199411 161309 199412
rect 161243 198388 161309 198389
rect 161243 198324 161244 198388
rect 161308 198324 161309 198388
rect 161243 198323 161309 198324
rect 161059 196484 161125 196485
rect 161059 196420 161060 196484
rect 161124 196420 161125 196484
rect 161059 196419 161125 196420
rect 160139 195396 160205 195397
rect 160139 195332 160140 195396
rect 160204 195332 160205 195396
rect 160139 195331 160205 195332
rect 159294 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 159914 160954
rect 159294 160634 159914 160718
rect 159294 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 159914 160634
rect 157195 146980 157261 146981
rect 157195 146916 157196 146980
rect 157260 146916 157261 146980
rect 157195 146915 157261 146916
rect 159294 142000 159914 160398
rect 161246 155277 161306 198323
rect 161430 196077 161490 199683
rect 161427 196076 161493 196077
rect 161427 196012 161428 196076
rect 161492 196012 161493 196076
rect 161427 196011 161493 196012
rect 161798 195805 161858 199819
rect 162531 199612 162597 199613
rect 162531 199548 162532 199612
rect 162596 199548 162597 199612
rect 162531 199547 162597 199548
rect 162347 197300 162413 197301
rect 162347 197236 162348 197300
rect 162412 197236 162413 197300
rect 162347 197235 162413 197236
rect 161795 195804 161861 195805
rect 161795 195740 161796 195804
rect 161860 195740 161861 195804
rect 161795 195739 161861 195740
rect 161243 155276 161309 155277
rect 161243 155212 161244 155276
rect 161308 155212 161309 155276
rect 161243 155211 161309 155212
rect 162350 151061 162410 197235
rect 162534 196893 162594 199547
rect 162531 196892 162597 196893
rect 162531 196828 162532 196892
rect 162596 196828 162597 196892
rect 162531 196827 162597 196828
rect 163086 196485 163146 199819
rect 163451 199748 163517 199749
rect 163451 199684 163452 199748
rect 163516 199684 163517 199748
rect 163451 199683 163517 199684
rect 163635 199748 163701 199749
rect 163635 199684 163636 199748
rect 163700 199684 163701 199748
rect 163635 199683 163701 199684
rect 163267 199612 163333 199613
rect 163267 199548 163268 199612
rect 163332 199548 163333 199612
rect 163267 199547 163333 199548
rect 163270 198797 163330 199547
rect 163267 198796 163333 198797
rect 163267 198732 163268 198796
rect 163332 198732 163333 198796
rect 163267 198731 163333 198732
rect 163454 196893 163514 199683
rect 163638 199477 163698 199683
rect 163635 199476 163701 199477
rect 163635 199412 163636 199476
rect 163700 199412 163701 199476
rect 163635 199411 163701 199412
rect 163451 196892 163517 196893
rect 163451 196828 163452 196892
rect 163516 196828 163517 196892
rect 163451 196827 163517 196828
rect 163083 196484 163149 196485
rect 163083 196420 163084 196484
rect 163148 196420 163149 196484
rect 163083 196419 163149 196420
rect 163822 196349 163882 199819
rect 164739 199748 164805 199749
rect 164739 199684 164740 199748
rect 164804 199684 164805 199748
rect 164739 199683 164805 199684
rect 164742 197437 164802 199683
rect 164926 197573 164986 199819
rect 165291 199748 165357 199749
rect 165291 199684 165292 199748
rect 165356 199684 165357 199748
rect 165291 199683 165357 199684
rect 165294 197981 165354 199683
rect 165291 197980 165357 197981
rect 165291 197916 165292 197980
rect 165356 197916 165357 197980
rect 165291 197915 165357 197916
rect 164923 197572 164989 197573
rect 164923 197508 164924 197572
rect 164988 197508 164989 197572
rect 164923 197507 164989 197508
rect 164739 197436 164805 197437
rect 164739 197372 164740 197436
rect 164804 197372 164805 197436
rect 164739 197371 164805 197372
rect 164923 196484 164989 196485
rect 164923 196420 164924 196484
rect 164988 196420 164989 196484
rect 164923 196419 164989 196420
rect 163819 196348 163885 196349
rect 163819 196284 163820 196348
rect 163884 196284 163885 196348
rect 163819 196283 163885 196284
rect 164926 191045 164986 196419
rect 165846 196077 165906 199819
rect 166030 196349 166090 199819
rect 166398 199477 166458 200091
rect 166579 199884 166645 199885
rect 166579 199820 166580 199884
rect 166644 199820 166645 199884
rect 166579 199819 166645 199820
rect 167499 199884 167565 199885
rect 167499 199820 167500 199884
rect 167564 199820 167565 199884
rect 167499 199819 167565 199820
rect 167683 199884 167749 199885
rect 167683 199820 167684 199884
rect 167748 199820 167749 199884
rect 167683 199819 167749 199820
rect 166395 199476 166461 199477
rect 166395 199412 166396 199476
rect 166460 199412 166461 199476
rect 166395 199411 166461 199412
rect 166027 196348 166093 196349
rect 166027 196284 166028 196348
rect 166092 196284 166093 196348
rect 166027 196283 166093 196284
rect 165843 196076 165909 196077
rect 165843 196012 165844 196076
rect 165908 196012 165909 196076
rect 165843 196011 165909 196012
rect 166582 195805 166642 199819
rect 167502 196213 167562 199819
rect 167686 196485 167746 199819
rect 168422 199613 168482 200227
rect 168974 200094 169770 200154
rect 168603 199884 168669 199885
rect 168603 199820 168604 199884
rect 168668 199820 168669 199884
rect 168603 199819 168669 199820
rect 168787 199884 168853 199885
rect 168787 199820 168788 199884
rect 168852 199820 168853 199884
rect 168787 199819 168853 199820
rect 168419 199612 168485 199613
rect 168419 199548 168420 199612
rect 168484 199548 168485 199612
rect 168419 199547 168485 199548
rect 168606 198389 168666 199819
rect 168603 198388 168669 198389
rect 168603 198324 168604 198388
rect 168668 198324 168669 198388
rect 168603 198323 168669 198324
rect 167683 196484 167749 196485
rect 167683 196420 167684 196484
rect 167748 196420 167749 196484
rect 167683 196419 167749 196420
rect 168790 196349 168850 199819
rect 168974 199341 169034 200094
rect 169523 200020 169589 200021
rect 169523 199956 169524 200020
rect 169588 199956 169589 200020
rect 169523 199955 169589 199956
rect 169155 199612 169221 199613
rect 169155 199548 169156 199612
rect 169220 199548 169221 199612
rect 169155 199547 169221 199548
rect 168971 199340 169037 199341
rect 168971 199276 168972 199340
rect 169036 199276 169037 199340
rect 168971 199275 169037 199276
rect 169158 198661 169218 199547
rect 169339 199476 169405 199477
rect 169339 199412 169340 199476
rect 169404 199412 169405 199476
rect 169339 199411 169405 199412
rect 169155 198660 169221 198661
rect 169155 198596 169156 198660
rect 169220 198596 169221 198660
rect 169155 198595 169221 198596
rect 169155 196484 169221 196485
rect 169155 196420 169156 196484
rect 169220 196420 169221 196484
rect 169155 196419 169221 196420
rect 168787 196348 168853 196349
rect 168787 196284 168788 196348
rect 168852 196284 168853 196348
rect 168787 196283 168853 196284
rect 167499 196212 167565 196213
rect 167499 196148 167500 196212
rect 167564 196148 167565 196212
rect 167499 196147 167565 196148
rect 166579 195804 166645 195805
rect 166579 195740 166580 195804
rect 166644 195740 166645 195804
rect 166579 195739 166645 195740
rect 164923 191044 164989 191045
rect 164923 190980 164924 191044
rect 164988 190980 164989 191044
rect 164923 190979 164989 190980
rect 169158 155685 169218 196419
rect 169155 155684 169221 155685
rect 169155 155620 169156 155684
rect 169220 155620 169221 155684
rect 169155 155619 169221 155620
rect 169342 155549 169402 199411
rect 169526 196213 169586 199955
rect 169710 199477 169770 200094
rect 170811 200020 170877 200021
rect 170811 199956 170812 200020
rect 170876 199956 170877 200020
rect 172835 200020 172901 200021
rect 172835 200018 172836 200020
rect 170811 199955 170877 199956
rect 172470 199958 172836 200018
rect 169891 199884 169957 199885
rect 169891 199820 169892 199884
rect 169956 199820 169957 199884
rect 169891 199819 169957 199820
rect 170627 199884 170693 199885
rect 170627 199820 170628 199884
rect 170692 199820 170693 199884
rect 170627 199819 170693 199820
rect 169707 199476 169773 199477
rect 169707 199412 169708 199476
rect 169772 199412 169773 199476
rect 169707 199411 169773 199412
rect 169523 196212 169589 196213
rect 169523 196148 169524 196212
rect 169588 196148 169589 196212
rect 169523 196147 169589 196148
rect 169894 196077 169954 199819
rect 170075 199748 170141 199749
rect 170075 199684 170076 199748
rect 170140 199684 170141 199748
rect 170075 199683 170141 199684
rect 170078 196349 170138 199683
rect 170075 196348 170141 196349
rect 170075 196284 170076 196348
rect 170140 196284 170141 196348
rect 170075 196283 170141 196284
rect 170630 196213 170690 199819
rect 170814 196485 170874 199955
rect 172470 199885 172530 199958
rect 172835 199956 172836 199958
rect 172900 199956 172901 200020
rect 172835 199955 172901 199956
rect 174123 200020 174189 200021
rect 174123 199956 174124 200020
rect 174188 199956 174189 200020
rect 174123 199955 174189 199956
rect 171363 199884 171429 199885
rect 171363 199820 171364 199884
rect 171428 199820 171429 199884
rect 171363 199819 171429 199820
rect 171547 199884 171613 199885
rect 171547 199820 171548 199884
rect 171612 199820 171613 199884
rect 171547 199819 171613 199820
rect 172467 199884 172533 199885
rect 172467 199820 172468 199884
rect 172532 199820 172533 199884
rect 172467 199819 172533 199820
rect 172651 199884 172717 199885
rect 172651 199820 172652 199884
rect 172716 199820 172717 199884
rect 172651 199819 172717 199820
rect 173387 199884 173453 199885
rect 173387 199820 173388 199884
rect 173452 199820 173453 199884
rect 173387 199819 173453 199820
rect 171366 196485 171426 199819
rect 171550 198661 171610 199819
rect 171731 199748 171797 199749
rect 171731 199684 171732 199748
rect 171796 199684 171797 199748
rect 171731 199683 171797 199684
rect 171915 199748 171981 199749
rect 171915 199684 171916 199748
rect 171980 199684 171981 199748
rect 171915 199683 171981 199684
rect 172467 199748 172533 199749
rect 172467 199684 172468 199748
rect 172532 199684 172533 199748
rect 172467 199683 172533 199684
rect 171734 199477 171794 199683
rect 171731 199476 171797 199477
rect 171731 199412 171732 199476
rect 171796 199412 171797 199476
rect 171731 199411 171797 199412
rect 171547 198660 171613 198661
rect 171547 198596 171548 198660
rect 171612 198596 171613 198660
rect 171547 198595 171613 198596
rect 170811 196484 170877 196485
rect 170811 196420 170812 196484
rect 170876 196420 170877 196484
rect 170811 196419 170877 196420
rect 171363 196484 171429 196485
rect 171363 196420 171364 196484
rect 171428 196420 171429 196484
rect 171363 196419 171429 196420
rect 171918 196213 171978 199683
rect 172283 197980 172349 197981
rect 172283 197916 172284 197980
rect 172348 197916 172349 197980
rect 172283 197915 172349 197916
rect 170627 196212 170693 196213
rect 170627 196148 170628 196212
rect 170692 196148 170693 196212
rect 170627 196147 170693 196148
rect 171915 196212 171981 196213
rect 171915 196148 171916 196212
rect 171980 196148 171981 196212
rect 171915 196147 171981 196148
rect 169891 196076 169957 196077
rect 169891 196012 169892 196076
rect 169956 196012 169957 196076
rect 169891 196011 169957 196012
rect 172286 190093 172346 197915
rect 172470 196349 172530 199683
rect 172467 196348 172533 196349
rect 172467 196284 172468 196348
rect 172532 196284 172533 196348
rect 172467 196283 172533 196284
rect 172654 194173 172714 199819
rect 172973 199748 173039 199749
rect 172973 199684 172974 199748
rect 173038 199746 173039 199748
rect 173038 199684 173082 199746
rect 172973 199683 173082 199684
rect 173022 194445 173082 199683
rect 173390 196349 173450 199819
rect 173571 199748 173637 199749
rect 173571 199684 173572 199748
rect 173636 199684 173637 199748
rect 173571 199683 173637 199684
rect 173387 196348 173453 196349
rect 173387 196284 173388 196348
rect 173452 196284 173453 196348
rect 173387 196283 173453 196284
rect 173019 194444 173085 194445
rect 173019 194380 173020 194444
rect 173084 194380 173085 194444
rect 173019 194379 173085 194380
rect 172651 194172 172717 194173
rect 172651 194108 172652 194172
rect 172716 194108 172717 194172
rect 172651 194107 172717 194108
rect 173574 194037 173634 199683
rect 174126 198933 174186 199955
rect 174859 199884 174925 199885
rect 174859 199820 174860 199884
rect 174924 199820 174925 199884
rect 174859 199819 174925 199820
rect 175411 199884 175477 199885
rect 175411 199820 175412 199884
rect 175476 199820 175477 199884
rect 175411 199819 175477 199820
rect 175963 199884 176029 199885
rect 175963 199820 175964 199884
rect 176028 199820 176029 199884
rect 175963 199819 176029 199820
rect 176515 199884 176581 199885
rect 176515 199820 176516 199884
rect 176580 199820 176581 199884
rect 176515 199819 176581 199820
rect 174307 199748 174373 199749
rect 174307 199684 174308 199748
rect 174372 199684 174373 199748
rect 174307 199683 174373 199684
rect 174123 198932 174189 198933
rect 174123 198868 174124 198932
rect 174188 198868 174189 198932
rect 174310 198930 174370 199683
rect 174862 199341 174922 199819
rect 174859 199340 174925 199341
rect 174859 199276 174860 199340
rect 174924 199276 174925 199340
rect 174859 199275 174925 199276
rect 174491 198932 174557 198933
rect 174491 198930 174492 198932
rect 174310 198870 174492 198930
rect 174123 198867 174189 198868
rect 174491 198868 174492 198870
rect 174556 198868 174557 198932
rect 174491 198867 174557 198868
rect 173755 197436 173821 197437
rect 173755 197372 173756 197436
rect 173820 197372 173821 197436
rect 173755 197371 173821 197372
rect 173571 194036 173637 194037
rect 173571 193972 173572 194036
rect 173636 193972 173637 194036
rect 173571 193971 173637 193972
rect 172283 190092 172349 190093
rect 172283 190028 172284 190092
rect 172348 190028 172349 190092
rect 172283 190027 172349 190028
rect 169339 155548 169405 155549
rect 169339 155484 169340 155548
rect 169404 155484 169405 155548
rect 169339 155483 169405 155484
rect 162347 151060 162413 151061
rect 162347 150996 162348 151060
rect 162412 150996 162413 151060
rect 162347 150995 162413 150996
rect 173758 149973 173818 197371
rect 175414 194853 175474 199819
rect 175595 198524 175661 198525
rect 175595 198460 175596 198524
rect 175660 198460 175661 198524
rect 175595 198459 175661 198460
rect 175411 194852 175477 194853
rect 175411 194788 175412 194852
rect 175476 194788 175477 194852
rect 175411 194787 175477 194788
rect 175598 194037 175658 198459
rect 175966 197437 176026 199819
rect 176331 197708 176397 197709
rect 176331 197644 176332 197708
rect 176396 197644 176397 197708
rect 176331 197643 176397 197644
rect 175963 197436 176029 197437
rect 175963 197372 175964 197436
rect 176028 197372 176029 197436
rect 175963 197371 176029 197372
rect 175595 194036 175661 194037
rect 175595 193972 175596 194036
rect 175660 193972 175661 194036
rect 175595 193971 175661 193972
rect 176334 155413 176394 197643
rect 176331 155412 176397 155413
rect 176331 155348 176332 155412
rect 176396 155348 176397 155412
rect 176331 155347 176397 155348
rect 176518 150245 176578 199819
rect 177294 178954 177914 198000
rect 177294 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 177914 178954
rect 177294 178634 177914 178718
rect 177294 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 177914 178634
rect 176515 150244 176581 150245
rect 176515 150180 176516 150244
rect 176580 150180 176581 150244
rect 176515 150179 176581 150180
rect 173755 149972 173821 149973
rect 173755 149908 173756 149972
rect 173820 149908 173821 149972
rect 173755 149907 173821 149908
rect 177294 142954 177914 178398
rect 177294 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 177914 142954
rect 177294 142634 177914 142718
rect 177294 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 177914 142634
rect 177294 142000 177914 142398
rect 181794 183454 182414 198000
rect 184059 195940 184125 195941
rect 184059 195876 184060 195940
rect 184124 195876 184125 195940
rect 184059 195875 184125 195876
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 142000 182414 146898
rect 146891 140044 146957 140045
rect 146891 139980 146892 140044
rect 146956 139980 146957 140044
rect 146891 139979 146957 139980
rect 129043 138684 129109 138685
rect 129043 138620 129044 138684
rect 129108 138620 129109 138684
rect 129043 138619 129109 138620
rect 127387 138276 127453 138277
rect 127387 138212 127388 138276
rect 127452 138212 127453 138276
rect 127387 138211 127453 138212
rect 184062 138005 184122 195875
rect 186083 192676 186149 192677
rect 186083 192612 186084 192676
rect 186148 192612 186149 192676
rect 186083 192611 186149 192612
rect 185347 191180 185413 191181
rect 185347 191116 185348 191180
rect 185412 191116 185413 191180
rect 185347 191115 185413 191116
rect 185350 138277 185410 191115
rect 185899 141540 185965 141541
rect 185899 141476 185900 141540
rect 185964 141476 185965 141540
rect 185899 141475 185965 141476
rect 185347 138276 185413 138277
rect 185347 138212 185348 138276
rect 185412 138212 185413 138276
rect 185347 138211 185413 138212
rect 185902 138141 185962 141475
rect 185899 138140 185965 138141
rect 185899 138076 185900 138140
rect 185964 138076 185965 138140
rect 185899 138075 185965 138076
rect 184059 138004 184125 138005
rect 184059 137940 184060 138004
rect 184124 137940 184125 138004
rect 184059 137939 184125 137940
rect 126835 137868 126901 137869
rect 126835 137804 126836 137868
rect 126900 137804 126901 137868
rect 126835 137803 126901 137804
rect 185347 137868 185413 137869
rect 185347 137804 185348 137868
rect 185412 137804 185413 137868
rect 185347 137803 185413 137804
rect 139568 115954 139888 115986
rect 139568 115718 139610 115954
rect 139846 115718 139888 115954
rect 139568 115634 139888 115718
rect 139568 115398 139610 115634
rect 139846 115398 139888 115634
rect 139568 115366 139888 115398
rect 170288 115954 170608 115986
rect 170288 115718 170330 115954
rect 170566 115718 170608 115954
rect 170288 115634 170608 115718
rect 170288 115398 170330 115634
rect 170566 115398 170608 115634
rect 170288 115366 170608 115398
rect 124208 111454 124528 111486
rect 124208 111218 124250 111454
rect 124486 111218 124528 111454
rect 124208 111134 124528 111218
rect 124208 110898 124250 111134
rect 124486 110898 124528 111134
rect 124208 110866 124528 110898
rect 154928 111454 155248 111486
rect 154928 111218 154970 111454
rect 155206 111218 155248 111454
rect 154928 111134 155248 111218
rect 154928 110898 154970 111134
rect 155206 110898 155248 111134
rect 154928 110866 155248 110898
rect 125547 81972 125613 81973
rect 125547 81908 125548 81972
rect 125612 81908 125613 81972
rect 125547 81907 125613 81908
rect 125550 75037 125610 81907
rect 184059 81700 184125 81701
rect 184059 81636 184060 81700
rect 184124 81636 184125 81700
rect 184059 81635 184125 81636
rect 181299 81564 181365 81565
rect 181299 81500 181300 81564
rect 181364 81500 181365 81564
rect 181299 81499 181365 81500
rect 176331 81292 176397 81293
rect 176331 81228 176332 81292
rect 176396 81228 176397 81292
rect 176331 81227 176397 81228
rect 129227 81156 129293 81157
rect 129227 81092 129228 81156
rect 129292 81092 129293 81156
rect 129227 81091 129293 81092
rect 170443 81156 170509 81157
rect 170443 81092 170444 81156
rect 170508 81092 170509 81156
rect 170443 81091 170509 81092
rect 129230 80613 129290 81091
rect 146891 81020 146957 81021
rect 146891 80956 146892 81020
rect 146956 80956 146957 81020
rect 146891 80955 146957 80956
rect 129227 80612 129293 80613
rect 129227 80548 129228 80612
rect 129292 80548 129293 80612
rect 129227 80547 129293 80548
rect 143395 80068 143461 80069
rect 139534 80006 140146 80066
rect 134011 79932 134077 79933
rect 134011 79868 134012 79932
rect 134076 79868 134077 79932
rect 134011 79867 134077 79868
rect 135483 79932 135549 79933
rect 135483 79868 135484 79932
rect 135548 79868 135549 79932
rect 135483 79867 135549 79868
rect 137691 79932 137757 79933
rect 137691 79868 137692 79932
rect 137756 79868 137757 79932
rect 137691 79867 137757 79868
rect 138059 79932 138125 79933
rect 138059 79868 138060 79932
rect 138124 79868 138125 79932
rect 138059 79867 138125 79868
rect 138979 79932 139045 79933
rect 138979 79868 138980 79932
rect 139044 79868 139045 79932
rect 138979 79867 139045 79868
rect 133827 79660 133893 79661
rect 133827 79596 133828 79660
rect 133892 79596 133893 79660
rect 133827 79595 133893 79596
rect 133459 79524 133525 79525
rect 133459 79460 133460 79524
rect 133524 79460 133525 79524
rect 133459 79459 133525 79460
rect 125547 75036 125613 75037
rect 125547 74972 125548 75036
rect 125612 74972 125613 75036
rect 125547 74971 125613 74972
rect 124075 66196 124141 66197
rect 124075 66132 124076 66196
rect 124140 66132 124141 66196
rect 124075 66131 124141 66132
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3226 123914 16398
rect 123294 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 123914 -3226
rect 123294 -3546 123914 -3462
rect 123294 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 123914 -3546
rect 123294 -7654 123914 -3782
rect 127794 57454 128414 78000
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -4186 128414 20898
rect 127794 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 128414 -4186
rect 127794 -4506 128414 -4422
rect 127794 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 128414 -4506
rect 127794 -7654 128414 -4742
rect 132294 61954 132914 78000
rect 133275 77756 133341 77757
rect 133275 77692 133276 77756
rect 133340 77692 133341 77756
rect 133275 77691 133341 77692
rect 133091 76668 133157 76669
rect 133091 76604 133092 76668
rect 133156 76604 133157 76668
rect 133091 76603 133157 76604
rect 132294 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 132914 61954
rect 132294 61634 132914 61718
rect 132294 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 132914 61634
rect 132294 25954 132914 61398
rect 133094 52461 133154 76603
rect 133278 56541 133338 77691
rect 133462 63341 133522 79459
rect 133459 63340 133525 63341
rect 133459 63276 133460 63340
rect 133524 63276 133525 63340
rect 133459 63275 133525 63276
rect 133275 56540 133341 56541
rect 133275 56476 133276 56540
rect 133340 56476 133341 56540
rect 133275 56475 133341 56476
rect 133091 52460 133157 52461
rect 133091 52396 133092 52460
rect 133156 52396 133157 52460
rect 133091 52395 133157 52396
rect 133830 49605 133890 79595
rect 134014 78437 134074 79867
rect 134195 78572 134261 78573
rect 134195 78508 134196 78572
rect 134260 78508 134261 78572
rect 134195 78507 134261 78508
rect 134011 78436 134077 78437
rect 134011 78372 134012 78436
rect 134076 78372 134077 78436
rect 134011 78371 134077 78372
rect 134011 78300 134077 78301
rect 134011 78236 134012 78300
rect 134076 78236 134077 78300
rect 134011 78235 134077 78236
rect 134014 50829 134074 78235
rect 134198 57765 134258 78507
rect 135299 77620 135365 77621
rect 135299 77556 135300 77620
rect 135364 77556 135365 77620
rect 135299 77555 135365 77556
rect 134379 77348 134445 77349
rect 134379 77284 134380 77348
rect 134444 77284 134445 77348
rect 134379 77283 134445 77284
rect 134382 74221 134442 77283
rect 134379 74220 134445 74221
rect 134379 74156 134380 74220
rect 134444 74156 134445 74220
rect 134379 74155 134445 74156
rect 134195 57764 134261 57765
rect 134195 57700 134196 57764
rect 134260 57700 134261 57764
rect 134195 57699 134261 57700
rect 134011 50828 134077 50829
rect 134011 50764 134012 50828
rect 134076 50764 134077 50828
rect 134011 50763 134077 50764
rect 133827 49604 133893 49605
rect 133827 49540 133828 49604
rect 133892 49540 133893 49604
rect 133827 49539 133893 49540
rect 135302 46885 135362 77555
rect 135486 48245 135546 79867
rect 137507 78300 137573 78301
rect 137507 78236 137508 78300
rect 137572 78236 137573 78300
rect 137507 78235 137573 78236
rect 135667 77348 135733 77349
rect 135667 77284 135668 77348
rect 135732 77284 135733 77348
rect 135667 77283 135733 77284
rect 135670 64837 135730 77283
rect 136794 66454 137414 78000
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 135667 64836 135733 64837
rect 135667 64772 135668 64836
rect 135732 64772 135733 64836
rect 135667 64771 135733 64772
rect 135483 48244 135549 48245
rect 135483 48180 135484 48244
rect 135548 48180 135549 48244
rect 135483 48179 135549 48180
rect 135299 46884 135365 46885
rect 135299 46820 135300 46884
rect 135364 46820 135365 46884
rect 135299 46819 135365 46820
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 132294 -5146 132914 25398
rect 132294 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 132914 -5146
rect 132294 -5466 132914 -5382
rect 132294 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 132914 -5466
rect 132294 -7654 132914 -5702
rect 136794 30454 137414 65898
rect 137510 53821 137570 78235
rect 137507 53820 137573 53821
rect 137507 53756 137508 53820
rect 137572 53756 137573 53820
rect 137507 53755 137573 53756
rect 137694 44165 137754 79867
rect 138062 50965 138122 79867
rect 138611 79796 138677 79797
rect 138611 79732 138612 79796
rect 138676 79732 138677 79796
rect 138611 79731 138677 79732
rect 138243 79660 138309 79661
rect 138243 79596 138244 79660
rect 138308 79596 138309 79660
rect 138243 79595 138309 79596
rect 138246 57901 138306 79595
rect 138427 78572 138493 78573
rect 138427 78508 138428 78572
rect 138492 78508 138493 78572
rect 138427 78507 138493 78508
rect 138430 63205 138490 78507
rect 138614 63477 138674 79731
rect 138982 78029 139042 79867
rect 139347 78572 139413 78573
rect 139347 78508 139348 78572
rect 139412 78508 139413 78572
rect 139347 78507 139413 78508
rect 138979 78028 139045 78029
rect 138979 77964 138980 78028
rect 139044 77964 139045 78028
rect 138979 77963 139045 77964
rect 138611 63476 138677 63477
rect 138611 63412 138612 63476
rect 138676 63412 138677 63476
rect 138611 63411 138677 63412
rect 138427 63204 138493 63205
rect 138427 63140 138428 63204
rect 138492 63140 138493 63204
rect 138427 63139 138493 63140
rect 138243 57900 138309 57901
rect 138243 57836 138244 57900
rect 138308 57836 138309 57900
rect 138243 57835 138309 57836
rect 139350 55045 139410 78507
rect 139534 55181 139594 80006
rect 140086 79933 140146 80006
rect 143395 80004 143396 80068
rect 143460 80004 143461 80068
rect 143395 80003 143461 80004
rect 139715 79932 139781 79933
rect 139715 79868 139716 79932
rect 139780 79868 139781 79932
rect 139715 79867 139781 79868
rect 140083 79932 140149 79933
rect 140083 79868 140084 79932
rect 140148 79868 140149 79932
rect 140083 79867 140149 79868
rect 141003 79932 141069 79933
rect 141003 79868 141004 79932
rect 141068 79868 141069 79932
rect 141003 79867 141069 79868
rect 142659 79932 142725 79933
rect 142659 79868 142660 79932
rect 142724 79868 142725 79932
rect 142659 79867 142725 79868
rect 139718 62117 139778 79867
rect 139899 79796 139965 79797
rect 139899 79732 139900 79796
rect 139964 79732 139965 79796
rect 139899 79731 139965 79732
rect 139902 65925 139962 79731
rect 140819 78300 140885 78301
rect 140819 78236 140820 78300
rect 140884 78236 140885 78300
rect 140819 78235 140885 78236
rect 140822 67285 140882 78235
rect 141006 77893 141066 79867
rect 141003 77892 141069 77893
rect 141003 77828 141004 77892
rect 141068 77828 141069 77892
rect 141003 77827 141069 77828
rect 141294 70954 141914 78000
rect 142662 77893 142722 79867
rect 142659 77892 142725 77893
rect 142659 77828 142660 77892
rect 142724 77828 142725 77892
rect 142659 77827 142725 77828
rect 143398 77310 143458 80003
rect 143579 79932 143645 79933
rect 143579 79868 143580 79932
rect 143644 79868 143645 79932
rect 143579 79867 143645 79868
rect 145603 79932 145669 79933
rect 145603 79868 145604 79932
rect 145668 79868 145669 79932
rect 145603 79867 145669 79868
rect 143582 78981 143642 79867
rect 144315 79660 144381 79661
rect 144315 79596 144316 79660
rect 144380 79596 144381 79660
rect 144315 79595 144381 79596
rect 143579 78980 143645 78981
rect 143579 78916 143580 78980
rect 143644 78916 143645 78980
rect 143579 78915 143645 78916
rect 143763 78028 143829 78029
rect 143763 77964 143764 78028
rect 143828 77964 143829 78028
rect 143763 77963 143829 77964
rect 143398 77250 143642 77310
rect 141294 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 141914 70954
rect 141294 70634 141914 70718
rect 141294 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 141914 70634
rect 140819 67284 140885 67285
rect 140819 67220 140820 67284
rect 140884 67220 140885 67284
rect 140819 67219 140885 67220
rect 139899 65924 139965 65925
rect 139899 65860 139900 65924
rect 139964 65860 139965 65924
rect 139899 65859 139965 65860
rect 139715 62116 139781 62117
rect 139715 62052 139716 62116
rect 139780 62052 139781 62116
rect 139715 62051 139781 62052
rect 139531 55180 139597 55181
rect 139531 55116 139532 55180
rect 139596 55116 139597 55180
rect 139531 55115 139597 55116
rect 139347 55044 139413 55045
rect 139347 54980 139348 55044
rect 139412 54980 139413 55044
rect 139347 54979 139413 54980
rect 138059 50964 138125 50965
rect 138059 50900 138060 50964
rect 138124 50900 138125 50964
rect 138059 50899 138125 50900
rect 137691 44164 137757 44165
rect 137691 44100 137692 44164
rect 137756 44100 137757 44164
rect 137691 44099 137757 44100
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 136794 -6106 137414 29898
rect 136794 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 137414 -6106
rect 136794 -6426 137414 -6342
rect 136794 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 137414 -6426
rect 136794 -7654 137414 -6662
rect 141294 34954 141914 70398
rect 143582 64837 143642 77250
rect 143579 64836 143645 64837
rect 143579 64772 143580 64836
rect 143644 64772 143645 64836
rect 143579 64771 143645 64772
rect 143582 64565 143642 64771
rect 143766 64701 143826 77963
rect 143947 77892 144013 77893
rect 143947 77828 143948 77892
rect 144012 77828 144013 77892
rect 143947 77827 144013 77828
rect 143950 70410 144010 77827
rect 143950 70350 144194 70410
rect 144134 68509 144194 70350
rect 144131 68508 144197 68509
rect 144131 68444 144132 68508
rect 144196 68444 144197 68508
rect 144131 68443 144197 68444
rect 143763 64700 143829 64701
rect 143763 64636 143764 64700
rect 143828 64636 143829 64700
rect 143763 64635 143829 64636
rect 143579 64564 143645 64565
rect 143579 64500 143580 64564
rect 143644 64500 143645 64564
rect 143579 64499 143645 64500
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141294 -7066 141914 34398
rect 144134 6221 144194 68443
rect 144318 67557 144378 79595
rect 145419 79524 145485 79525
rect 145419 79460 145420 79524
rect 145484 79460 145485 79524
rect 145419 79459 145485 79460
rect 145422 73133 145482 79459
rect 145606 75445 145666 79867
rect 146523 79796 146589 79797
rect 146523 79732 146524 79796
rect 146588 79732 146589 79796
rect 146523 79731 146589 79732
rect 145794 75454 146414 78000
rect 145603 75444 145669 75445
rect 145603 75380 145604 75444
rect 145668 75380 145669 75444
rect 145603 75379 145669 75380
rect 145419 73132 145485 73133
rect 145419 73068 145420 73132
rect 145484 73068 145485 73132
rect 145419 73067 145485 73068
rect 144315 67556 144381 67557
rect 144315 67492 144316 67556
rect 144380 67492 144381 67556
rect 144315 67491 144381 67492
rect 144315 64836 144381 64837
rect 144315 64772 144316 64836
rect 144380 64772 144381 64836
rect 144315 64771 144381 64772
rect 144318 8941 144378 64771
rect 144499 64700 144565 64701
rect 144499 64636 144500 64700
rect 144564 64636 144565 64700
rect 144499 64635 144565 64636
rect 144502 35189 144562 64635
rect 144499 35188 144565 35189
rect 144499 35124 144500 35188
rect 144564 35124 144565 35188
rect 144499 35123 144565 35124
rect 145422 22677 145482 73067
rect 145606 67693 145666 75379
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145603 67692 145669 67693
rect 145603 67628 145604 67692
rect 145668 67628 145669 67692
rect 145603 67627 145669 67628
rect 145794 39454 146414 74898
rect 146526 72997 146586 79731
rect 146894 79661 146954 80955
rect 149835 80884 149901 80885
rect 149835 80820 149836 80884
rect 149900 80820 149901 80884
rect 149835 80819 149901 80820
rect 149838 79933 149898 80819
rect 151307 80204 151373 80205
rect 151307 80140 151308 80204
rect 151372 80140 151373 80204
rect 151307 80139 151373 80140
rect 147075 79932 147141 79933
rect 147075 79868 147076 79932
rect 147140 79868 147141 79932
rect 147075 79867 147141 79868
rect 147811 79932 147877 79933
rect 147811 79868 147812 79932
rect 147876 79868 147877 79932
rect 147811 79867 147877 79868
rect 148179 79932 148245 79933
rect 148179 79868 148180 79932
rect 148244 79868 148245 79932
rect 148179 79867 148245 79868
rect 149835 79932 149901 79933
rect 149835 79868 149836 79932
rect 149900 79868 149901 79932
rect 149835 79867 149901 79868
rect 146891 79660 146957 79661
rect 146891 79596 146892 79660
rect 146956 79596 146957 79660
rect 146891 79595 146957 79596
rect 146891 77484 146957 77485
rect 146891 77420 146892 77484
rect 146956 77420 146957 77484
rect 146891 77419 146957 77420
rect 146523 72996 146589 72997
rect 146523 72932 146524 72996
rect 146588 72932 146589 72996
rect 146523 72931 146589 72932
rect 146526 68237 146586 72931
rect 146894 71365 146954 77419
rect 147078 72861 147138 79867
rect 147814 79389 147874 79867
rect 148182 79389 148242 79867
rect 147811 79388 147877 79389
rect 147811 79324 147812 79388
rect 147876 79324 147877 79388
rect 147811 79323 147877 79324
rect 148179 79388 148245 79389
rect 148179 79324 148180 79388
rect 148244 79324 148245 79388
rect 148179 79323 148245 79324
rect 148363 78572 148429 78573
rect 148363 78508 148364 78572
rect 148428 78508 148429 78572
rect 148363 78507 148429 78508
rect 149467 78572 149533 78573
rect 149467 78508 149468 78572
rect 149532 78508 149533 78572
rect 149467 78507 149533 78508
rect 147995 77620 148061 77621
rect 147995 77556 147996 77620
rect 148060 77556 148061 77620
rect 147995 77555 148061 77556
rect 147443 77348 147509 77349
rect 147443 77284 147444 77348
rect 147508 77284 147509 77348
rect 147443 77283 147509 77284
rect 147811 77348 147877 77349
rect 147811 77284 147812 77348
rect 147876 77284 147877 77348
rect 147811 77283 147877 77284
rect 147446 75717 147506 77283
rect 147443 75716 147509 75717
rect 147443 75652 147444 75716
rect 147508 75652 147509 75716
rect 147443 75651 147509 75652
rect 147075 72860 147141 72861
rect 147075 72796 147076 72860
rect 147140 72796 147141 72860
rect 147075 72795 147141 72796
rect 146891 71364 146957 71365
rect 146891 71300 146892 71364
rect 146956 71300 146957 71364
rect 146891 71299 146957 71300
rect 146523 68236 146589 68237
rect 146523 68172 146524 68236
rect 146588 68172 146589 68236
rect 146523 68171 146589 68172
rect 146894 53141 146954 71299
rect 147078 57221 147138 72795
rect 147446 68373 147506 75651
rect 147814 69733 147874 77283
rect 147811 69732 147877 69733
rect 147811 69668 147812 69732
rect 147876 69668 147877 69732
rect 147811 69667 147877 69668
rect 147443 68372 147509 68373
rect 147443 68308 147444 68372
rect 147508 68308 147509 68372
rect 147443 68307 147509 68308
rect 147998 67421 148058 77555
rect 148366 72725 148426 78507
rect 148547 77484 148613 77485
rect 148547 77420 148548 77484
rect 148612 77420 148613 77484
rect 148547 77419 148613 77420
rect 148550 74357 148610 77419
rect 148547 74356 148613 74357
rect 148547 74292 148548 74356
rect 148612 74292 148613 74356
rect 148547 74291 148613 74292
rect 149470 74221 149530 78507
rect 149838 78165 149898 79867
rect 149835 78164 149901 78165
rect 149835 78100 149836 78164
rect 149900 78100 149901 78164
rect 149835 78099 149901 78100
rect 150019 77484 150085 77485
rect 150019 77420 150020 77484
rect 150084 77420 150085 77484
rect 150019 77419 150085 77420
rect 149651 77348 149717 77349
rect 149651 77284 149652 77348
rect 149716 77284 149717 77348
rect 149651 77283 149717 77284
rect 149835 77348 149901 77349
rect 149835 77284 149836 77348
rect 149900 77284 149901 77348
rect 149835 77283 149901 77284
rect 149467 74220 149533 74221
rect 149467 74156 149468 74220
rect 149532 74156 149533 74220
rect 149467 74155 149533 74156
rect 148363 72724 148429 72725
rect 148363 72660 148364 72724
rect 148428 72660 148429 72724
rect 148363 72659 148429 72660
rect 148366 70410 148426 72659
rect 148366 70350 148610 70410
rect 148363 69732 148429 69733
rect 148363 69668 148364 69732
rect 148428 69668 148429 69732
rect 148363 69667 148429 69668
rect 147995 67420 148061 67421
rect 147995 67356 147996 67420
rect 148060 67356 148061 67420
rect 147995 67355 148061 67356
rect 147998 64890 148058 67355
rect 147998 64830 148242 64890
rect 147075 57220 147141 57221
rect 147075 57156 147076 57220
rect 147140 57156 147141 57220
rect 147075 57155 147141 57156
rect 146891 53140 146957 53141
rect 146891 53076 146892 53140
rect 146956 53076 146957 53140
rect 146891 53075 146957 53076
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145419 22676 145485 22677
rect 145419 22612 145420 22676
rect 145484 22612 145485 22676
rect 145419 22611 145485 22612
rect 144315 8940 144381 8941
rect 144315 8876 144316 8940
rect 144380 8876 144381 8940
rect 144315 8875 144381 8876
rect 144131 6220 144197 6221
rect 144131 6156 144132 6220
rect 144196 6156 144197 6220
rect 144131 6155 144197 6156
rect 141294 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 141914 -7066
rect 141294 -7386 141914 -7302
rect 141294 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 141914 -7386
rect 141294 -7654 141914 -7622
rect 145794 3454 146414 38898
rect 148182 30973 148242 64830
rect 148366 45389 148426 69667
rect 148550 62797 148610 70350
rect 149654 68509 149714 77283
rect 149651 68508 149717 68509
rect 149651 68444 149652 68508
rect 149716 68444 149717 68508
rect 149651 68443 149717 68444
rect 149838 67557 149898 77283
rect 149835 67556 149901 67557
rect 149835 67492 149836 67556
rect 149900 67492 149901 67556
rect 149835 67491 149901 67492
rect 148547 62796 148613 62797
rect 148547 62732 148548 62796
rect 148612 62732 148613 62796
rect 148547 62731 148613 62732
rect 150022 60485 150082 77419
rect 150019 60484 150085 60485
rect 150019 60420 150020 60484
rect 150084 60420 150085 60484
rect 150019 60419 150085 60420
rect 148363 45388 148429 45389
rect 148363 45324 148364 45388
rect 148428 45324 148429 45388
rect 148363 45323 148429 45324
rect 150294 43954 150914 78000
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 148179 30972 148245 30973
rect 148179 30908 148180 30972
rect 148244 30908 148245 30972
rect 148179 30907 148245 30908
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 150294 7954 150914 43398
rect 151310 34509 151370 80139
rect 170446 80069 170506 81091
rect 174675 81020 174741 81021
rect 174675 80956 174676 81020
rect 174740 80956 174741 81020
rect 174675 80955 174741 80956
rect 170627 80748 170693 80749
rect 170627 80684 170628 80748
rect 170692 80684 170693 80748
rect 170627 80683 170693 80684
rect 170443 80068 170509 80069
rect 170443 80004 170444 80068
rect 170508 80004 170509 80068
rect 170443 80003 170509 80004
rect 153883 79932 153949 79933
rect 153883 79868 153884 79932
rect 153948 79868 153949 79932
rect 153883 79867 153949 79868
rect 154987 79932 155053 79933
rect 154987 79868 154988 79932
rect 155052 79868 155053 79932
rect 154987 79867 155053 79868
rect 155907 79932 155973 79933
rect 155907 79868 155908 79932
rect 155972 79868 155973 79932
rect 155907 79867 155973 79868
rect 157931 79932 157997 79933
rect 157931 79868 157932 79932
rect 157996 79868 157997 79932
rect 157931 79867 157997 79868
rect 159955 79932 160021 79933
rect 159955 79868 159956 79932
rect 160020 79868 160021 79932
rect 159955 79867 160021 79868
rect 161059 79932 161125 79933
rect 161059 79868 161060 79932
rect 161124 79868 161125 79932
rect 161059 79867 161125 79868
rect 162163 79932 162229 79933
rect 162163 79868 162164 79932
rect 162228 79868 162229 79932
rect 162163 79867 162229 79868
rect 163267 79932 163333 79933
rect 163267 79868 163268 79932
rect 163332 79868 163333 79932
rect 163267 79867 163333 79868
rect 163451 79932 163517 79933
rect 163451 79868 163452 79932
rect 163516 79868 163517 79932
rect 163451 79867 163517 79868
rect 164555 79932 164621 79933
rect 164555 79868 164556 79932
rect 164620 79868 164621 79932
rect 164555 79867 164621 79868
rect 165291 79932 165357 79933
rect 165291 79868 165292 79932
rect 165356 79868 165357 79932
rect 165291 79867 165357 79868
rect 166027 79932 166093 79933
rect 166027 79868 166028 79932
rect 166092 79868 166093 79932
rect 166027 79867 166093 79868
rect 166579 79932 166645 79933
rect 166579 79868 166580 79932
rect 166644 79868 166645 79932
rect 166579 79867 166645 79868
rect 167867 79932 167933 79933
rect 167867 79868 167868 79932
rect 167932 79868 167933 79932
rect 167867 79867 167933 79868
rect 170075 79932 170141 79933
rect 170075 79868 170076 79932
rect 170140 79930 170141 79932
rect 170140 79870 170506 79930
rect 170140 79868 170141 79870
rect 170075 79867 170141 79868
rect 152779 79796 152845 79797
rect 152779 79732 152780 79796
rect 152844 79732 152845 79796
rect 152779 79731 152845 79732
rect 151675 77484 151741 77485
rect 151675 77420 151676 77484
rect 151740 77420 151741 77484
rect 151675 77419 151741 77420
rect 152595 77484 152661 77485
rect 152595 77420 152596 77484
rect 152660 77420 152661 77484
rect 152595 77419 152661 77420
rect 151678 73405 151738 77419
rect 152411 76804 152477 76805
rect 152411 76740 152412 76804
rect 152476 76740 152477 76804
rect 152411 76739 152477 76740
rect 151675 73404 151741 73405
rect 151675 73340 151676 73404
rect 151740 73340 151741 73404
rect 151675 73339 151741 73340
rect 152414 46885 152474 76739
rect 152598 57901 152658 77419
rect 152595 57900 152661 57901
rect 152595 57836 152596 57900
rect 152660 57836 152661 57900
rect 152595 57835 152661 57836
rect 152782 52053 152842 79731
rect 153886 76125 153946 79867
rect 154435 79388 154501 79389
rect 154435 79324 154436 79388
rect 154500 79324 154501 79388
rect 154435 79323 154501 79324
rect 154251 76396 154317 76397
rect 154251 76332 154252 76396
rect 154316 76332 154317 76396
rect 154251 76331 154317 76332
rect 153883 76124 153949 76125
rect 153883 76060 153884 76124
rect 153948 76060 153949 76124
rect 153883 76059 153949 76060
rect 154254 56269 154314 76331
rect 154251 56268 154317 56269
rect 154251 56204 154252 56268
rect 154316 56204 154317 56268
rect 154251 56203 154317 56204
rect 152779 52052 152845 52053
rect 152779 51988 152780 52052
rect 152844 51988 152845 52052
rect 152779 51987 152845 51988
rect 152411 46884 152477 46885
rect 152411 46820 152412 46884
rect 152476 46820 152477 46884
rect 152411 46819 152477 46820
rect 154438 44165 154498 79323
rect 154990 78165 155050 79867
rect 155539 79796 155605 79797
rect 155539 79732 155540 79796
rect 155604 79732 155605 79796
rect 155539 79731 155605 79732
rect 154987 78164 155053 78165
rect 154987 78100 154988 78164
rect 155052 78100 155053 78164
rect 154987 78099 155053 78100
rect 154794 48454 155414 78000
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 154435 44164 154501 44165
rect 154435 44100 154436 44164
rect 154500 44100 154501 44164
rect 154435 44099 154501 44100
rect 151307 34508 151373 34509
rect 151307 34444 151308 34508
rect 151372 34444 151373 34508
rect 151307 34443 151373 34444
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150294 -1306 150914 7398
rect 150294 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 150914 -1306
rect 150294 -1626 150914 -1542
rect 150294 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 150914 -1626
rect 150294 -7654 150914 -1862
rect 154794 12454 155414 47898
rect 155542 38589 155602 79731
rect 155910 79117 155970 79867
rect 156643 79252 156709 79253
rect 156643 79188 156644 79252
rect 156708 79188 156709 79252
rect 156643 79187 156709 79188
rect 155907 79116 155973 79117
rect 155907 79052 155908 79116
rect 155972 79052 155973 79116
rect 155907 79051 155973 79052
rect 155723 78028 155789 78029
rect 155723 77964 155724 78028
rect 155788 77964 155789 78028
rect 155723 77963 155789 77964
rect 155539 38588 155605 38589
rect 155539 38524 155540 38588
rect 155604 38524 155605 38588
rect 155539 38523 155605 38524
rect 155726 17917 155786 77963
rect 156646 64429 156706 79187
rect 157011 78300 157077 78301
rect 157011 78236 157012 78300
rect 157076 78236 157077 78300
rect 157011 78235 157077 78236
rect 156827 75716 156893 75717
rect 156827 75652 156828 75716
rect 156892 75652 156893 75716
rect 156827 75651 156893 75652
rect 156643 64428 156709 64429
rect 156643 64364 156644 64428
rect 156708 64364 156709 64428
rect 156643 64363 156709 64364
rect 156830 52325 156890 75651
rect 156827 52324 156893 52325
rect 156827 52260 156828 52324
rect 156892 52260 156893 52324
rect 156827 52259 156893 52260
rect 157014 37093 157074 78235
rect 157195 75308 157261 75309
rect 157195 75244 157196 75308
rect 157260 75244 157261 75308
rect 157195 75243 157261 75244
rect 157011 37092 157077 37093
rect 157011 37028 157012 37092
rect 157076 37028 157077 37092
rect 157011 37027 157077 37028
rect 157198 35869 157258 75243
rect 157934 56541 157994 79867
rect 158483 79796 158549 79797
rect 158483 79732 158484 79796
rect 158548 79732 158549 79796
rect 158483 79731 158549 79732
rect 158115 79252 158181 79253
rect 158115 79188 158116 79252
rect 158180 79188 158181 79252
rect 158115 79187 158181 79188
rect 157931 56540 157997 56541
rect 157931 56476 157932 56540
rect 157996 56476 157997 56540
rect 157931 56475 157997 56476
rect 158118 53685 158178 79187
rect 158299 78708 158365 78709
rect 158299 78644 158300 78708
rect 158364 78644 158365 78708
rect 158299 78643 158365 78644
rect 158115 53684 158181 53685
rect 158115 53620 158116 53684
rect 158180 53620 158181 53684
rect 158115 53619 158181 53620
rect 158302 50829 158362 78643
rect 158299 50828 158365 50829
rect 158299 50764 158300 50828
rect 158364 50764 158365 50828
rect 158299 50763 158365 50764
rect 157195 35868 157261 35869
rect 157195 35804 157196 35868
rect 157260 35804 157261 35868
rect 157195 35803 157261 35804
rect 158486 21997 158546 79731
rect 158851 78844 158917 78845
rect 158851 78780 158852 78844
rect 158916 78780 158917 78844
rect 158851 78779 158917 78780
rect 158483 21996 158549 21997
rect 158483 21932 158484 21996
rect 158548 21932 158549 21996
rect 158483 21931 158549 21932
rect 158854 21861 158914 78779
rect 159958 78709 160018 79867
rect 159955 78708 160021 78709
rect 159955 78644 159956 78708
rect 160020 78644 160021 78708
rect 159955 78643 160021 78644
rect 159035 75308 159101 75309
rect 159035 75244 159036 75308
rect 159100 75244 159101 75308
rect 159035 75243 159101 75244
rect 158851 21860 158917 21861
rect 158851 21796 158852 21860
rect 158916 21796 158917 21860
rect 158851 21795 158917 21796
rect 159038 21725 159098 75243
rect 159294 52954 159914 78000
rect 160691 76940 160757 76941
rect 160691 76876 160692 76940
rect 160756 76876 160757 76940
rect 160691 76875 160757 76876
rect 160694 63477 160754 76875
rect 160875 76804 160941 76805
rect 160875 76740 160876 76804
rect 160940 76740 160941 76804
rect 160875 76739 160941 76740
rect 160691 63476 160757 63477
rect 160691 63412 160692 63476
rect 160756 63412 160757 63476
rect 160691 63411 160757 63412
rect 160878 55045 160938 76739
rect 160875 55044 160941 55045
rect 160875 54980 160876 55044
rect 160940 54980 160941 55044
rect 160875 54979 160941 54980
rect 161062 53821 161122 79867
rect 161243 79796 161309 79797
rect 161243 79732 161244 79796
rect 161308 79732 161309 79796
rect 161243 79731 161309 79732
rect 161059 53820 161125 53821
rect 161059 53756 161060 53820
rect 161124 53756 161125 53820
rect 161059 53755 161125 53756
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159035 21724 159101 21725
rect 159035 21660 159036 21724
rect 159100 21660 159101 21724
rect 159035 21659 159101 21660
rect 155723 17916 155789 17917
rect 155723 17852 155724 17916
rect 155788 17852 155789 17916
rect 155723 17851 155789 17852
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 154794 -2266 155414 11898
rect 154794 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 155414 -2266
rect 154794 -2586 155414 -2502
rect 154794 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 155414 -2586
rect 154794 -7654 155414 -2822
rect 159294 16954 159914 52398
rect 161246 50557 161306 79731
rect 161243 50556 161309 50557
rect 161243 50492 161244 50556
rect 161308 50492 161309 50556
rect 161243 50491 161309 50492
rect 162166 45253 162226 79867
rect 162531 79796 162597 79797
rect 162531 79732 162532 79796
rect 162596 79732 162597 79796
rect 162531 79731 162597 79732
rect 162347 76804 162413 76805
rect 162347 76740 162348 76804
rect 162412 76740 162413 76804
rect 162347 76739 162413 76740
rect 162350 56405 162410 76739
rect 162347 56404 162413 56405
rect 162347 56340 162348 56404
rect 162412 56340 162413 56404
rect 162347 56339 162413 56340
rect 162534 49605 162594 79731
rect 163270 60621 163330 79867
rect 163267 60620 163333 60621
rect 163267 60556 163268 60620
rect 163332 60556 163333 60620
rect 163267 60555 163333 60556
rect 162531 49604 162597 49605
rect 162531 49540 162532 49604
rect 162596 49540 162597 49604
rect 162531 49539 162597 49540
rect 163454 48109 163514 79867
rect 163635 79660 163701 79661
rect 163635 79596 163636 79660
rect 163700 79596 163701 79660
rect 163635 79595 163701 79596
rect 163451 48108 163517 48109
rect 163451 48044 163452 48108
rect 163516 48044 163517 48108
rect 163451 48043 163517 48044
rect 162163 45252 162229 45253
rect 162163 45188 162164 45252
rect 162228 45188 162229 45252
rect 162163 45187 162229 45188
rect 163638 43893 163698 79595
rect 163794 57454 164414 78000
rect 164558 76941 164618 79867
rect 165107 79796 165173 79797
rect 165107 79732 165108 79796
rect 165172 79732 165173 79796
rect 165107 79731 165173 79732
rect 164923 77348 164989 77349
rect 164923 77284 164924 77348
rect 164988 77284 164989 77348
rect 164923 77283 164989 77284
rect 164555 76940 164621 76941
rect 164555 76876 164556 76940
rect 164620 76876 164621 76940
rect 164555 76875 164621 76876
rect 164926 60349 164986 77283
rect 164923 60348 164989 60349
rect 164923 60284 164924 60348
rect 164988 60284 164989 60348
rect 164923 60283 164989 60284
rect 165110 57493 165170 79731
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 165107 57492 165173 57493
rect 165107 57428 165108 57492
rect 165172 57428 165173 57492
rect 165107 57427 165173 57428
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163635 43892 163701 43893
rect 163635 43828 163636 43892
rect 163700 43828 163701 43892
rect 163635 43827 163701 43828
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 159294 -3226 159914 16398
rect 159294 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 159914 -3226
rect 159294 -3546 159914 -3462
rect 159294 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 159914 -3546
rect 159294 -7654 159914 -3782
rect 163794 21454 164414 56898
rect 165294 50421 165354 79867
rect 166030 76805 166090 79867
rect 166395 79660 166461 79661
rect 166395 79596 166396 79660
rect 166460 79596 166461 79660
rect 166395 79595 166461 79596
rect 165475 76804 165541 76805
rect 165475 76740 165476 76804
rect 165540 76740 165541 76804
rect 165475 76739 165541 76740
rect 166027 76804 166093 76805
rect 166027 76740 166028 76804
rect 166092 76740 166093 76804
rect 166027 76739 166093 76740
rect 165291 50420 165357 50421
rect 165291 50356 165292 50420
rect 165356 50356 165357 50420
rect 165291 50355 165357 50356
rect 165478 26213 165538 76739
rect 166398 55181 166458 79595
rect 166395 55180 166461 55181
rect 166395 55116 166396 55180
rect 166460 55116 166461 55180
rect 166395 55115 166461 55116
rect 166582 45117 166642 79867
rect 166763 79796 166829 79797
rect 166763 79732 166764 79796
rect 166828 79732 166829 79796
rect 166763 79731 166829 79732
rect 167683 79796 167749 79797
rect 167683 79732 167684 79796
rect 167748 79732 167749 79796
rect 167683 79731 167749 79732
rect 166579 45116 166645 45117
rect 166579 45052 166580 45116
rect 166644 45052 166645 45116
rect 166579 45051 166645 45052
rect 166766 44029 166826 79731
rect 167686 46749 167746 79731
rect 167870 76941 167930 79867
rect 168051 79796 168117 79797
rect 168051 79732 168052 79796
rect 168116 79732 168117 79796
rect 168051 79731 168117 79732
rect 170075 79796 170141 79797
rect 170075 79732 170076 79796
rect 170140 79732 170141 79796
rect 170075 79731 170141 79732
rect 167867 76940 167933 76941
rect 167867 76876 167868 76940
rect 167932 76876 167933 76940
rect 167867 76875 167933 76876
rect 167867 76804 167933 76805
rect 167867 76740 167868 76804
rect 167932 76740 167933 76804
rect 167867 76739 167933 76740
rect 167683 46748 167749 46749
rect 167683 46684 167684 46748
rect 167748 46684 167749 46748
rect 167683 46683 167749 46684
rect 167870 46613 167930 76739
rect 167867 46612 167933 46613
rect 167867 46548 167868 46612
rect 167932 46548 167933 46612
rect 167867 46547 167933 46548
rect 166763 44028 166829 44029
rect 166763 43964 166764 44028
rect 166828 43964 166829 44028
rect 166763 43963 166829 43964
rect 168054 43485 168114 79731
rect 169523 79524 169589 79525
rect 169523 79460 169524 79524
rect 169588 79460 169589 79524
rect 169523 79459 169589 79460
rect 168294 61954 168914 78000
rect 169339 76804 169405 76805
rect 169339 76740 169340 76804
rect 169404 76740 169405 76804
rect 169339 76739 169405 76740
rect 168294 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 168914 61954
rect 168294 61634 168914 61718
rect 168294 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 168914 61634
rect 168051 43484 168117 43485
rect 168051 43420 168052 43484
rect 168116 43420 168117 43484
rect 168051 43419 168117 43420
rect 165475 26212 165541 26213
rect 165475 26148 165476 26212
rect 165540 26148 165541 26212
rect 165475 26147 165541 26148
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -4186 164414 20898
rect 163794 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 164414 -4186
rect 163794 -4506 164414 -4422
rect 163794 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 164414 -4506
rect 163794 -7654 164414 -4742
rect 168294 25954 168914 61398
rect 169342 57629 169402 76739
rect 169339 57628 169405 57629
rect 169339 57564 169340 57628
rect 169404 57564 169405 57628
rect 169339 57563 169405 57564
rect 169526 47973 169586 79459
rect 170078 75037 170138 79731
rect 170446 76805 170506 79870
rect 170630 79525 170690 80683
rect 173203 80340 173269 80341
rect 173203 80276 173204 80340
rect 173268 80276 173269 80340
rect 173203 80275 173269 80276
rect 170995 79932 171061 79933
rect 170995 79868 170996 79932
rect 171060 79868 171061 79932
rect 170995 79867 171061 79868
rect 171915 79932 171981 79933
rect 171915 79868 171916 79932
rect 171980 79868 171981 79932
rect 171915 79867 171981 79868
rect 172099 79932 172165 79933
rect 172099 79868 172100 79932
rect 172164 79868 172165 79932
rect 172099 79867 172165 79868
rect 170627 79524 170693 79525
rect 170627 79460 170628 79524
rect 170692 79460 170693 79524
rect 170627 79459 170693 79460
rect 170998 78573 171058 79867
rect 171179 79796 171245 79797
rect 171179 79732 171180 79796
rect 171244 79732 171245 79796
rect 171179 79731 171245 79732
rect 170811 78572 170877 78573
rect 170811 78508 170812 78572
rect 170876 78508 170877 78572
rect 170811 78507 170877 78508
rect 170995 78572 171061 78573
rect 170995 78508 170996 78572
rect 171060 78508 171061 78572
rect 170995 78507 171061 78508
rect 170443 76804 170509 76805
rect 170443 76740 170444 76804
rect 170508 76740 170509 76804
rect 170443 76739 170509 76740
rect 170627 75988 170693 75989
rect 170627 75924 170628 75988
rect 170692 75924 170693 75988
rect 170627 75923 170693 75924
rect 170075 75036 170141 75037
rect 170075 74972 170076 75036
rect 170140 74972 170141 75036
rect 170075 74971 170141 74972
rect 170630 67421 170690 75923
rect 170627 67420 170693 67421
rect 170627 67356 170628 67420
rect 170692 67356 170693 67420
rect 170627 67355 170693 67356
rect 170814 66197 170874 78507
rect 171182 77310 171242 79731
rect 170998 77250 171242 77310
rect 170811 66196 170877 66197
rect 170811 66132 170812 66196
rect 170876 66132 170877 66196
rect 170811 66131 170877 66132
rect 170998 48245 171058 77250
rect 171918 55861 171978 79867
rect 172102 59261 172162 79867
rect 173206 78981 173266 80275
rect 174678 79933 174738 80955
rect 173571 79932 173637 79933
rect 173571 79868 173572 79932
rect 173636 79868 173637 79932
rect 173571 79867 173637 79868
rect 174675 79932 174741 79933
rect 174675 79868 174676 79932
rect 174740 79868 174741 79932
rect 174675 79867 174741 79868
rect 175963 79932 176029 79933
rect 175963 79868 175964 79932
rect 176028 79868 176029 79932
rect 175963 79867 176029 79868
rect 173203 78980 173269 78981
rect 173203 78916 173204 78980
rect 173268 78916 173269 78980
rect 173203 78915 173269 78916
rect 172794 66454 173414 78000
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 172099 59260 172165 59261
rect 172099 59196 172100 59260
rect 172164 59196 172165 59260
rect 172099 59195 172165 59196
rect 171915 55860 171981 55861
rect 171915 55796 171916 55860
rect 171980 55796 171981 55860
rect 171915 55795 171981 55796
rect 170995 48244 171061 48245
rect 170995 48180 170996 48244
rect 171060 48180 171061 48244
rect 170995 48179 171061 48180
rect 169523 47972 169589 47973
rect 169523 47908 169524 47972
rect 169588 47908 169589 47972
rect 169523 47907 169589 47908
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168294 -5146 168914 25398
rect 168294 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 168914 -5146
rect 168294 -5466 168914 -5382
rect 168294 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 168914 -5466
rect 168294 -7654 168914 -5702
rect 172794 30454 173414 65898
rect 173574 62117 173634 79867
rect 174491 79796 174557 79797
rect 174491 79732 174492 79796
rect 174556 79732 174557 79796
rect 174491 79731 174557 79732
rect 173755 79660 173821 79661
rect 173755 79596 173756 79660
rect 173820 79596 173821 79660
rect 173755 79595 173821 79596
rect 173571 62116 173637 62117
rect 173571 62052 173572 62116
rect 173636 62052 173637 62116
rect 173571 62051 173637 62052
rect 173758 44981 173818 79595
rect 174494 64701 174554 79731
rect 175043 79660 175109 79661
rect 175043 79596 175044 79660
rect 175108 79596 175109 79660
rect 175043 79595 175109 79596
rect 174675 77212 174741 77213
rect 174675 77148 174676 77212
rect 174740 77148 174741 77212
rect 174675 77147 174741 77148
rect 174491 64700 174557 64701
rect 174491 64636 174492 64700
rect 174556 64636 174557 64700
rect 174491 64635 174557 64636
rect 174678 63341 174738 77147
rect 174859 76260 174925 76261
rect 174859 76196 174860 76260
rect 174924 76196 174925 76260
rect 174859 76195 174925 76196
rect 174675 63340 174741 63341
rect 174675 63276 174676 63340
rect 174740 63276 174741 63340
rect 174675 63275 174741 63276
rect 174862 52189 174922 76195
rect 174859 52188 174925 52189
rect 174859 52124 174860 52188
rect 174924 52124 174925 52188
rect 174859 52123 174925 52124
rect 175046 45525 175106 79595
rect 175966 57765 176026 79867
rect 176334 79661 176394 81227
rect 176515 80068 176581 80069
rect 176515 80004 176516 80068
rect 176580 80004 176581 80068
rect 176515 80003 176581 80004
rect 176331 79660 176397 79661
rect 176331 79596 176332 79660
rect 176396 79596 176397 79660
rect 176331 79595 176397 79596
rect 176331 78572 176397 78573
rect 176331 78508 176332 78572
rect 176396 78508 176397 78572
rect 176331 78507 176397 78508
rect 176147 77756 176213 77757
rect 176147 77692 176148 77756
rect 176212 77692 176213 77756
rect 176147 77691 176213 77692
rect 175963 57764 176029 57765
rect 175963 57700 175964 57764
rect 176028 57700 176029 57764
rect 175963 57699 176029 57700
rect 176150 50285 176210 77691
rect 176147 50284 176213 50285
rect 176147 50220 176148 50284
rect 176212 50220 176213 50284
rect 176147 50219 176213 50220
rect 176334 49469 176394 78507
rect 176331 49468 176397 49469
rect 176331 49404 176332 49468
rect 176396 49404 176397 49468
rect 176331 49403 176397 49404
rect 175043 45524 175109 45525
rect 175043 45460 175044 45524
rect 175108 45460 175109 45524
rect 175043 45459 175109 45460
rect 173755 44980 173821 44981
rect 173755 44916 173756 44980
rect 173820 44916 173821 44980
rect 173755 44915 173821 44916
rect 176518 37229 176578 80003
rect 177294 70954 177914 78000
rect 177294 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 177914 70954
rect 177294 70634 177914 70718
rect 177294 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 177914 70634
rect 176515 37228 176581 37229
rect 176515 37164 176516 37228
rect 176580 37164 176581 37228
rect 176515 37163 176581 37164
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 172794 -6106 173414 29898
rect 172794 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 173414 -6106
rect 172794 -6426 173414 -6342
rect 172794 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 173414 -6426
rect 172794 -7654 173414 -6662
rect 177294 34954 177914 70398
rect 181302 68781 181362 81499
rect 181794 75454 182414 78000
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181299 68780 181365 68781
rect 181299 68716 181300 68780
rect 181364 68716 181365 68780
rect 181299 68715 181365 68716
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 177294 -7066 177914 34398
rect 177294 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 177914 -7066
rect 177294 -7386 177914 -7302
rect 177294 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 177914 -7386
rect 177294 -7654 177914 -7622
rect 181794 39454 182414 74898
rect 184062 71365 184122 81635
rect 185350 81429 185410 137803
rect 185648 111454 185968 111486
rect 185648 111218 185690 111454
rect 185926 111218 185968 111454
rect 185648 111134 185968 111218
rect 185648 110898 185690 111134
rect 185926 110898 185968 111134
rect 185648 110866 185968 110898
rect 186086 93805 186146 192611
rect 186294 187954 186914 198000
rect 187003 197844 187069 197845
rect 187003 197780 187004 197844
rect 187068 197780 187069 197844
rect 187003 197779 187069 197780
rect 186294 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 186914 187954
rect 186294 187634 186914 187718
rect 186294 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 186914 187634
rect 186294 151954 186914 187398
rect 186294 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 186914 151954
rect 186294 151634 186914 151718
rect 186294 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 186914 151634
rect 186294 142000 186914 151398
rect 186267 140180 186333 140181
rect 186267 140116 186268 140180
rect 186332 140116 186333 140180
rect 186267 140115 186333 140116
rect 186270 93870 186330 140115
rect 186635 138276 186701 138277
rect 186635 138212 186636 138276
rect 186700 138212 186701 138276
rect 186635 138211 186701 138212
rect 186451 138140 186517 138141
rect 186451 138076 186452 138140
rect 186516 138076 186517 138140
rect 186451 138075 186517 138076
rect 186454 136101 186514 138075
rect 186451 136100 186517 136101
rect 186451 136036 186452 136100
rect 186516 136036 186517 136100
rect 186451 136035 186517 136036
rect 186638 135965 186698 138211
rect 186635 135964 186701 135965
rect 186635 135900 186636 135964
rect 186700 135900 186701 135964
rect 186635 135899 186701 135900
rect 186270 93810 186698 93870
rect 186083 93804 186149 93805
rect 186083 93740 186084 93804
rect 186148 93740 186149 93804
rect 186083 93739 186149 93740
rect 186083 90404 186149 90405
rect 186083 90340 186084 90404
rect 186148 90340 186149 90404
rect 186083 90339 186149 90340
rect 186086 84693 186146 90339
rect 186083 84692 186149 84693
rect 186083 84628 186084 84692
rect 186148 84628 186149 84692
rect 186083 84627 186149 84628
rect 186638 84210 186698 93810
rect 186819 84692 186885 84693
rect 186819 84628 186820 84692
rect 186884 84628 186885 84692
rect 186819 84627 186885 84628
rect 186086 84150 186698 84210
rect 185715 81836 185781 81837
rect 185715 81772 185716 81836
rect 185780 81772 185781 81836
rect 185715 81771 185781 81772
rect 185347 81428 185413 81429
rect 185347 81364 185348 81428
rect 185412 81364 185413 81428
rect 185347 81363 185413 81364
rect 185718 80070 185778 81771
rect 186086 81290 186146 84150
rect 186451 82108 186517 82109
rect 186451 82044 186452 82108
rect 186516 82044 186517 82108
rect 186451 82043 186517 82044
rect 186267 81836 186333 81837
rect 186267 81772 186268 81836
rect 186332 81772 186333 81836
rect 186267 81771 186333 81772
rect 186270 81565 186330 81771
rect 186267 81564 186333 81565
rect 186267 81500 186268 81564
rect 186332 81500 186333 81564
rect 186267 81499 186333 81500
rect 186086 81230 186330 81290
rect 185718 80010 185962 80070
rect 185902 75309 185962 80010
rect 186270 79525 186330 81230
rect 186267 79524 186333 79525
rect 186267 79460 186268 79524
rect 186332 79460 186333 79524
rect 186267 79459 186333 79460
rect 186454 79386 186514 82043
rect 186822 81429 186882 84627
rect 186819 81428 186885 81429
rect 186819 81364 186820 81428
rect 186884 81364 186885 81428
rect 186819 81363 186885 81364
rect 186086 79326 186514 79386
rect 185899 75308 185965 75309
rect 185899 75244 185900 75308
rect 185964 75244 185965 75308
rect 185899 75243 185965 75244
rect 185902 74493 185962 75243
rect 185899 74492 185965 74493
rect 185899 74428 185900 74492
rect 185964 74428 185965 74492
rect 185899 74427 185965 74428
rect 184059 71364 184125 71365
rect 184059 71300 184060 71364
rect 184124 71300 184125 71364
rect 184059 71299 184125 71300
rect 186086 64565 186146 79326
rect 186083 64564 186149 64565
rect 186083 64500 186084 64564
rect 186148 64500 186149 64564
rect 186083 64499 186149 64500
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 186294 43954 186914 78000
rect 187006 75173 187066 197779
rect 187190 143445 187250 212467
rect 187742 151333 187802 274619
rect 190794 264454 191414 299898
rect 190794 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 191414 264454
rect 190794 264134 191414 264218
rect 190794 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 191414 264134
rect 189211 262308 189277 262309
rect 189211 262244 189212 262308
rect 189276 262244 189277 262308
rect 189211 262243 189277 262244
rect 189027 198796 189093 198797
rect 189027 198732 189028 198796
rect 189092 198732 189093 198796
rect 189027 198731 189093 198732
rect 187923 198660 187989 198661
rect 187923 198596 187924 198660
rect 187988 198596 187989 198660
rect 187923 198595 187989 198596
rect 187739 151332 187805 151333
rect 187739 151268 187740 151332
rect 187804 151268 187805 151332
rect 187739 151267 187805 151268
rect 187739 149564 187805 149565
rect 187739 149500 187740 149564
rect 187804 149500 187805 149564
rect 187739 149499 187805 149500
rect 187187 143444 187253 143445
rect 187187 143380 187188 143444
rect 187252 143380 187253 143444
rect 187187 143379 187253 143380
rect 187187 138140 187253 138141
rect 187187 138076 187188 138140
rect 187252 138076 187253 138140
rect 187187 138075 187253 138076
rect 187003 75172 187069 75173
rect 187003 75108 187004 75172
rect 187068 75108 187069 75172
rect 187003 75107 187069 75108
rect 187190 64565 187250 138075
rect 187742 80205 187802 149499
rect 187739 80204 187805 80205
rect 187739 80140 187740 80204
rect 187804 80140 187805 80204
rect 187739 80139 187805 80140
rect 187926 76261 187986 198595
rect 188107 197572 188173 197573
rect 188107 197508 188108 197572
rect 188172 197508 188173 197572
rect 188107 197507 188173 197508
rect 188110 77757 188170 197507
rect 188291 139636 188357 139637
rect 188291 139572 188292 139636
rect 188356 139572 188357 139636
rect 188291 139571 188357 139572
rect 188294 138141 188354 139571
rect 188291 138140 188357 138141
rect 188291 138076 188292 138140
rect 188356 138076 188357 138140
rect 188291 138075 188357 138076
rect 189030 80341 189090 198731
rect 189214 144261 189274 262243
rect 190794 262000 191414 263898
rect 195294 707718 195914 711590
rect 195294 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 195914 707718
rect 195294 707398 195914 707482
rect 195294 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 195914 707398
rect 195294 700954 195914 707162
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 664954 195914 700398
rect 195294 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 195914 664954
rect 195294 664634 195914 664718
rect 195294 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 195914 664634
rect 195294 628954 195914 664398
rect 195294 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 195914 628954
rect 195294 628634 195914 628718
rect 195294 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 195914 628634
rect 195294 592954 195914 628398
rect 195294 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 195914 592954
rect 195294 592634 195914 592718
rect 195294 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 195914 592634
rect 195294 556954 195914 592398
rect 195294 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 195914 556954
rect 195294 556634 195914 556718
rect 195294 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 195914 556634
rect 195294 520954 195914 556398
rect 195294 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 195914 520954
rect 195294 520634 195914 520718
rect 195294 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 195914 520634
rect 195294 484954 195914 520398
rect 195294 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 195914 484954
rect 195294 484634 195914 484718
rect 195294 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 195914 484634
rect 195294 448954 195914 484398
rect 195294 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 195914 448954
rect 195294 448634 195914 448718
rect 195294 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 195914 448634
rect 195294 412954 195914 448398
rect 195294 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 195914 412954
rect 195294 412634 195914 412718
rect 195294 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 195914 412634
rect 195294 376954 195914 412398
rect 195294 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 195914 376954
rect 195294 376634 195914 376718
rect 195294 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 195914 376634
rect 195294 340954 195914 376398
rect 195294 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 195914 340954
rect 195294 340634 195914 340718
rect 195294 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 195914 340634
rect 195294 304954 195914 340398
rect 195294 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 195914 304954
rect 195294 304634 195914 304718
rect 195294 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 195914 304634
rect 195294 268954 195914 304398
rect 195294 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 195914 268954
rect 195294 268634 195914 268718
rect 195294 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 195914 268634
rect 193627 262716 193693 262717
rect 193627 262652 193628 262716
rect 193692 262652 193693 262716
rect 193627 262651 193693 262652
rect 193443 262580 193509 262581
rect 193443 262516 193444 262580
rect 193508 262516 193509 262580
rect 193443 262515 193509 262516
rect 190794 192454 191414 198000
rect 193259 196484 193325 196485
rect 193259 196420 193260 196484
rect 193324 196420 193325 196484
rect 193259 196419 193325 196420
rect 190794 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 191414 192454
rect 190794 192134 191414 192218
rect 190794 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 191414 192134
rect 190794 156454 191414 191898
rect 190794 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 191414 156454
rect 190794 156134 191414 156218
rect 190794 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 191414 156134
rect 190499 151468 190565 151469
rect 190499 151404 190500 151468
rect 190564 151404 190565 151468
rect 190499 151403 190565 151404
rect 189579 144668 189645 144669
rect 189579 144604 189580 144668
rect 189644 144604 189645 144668
rect 189579 144603 189645 144604
rect 189211 144260 189277 144261
rect 189211 144196 189212 144260
rect 189276 144196 189277 144260
rect 189211 144195 189277 144196
rect 189395 140044 189461 140045
rect 189395 139980 189396 140044
rect 189460 139980 189461 140044
rect 189395 139979 189461 139980
rect 189027 80340 189093 80341
rect 189027 80276 189028 80340
rect 189092 80276 189093 80340
rect 189027 80275 189093 80276
rect 188291 80204 188357 80205
rect 188291 80140 188292 80204
rect 188356 80140 188357 80204
rect 188291 80139 188357 80140
rect 188107 77756 188173 77757
rect 188107 77692 188108 77756
rect 188172 77692 188173 77756
rect 188107 77691 188173 77692
rect 187923 76260 187989 76261
rect 187923 76196 187924 76260
rect 187988 76196 187989 76260
rect 187923 76195 187989 76196
rect 187926 68917 187986 76195
rect 188294 72453 188354 80139
rect 189398 79389 189458 139979
rect 189395 79388 189461 79389
rect 189395 79324 189396 79388
rect 189460 79324 189461 79388
rect 189395 79323 189461 79324
rect 188291 72452 188357 72453
rect 188291 72388 188292 72452
rect 188356 72388 188357 72452
rect 188291 72387 188357 72388
rect 189582 68917 189642 144603
rect 190502 78301 190562 151403
rect 190794 142000 191414 155898
rect 191971 150516 192037 150517
rect 191971 150452 191972 150516
rect 192036 150452 192037 150516
rect 191971 150451 192037 150452
rect 191603 140452 191669 140453
rect 191603 140388 191604 140452
rect 191668 140388 191669 140452
rect 191603 140387 191669 140388
rect 190867 140316 190933 140317
rect 190867 140252 190868 140316
rect 190932 140252 190933 140316
rect 190867 140251 190933 140252
rect 190870 79253 190930 140251
rect 190867 79252 190933 79253
rect 190867 79188 190868 79252
rect 190932 79188 190933 79252
rect 190867 79187 190933 79188
rect 190499 78300 190565 78301
rect 190499 78236 190500 78300
rect 190564 78236 190565 78300
rect 190499 78235 190565 78236
rect 187923 68916 187989 68917
rect 187923 68852 187924 68916
rect 187988 68852 187989 68916
rect 187923 68851 187989 68852
rect 189579 68916 189645 68917
rect 189579 68852 189580 68916
rect 189644 68852 189645 68916
rect 189579 68851 189645 68852
rect 187187 64564 187253 64565
rect 187187 64500 187188 64564
rect 187252 64500 187253 64564
rect 187187 64499 187253 64500
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 186294 7954 186914 43398
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1306 186914 7398
rect 186294 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 186914 -1306
rect 186294 -1626 186914 -1542
rect 186294 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 186914 -1626
rect 186294 -7654 186914 -1862
rect 190794 48454 191414 78000
rect 191606 76397 191666 140387
rect 191787 139500 191853 139501
rect 191787 139436 191788 139500
rect 191852 139436 191853 139500
rect 191787 139435 191853 139436
rect 191603 76396 191669 76397
rect 191603 76332 191604 76396
rect 191668 76332 191669 76396
rect 191603 76331 191669 76332
rect 191790 59941 191850 139435
rect 191974 76669 192034 150451
rect 192155 147660 192221 147661
rect 192155 147596 192156 147660
rect 192220 147596 192221 147660
rect 192155 147595 192221 147596
rect 192158 81157 192218 147595
rect 192155 81156 192221 81157
rect 192155 81092 192156 81156
rect 192220 81092 192221 81156
rect 192155 81091 192221 81092
rect 191971 76668 192037 76669
rect 191971 76604 191972 76668
rect 192036 76604 192037 76668
rect 191971 76603 192037 76604
rect 191787 59940 191853 59941
rect 191787 59876 191788 59940
rect 191852 59876 191853 59940
rect 191787 59875 191853 59876
rect 193262 52461 193322 196419
rect 193446 144397 193506 262515
rect 193443 144396 193509 144397
rect 193443 144332 193444 144396
rect 193508 144332 193509 144396
rect 193443 144331 193509 144332
rect 193630 144125 193690 262651
rect 195294 232954 195914 268398
rect 199794 708678 200414 711590
rect 199794 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 200414 708678
rect 199794 708358 200414 708442
rect 199794 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 200414 708358
rect 199794 669454 200414 708122
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 197675 265300 197741 265301
rect 197675 265236 197676 265300
rect 197740 265236 197741 265300
rect 197675 265235 197741 265236
rect 197491 265028 197557 265029
rect 197491 264964 197492 265028
rect 197556 264964 197557 265028
rect 197491 264963 197557 264964
rect 195294 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 195914 232954
rect 195294 232634 195914 232718
rect 195294 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 195914 232634
rect 195294 196954 195914 232398
rect 195294 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 195914 196954
rect 197307 196892 197373 196893
rect 197307 196828 197308 196892
rect 197372 196828 197373 196892
rect 197307 196827 197373 196828
rect 195294 196634 195914 196718
rect 195294 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 195914 196634
rect 194547 195396 194613 195397
rect 194547 195332 194548 195396
rect 194612 195332 194613 195396
rect 194547 195331 194613 195332
rect 193811 147388 193877 147389
rect 193811 147324 193812 147388
rect 193876 147324 193877 147388
rect 193811 147323 193877 147324
rect 193627 144124 193693 144125
rect 193627 144060 193628 144124
rect 193692 144060 193693 144124
rect 193627 144059 193693 144060
rect 193814 76805 193874 147323
rect 193995 144804 194061 144805
rect 193995 144740 193996 144804
rect 194060 144740 194061 144804
rect 193995 144739 194061 144740
rect 193811 76804 193877 76805
rect 193811 76740 193812 76804
rect 193876 76740 193877 76804
rect 193811 76739 193877 76740
rect 193259 52460 193325 52461
rect 193259 52396 193260 52460
rect 193324 52396 193325 52460
rect 193259 52395 193325 52396
rect 193998 50557 194058 144739
rect 194550 53821 194610 195331
rect 195294 160954 195914 196398
rect 195294 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 195914 160954
rect 195294 160634 195914 160718
rect 195294 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 195914 160634
rect 194731 147524 194797 147525
rect 194731 147460 194732 147524
rect 194796 147460 194797 147524
rect 194731 147459 194797 147460
rect 194734 79117 194794 147459
rect 195294 124954 195914 160398
rect 196571 147524 196637 147525
rect 196571 147460 196572 147524
rect 196636 147460 196637 147524
rect 196571 147459 196637 147460
rect 196203 147252 196269 147253
rect 196203 147188 196204 147252
rect 196268 147188 196269 147252
rect 196203 147187 196269 147188
rect 196019 146028 196085 146029
rect 196019 145964 196020 146028
rect 196084 145964 196085 146028
rect 196019 145963 196085 145964
rect 195294 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 195914 124954
rect 195294 124634 195914 124718
rect 195294 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 195914 124634
rect 195294 88954 195914 124398
rect 195294 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 195914 88954
rect 195294 88634 195914 88718
rect 195294 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 195914 88634
rect 194731 79116 194797 79117
rect 194731 79052 194732 79116
rect 194796 79052 194797 79116
rect 194731 79051 194797 79052
rect 194547 53820 194613 53821
rect 194547 53756 194548 53820
rect 194612 53756 194613 53820
rect 194547 53755 194613 53756
rect 194550 53141 194610 53755
rect 194547 53140 194613 53141
rect 194547 53076 194548 53140
rect 194612 53076 194613 53140
rect 194547 53075 194613 53076
rect 195294 52954 195914 88398
rect 196022 73677 196082 145963
rect 196206 80885 196266 147187
rect 196203 80884 196269 80885
rect 196203 80820 196204 80884
rect 196268 80820 196269 80884
rect 196203 80819 196269 80820
rect 196019 73676 196085 73677
rect 196019 73612 196020 73676
rect 196084 73612 196085 73676
rect 196019 73611 196085 73612
rect 196574 57357 196634 147459
rect 196571 57356 196637 57357
rect 196571 57292 196572 57356
rect 196636 57292 196637 57356
rect 196571 57291 196637 57292
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 193995 50556 194061 50557
rect 193995 50492 193996 50556
rect 194060 50492 194061 50556
rect 193995 50491 194061 50492
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 190794 12454 191414 47898
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2266 191414 11898
rect 190794 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 191414 -2266
rect 190794 -2586 191414 -2502
rect 190794 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 191414 -2586
rect 190794 -7654 191414 -2822
rect 195294 16954 195914 52398
rect 197310 43893 197370 196827
rect 197494 139773 197554 264963
rect 197678 146845 197738 265235
rect 198963 265164 199029 265165
rect 198963 265100 198964 265164
rect 199028 265100 199029 265164
rect 198963 265099 199029 265100
rect 198779 193084 198845 193085
rect 198779 193020 198780 193084
rect 198844 193020 198845 193084
rect 198779 193019 198845 193020
rect 197859 147116 197925 147117
rect 197859 147052 197860 147116
rect 197924 147052 197925 147116
rect 197859 147051 197925 147052
rect 197675 146844 197741 146845
rect 197675 146780 197676 146844
rect 197740 146780 197741 146844
rect 197675 146779 197741 146780
rect 197675 146164 197741 146165
rect 197675 146100 197676 146164
rect 197740 146100 197741 146164
rect 197675 146099 197741 146100
rect 197491 139772 197557 139773
rect 197491 139708 197492 139772
rect 197556 139708 197557 139772
rect 197491 139707 197557 139708
rect 197678 81293 197738 146099
rect 197675 81292 197741 81293
rect 197675 81228 197676 81292
rect 197740 81228 197741 81292
rect 197675 81227 197741 81228
rect 197862 73949 197922 147051
rect 197859 73948 197925 73949
rect 197859 73884 197860 73948
rect 197924 73884 197925 73948
rect 197859 73883 197925 73884
rect 198782 45117 198842 193019
rect 198966 144533 199026 265099
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199331 195124 199397 195125
rect 199331 195060 199332 195124
rect 199396 195060 199397 195124
rect 199331 195059 199397 195060
rect 199334 146301 199394 195059
rect 199794 165454 200414 200898
rect 204294 709638 204914 711590
rect 204294 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 204914 709638
rect 204294 709318 204914 709402
rect 204294 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 204914 709318
rect 204294 673954 204914 709082
rect 204294 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 204914 673954
rect 204294 673634 204914 673718
rect 204294 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 204914 673634
rect 204294 637954 204914 673398
rect 204294 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 204914 637954
rect 204294 637634 204914 637718
rect 204294 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 204914 637634
rect 204294 601954 204914 637398
rect 204294 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 204914 601954
rect 204294 601634 204914 601718
rect 204294 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 204914 601634
rect 204294 565954 204914 601398
rect 204294 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 204914 565954
rect 204294 565634 204914 565718
rect 204294 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 204914 565634
rect 204294 529954 204914 565398
rect 204294 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 204914 529954
rect 204294 529634 204914 529718
rect 204294 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 204914 529634
rect 204294 493954 204914 529398
rect 204294 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 204914 493954
rect 204294 493634 204914 493718
rect 204294 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 204914 493634
rect 204294 457954 204914 493398
rect 204294 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 204914 457954
rect 204294 457634 204914 457718
rect 204294 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 204914 457634
rect 204294 421954 204914 457398
rect 204294 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 204914 421954
rect 204294 421634 204914 421718
rect 204294 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 204914 421634
rect 204294 385954 204914 421398
rect 204294 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 204914 385954
rect 204294 385634 204914 385718
rect 204294 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 204914 385634
rect 204294 349954 204914 385398
rect 204294 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 204914 349954
rect 204294 349634 204914 349718
rect 204294 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 204914 349634
rect 204294 313954 204914 349398
rect 204294 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 204914 313954
rect 204294 313634 204914 313718
rect 204294 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 204914 313634
rect 204294 277954 204914 313398
rect 204294 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 204914 277954
rect 204294 277634 204914 277718
rect 204294 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 204914 277634
rect 204294 241954 204914 277398
rect 204294 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 204914 241954
rect 204294 241634 204914 241718
rect 204294 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 204914 241634
rect 204294 205954 204914 241398
rect 204294 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 204914 205954
rect 204294 205634 204914 205718
rect 204294 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 204914 205634
rect 200803 199204 200869 199205
rect 200803 199140 200804 199204
rect 200868 199140 200869 199204
rect 200803 199139 200869 199140
rect 200619 199068 200685 199069
rect 200619 199004 200620 199068
rect 200684 199004 200685 199068
rect 200619 199003 200685 199004
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199515 146844 199581 146845
rect 199515 146780 199516 146844
rect 199580 146780 199581 146844
rect 199515 146779 199581 146780
rect 199331 146300 199397 146301
rect 199331 146236 199332 146300
rect 199396 146236 199397 146300
rect 199331 146235 199397 146236
rect 199147 145892 199213 145893
rect 199147 145828 199148 145892
rect 199212 145828 199213 145892
rect 199147 145827 199213 145828
rect 198963 144532 199029 144533
rect 198963 144468 198964 144532
rect 199028 144468 199029 144532
rect 198963 144467 199029 144468
rect 199150 81021 199210 145827
rect 199331 137324 199397 137325
rect 199331 137260 199332 137324
rect 199396 137260 199397 137324
rect 199331 137259 199397 137260
rect 199147 81020 199213 81021
rect 199147 80956 199148 81020
rect 199212 80956 199213 81020
rect 199147 80955 199213 80956
rect 199334 61981 199394 137259
rect 199518 76941 199578 146779
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199515 76940 199581 76941
rect 199515 76876 199516 76940
rect 199580 76876 199581 76940
rect 199515 76875 199581 76876
rect 199331 61980 199397 61981
rect 199331 61916 199332 61980
rect 199396 61916 199397 61980
rect 199331 61915 199397 61916
rect 199794 57454 200414 92898
rect 200622 64701 200682 199003
rect 200806 68917 200866 199139
rect 200987 198932 201053 198933
rect 200987 198868 200988 198932
rect 201052 198868 201053 198932
rect 200987 198867 201053 198868
rect 200990 71365 201050 198867
rect 201171 198388 201237 198389
rect 201171 198324 201172 198388
rect 201236 198324 201237 198388
rect 201171 198323 201237 198324
rect 201174 81429 201234 198323
rect 201723 194580 201789 194581
rect 201723 194516 201724 194580
rect 201788 194516 201789 194580
rect 201723 194515 201789 194516
rect 201539 192948 201605 192949
rect 201539 192884 201540 192948
rect 201604 192884 201605 192948
rect 201539 192883 201605 192884
rect 201171 81428 201237 81429
rect 201171 81364 201172 81428
rect 201236 81364 201237 81428
rect 201171 81363 201237 81364
rect 200987 71364 201053 71365
rect 200987 71300 200988 71364
rect 201052 71300 201053 71364
rect 200987 71299 201053 71300
rect 200803 68916 200869 68917
rect 200803 68852 200804 68916
rect 200868 68852 200869 68916
rect 200803 68851 200869 68852
rect 200619 64700 200685 64701
rect 200619 64636 200620 64700
rect 200684 64636 200685 64700
rect 200619 64635 200685 64636
rect 201355 64700 201421 64701
rect 201355 64636 201356 64700
rect 201420 64636 201421 64700
rect 201355 64635 201421 64636
rect 201358 64157 201418 64635
rect 201355 64156 201421 64157
rect 201355 64092 201356 64156
rect 201420 64092 201421 64156
rect 201355 64091 201421 64092
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 198779 45116 198845 45117
rect 198779 45052 198780 45116
rect 198844 45052 198845 45116
rect 198779 45051 198845 45052
rect 197307 43892 197373 43893
rect 197307 43828 197308 43892
rect 197372 43828 197373 43892
rect 197307 43827 197373 43828
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3226 195914 16398
rect 195294 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 195914 -3226
rect 195294 -3546 195914 -3462
rect 195294 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 195914 -3546
rect 195294 -7654 195914 -3782
rect 199794 21454 200414 56898
rect 201542 43485 201602 192883
rect 201726 46205 201786 194515
rect 201907 193220 201973 193221
rect 201907 193156 201908 193220
rect 201972 193156 201973 193220
rect 201907 193155 201973 193156
rect 201910 52461 201970 193155
rect 204294 169954 204914 205398
rect 208794 710598 209414 711590
rect 208794 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 209414 710598
rect 208794 710278 209414 710362
rect 208794 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 209414 710278
rect 208794 678454 209414 710042
rect 208794 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 209414 678454
rect 208794 678134 209414 678218
rect 208794 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 209414 678134
rect 208794 642454 209414 677898
rect 208794 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 209414 642454
rect 208794 642134 209414 642218
rect 208794 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 209414 642134
rect 208794 606454 209414 641898
rect 208794 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 209414 606454
rect 208794 606134 209414 606218
rect 208794 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 209414 606134
rect 208794 570454 209414 605898
rect 208794 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 209414 570454
rect 208794 570134 209414 570218
rect 208794 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 209414 570134
rect 208794 534454 209414 569898
rect 208794 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 209414 534454
rect 208794 534134 209414 534218
rect 208794 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 209414 534134
rect 208794 498454 209414 533898
rect 208794 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 209414 498454
rect 208794 498134 209414 498218
rect 208794 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 209414 498134
rect 208794 462454 209414 497898
rect 208794 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 209414 462454
rect 208794 462134 209414 462218
rect 208794 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 209414 462134
rect 208794 426454 209414 461898
rect 208794 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 209414 426454
rect 208794 426134 209414 426218
rect 208794 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 209414 426134
rect 208794 390454 209414 425898
rect 208794 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 209414 390454
rect 208794 390134 209414 390218
rect 208794 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 209414 390134
rect 208794 354454 209414 389898
rect 208794 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 209414 354454
rect 208794 354134 209414 354218
rect 208794 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 209414 354134
rect 208794 318454 209414 353898
rect 208794 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 209414 318454
rect 208794 318134 209414 318218
rect 208794 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 209414 318134
rect 208794 282454 209414 317898
rect 208794 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 209414 282454
rect 208794 282134 209414 282218
rect 208794 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 209414 282134
rect 208794 246454 209414 281898
rect 208794 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 209414 246454
rect 208794 246134 209414 246218
rect 208794 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 209414 246134
rect 208794 210454 209414 245898
rect 208794 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 209414 210454
rect 208794 210134 209414 210218
rect 208794 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 209414 210134
rect 207059 200564 207125 200565
rect 207059 200500 207060 200564
rect 207124 200500 207125 200564
rect 207059 200499 207125 200500
rect 204294 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 204914 169954
rect 204294 169634 204914 169718
rect 204294 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 204914 169634
rect 202091 150380 202157 150381
rect 202091 150316 202092 150380
rect 202156 150316 202157 150380
rect 202091 150315 202157 150316
rect 202094 75445 202154 150315
rect 203011 150108 203077 150109
rect 203011 150044 203012 150108
rect 203076 150044 203077 150108
rect 203011 150043 203077 150044
rect 202827 149972 202893 149973
rect 202827 149908 202828 149972
rect 202892 149908 202893 149972
rect 202827 149907 202893 149908
rect 202091 75444 202157 75445
rect 202091 75380 202092 75444
rect 202156 75380 202157 75444
rect 202091 75379 202157 75380
rect 202830 74550 202890 149907
rect 203014 78981 203074 150043
rect 203379 149156 203445 149157
rect 203379 149092 203380 149156
rect 203444 149092 203445 149156
rect 203379 149091 203445 149092
rect 203011 78980 203077 78981
rect 203011 78916 203012 78980
rect 203076 78916 203077 78980
rect 203011 78915 203077 78916
rect 202830 74490 203074 74550
rect 201907 52460 201973 52461
rect 201907 52396 201908 52460
rect 201972 52396 201973 52460
rect 201907 52395 201973 52396
rect 201723 46204 201789 46205
rect 201723 46140 201724 46204
rect 201788 46140 201789 46204
rect 201723 46139 201789 46140
rect 203014 44981 203074 74490
rect 203382 54773 203442 149091
rect 203563 136644 203629 136645
rect 203563 136580 203564 136644
rect 203628 136580 203629 136644
rect 203563 136579 203629 136580
rect 203566 66061 203626 136579
rect 204294 133954 204914 169398
rect 205771 149836 205837 149837
rect 205771 149772 205772 149836
rect 205836 149772 205837 149836
rect 205771 149771 205837 149772
rect 205587 149700 205653 149701
rect 205587 149636 205588 149700
rect 205652 149636 205653 149700
rect 205587 149635 205653 149636
rect 204294 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 204914 133954
rect 204294 133634 204914 133718
rect 204294 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 204914 133634
rect 204294 97954 204914 133398
rect 204294 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 204914 97954
rect 204294 97634 204914 97718
rect 204294 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 204914 97634
rect 203563 66060 203629 66061
rect 203563 65996 203564 66060
rect 203628 65996 203629 66060
rect 203563 65995 203629 65996
rect 204294 61954 204914 97398
rect 205590 79250 205650 149635
rect 205774 80069 205834 149771
rect 205771 80068 205837 80069
rect 205771 80004 205772 80068
rect 205836 80004 205837 80068
rect 205771 80003 205837 80004
rect 205590 79190 205834 79250
rect 205774 72725 205834 79190
rect 205771 72724 205837 72725
rect 205771 72660 205772 72724
rect 205836 72660 205837 72724
rect 205771 72659 205837 72660
rect 204294 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 204914 61954
rect 204294 61634 204914 61718
rect 204294 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 204914 61634
rect 203379 54772 203445 54773
rect 203379 54708 203380 54772
rect 203444 54708 203445 54772
rect 203379 54707 203445 54708
rect 203011 44980 203077 44981
rect 203011 44916 203012 44980
rect 203076 44916 203077 44980
rect 203011 44915 203077 44916
rect 201539 43484 201605 43485
rect 201539 43420 201540 43484
rect 201604 43420 201605 43484
rect 201539 43419 201605 43420
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4186 200414 20898
rect 199794 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 200414 -4186
rect 199794 -4506 200414 -4422
rect 199794 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 200414 -4506
rect 199794 -7654 200414 -4742
rect 204294 25954 204914 61398
rect 207062 50965 207122 200499
rect 208794 174454 209414 209898
rect 213294 711558 213914 711590
rect 213294 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 213914 711558
rect 213294 711238 213914 711322
rect 213294 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 213914 711238
rect 213294 682954 213914 711002
rect 213294 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 213914 682954
rect 213294 682634 213914 682718
rect 213294 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 213914 682634
rect 213294 646954 213914 682398
rect 213294 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 213914 646954
rect 213294 646634 213914 646718
rect 213294 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 213914 646634
rect 213294 610954 213914 646398
rect 213294 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 213914 610954
rect 213294 610634 213914 610718
rect 213294 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 213914 610634
rect 213294 574954 213914 610398
rect 213294 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 213914 574954
rect 213294 574634 213914 574718
rect 213294 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 213914 574634
rect 213294 538954 213914 574398
rect 213294 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 213914 538954
rect 213294 538634 213914 538718
rect 213294 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 213914 538634
rect 213294 502954 213914 538398
rect 213294 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 213914 502954
rect 213294 502634 213914 502718
rect 213294 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 213914 502634
rect 213294 466954 213914 502398
rect 213294 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 213914 466954
rect 213294 466634 213914 466718
rect 213294 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 213914 466634
rect 213294 430954 213914 466398
rect 213294 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 213914 430954
rect 213294 430634 213914 430718
rect 213294 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 213914 430634
rect 213294 394954 213914 430398
rect 213294 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 213914 394954
rect 213294 394634 213914 394718
rect 213294 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 213914 394634
rect 213294 358954 213914 394398
rect 213294 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 213914 358954
rect 213294 358634 213914 358718
rect 213294 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 213914 358634
rect 213294 322954 213914 358398
rect 213294 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 213914 322954
rect 213294 322634 213914 322718
rect 213294 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 213914 322634
rect 213294 286954 213914 322398
rect 213294 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 213914 286954
rect 213294 286634 213914 286718
rect 213294 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 213914 286634
rect 213294 250954 213914 286398
rect 213294 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 213914 250954
rect 213294 250634 213914 250718
rect 213294 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 213914 250634
rect 213294 214954 213914 250398
rect 213294 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 213914 214954
rect 213294 214634 213914 214718
rect 213294 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 213914 214634
rect 210003 194036 210069 194037
rect 210003 193972 210004 194036
rect 210068 193972 210069 194036
rect 210003 193971 210069 193972
rect 209819 193900 209885 193901
rect 209819 193836 209820 193900
rect 209884 193836 209885 193900
rect 209819 193835 209885 193836
rect 208794 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 209414 174454
rect 208794 174134 209414 174218
rect 208794 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 209414 174134
rect 207611 150380 207677 150381
rect 207611 150316 207612 150380
rect 207676 150316 207677 150380
rect 207611 150315 207677 150316
rect 207059 50964 207125 50965
rect 207059 50900 207060 50964
rect 207124 50900 207125 50964
rect 207059 50899 207125 50900
rect 207614 46749 207674 150315
rect 208794 138454 209414 173898
rect 208794 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 209414 138454
rect 208794 138134 209414 138218
rect 208794 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 209414 138134
rect 208794 102454 209414 137898
rect 208794 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 209414 102454
rect 208794 102134 209414 102218
rect 208794 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 209414 102134
rect 208794 66454 209414 101898
rect 208794 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 209414 66454
rect 208794 66134 209414 66218
rect 208794 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 209414 66134
rect 207611 46748 207677 46749
rect 207611 46684 207612 46748
rect 207676 46684 207677 46748
rect 207611 46683 207677 46684
rect 207614 45661 207674 46683
rect 207611 45660 207677 45661
rect 207611 45596 207612 45660
rect 207676 45596 207677 45660
rect 207611 45595 207677 45596
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5146 204914 25398
rect 204294 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 204914 -5146
rect 204294 -5466 204914 -5382
rect 204294 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 204914 -5466
rect 204294 -7654 204914 -5702
rect 208794 30454 209414 65898
rect 209822 50285 209882 193835
rect 210006 77213 210066 193971
rect 213294 178954 213914 214398
rect 213294 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 213914 178954
rect 213294 178634 213914 178718
rect 213294 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 213914 178634
rect 213294 142954 213914 178398
rect 213294 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 213914 142954
rect 213294 142634 213914 142718
rect 213294 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 213914 142634
rect 213294 106954 213914 142398
rect 213294 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 213914 106954
rect 213294 106634 213914 106718
rect 213294 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 213914 106634
rect 210003 77212 210069 77213
rect 210003 77148 210004 77212
rect 210068 77148 210069 77212
rect 210003 77147 210069 77148
rect 213294 70954 213914 106398
rect 213294 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 213914 70954
rect 213294 70634 213914 70718
rect 213294 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 213914 70634
rect 209819 50284 209885 50285
rect 209819 50220 209820 50284
rect 209884 50220 209885 50284
rect 209819 50219 209885 50220
rect 208794 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 209414 30454
rect 208794 30134 209414 30218
rect 208794 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 209414 30134
rect 208794 -6106 209414 29898
rect 208794 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 209414 -6106
rect 208794 -6426 209414 -6342
rect 208794 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 209414 -6426
rect 208794 -7654 209414 -6662
rect 213294 34954 213914 70398
rect 213294 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 213914 34954
rect 213294 34634 213914 34718
rect 213294 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 213914 34634
rect 213294 -7066 213914 34398
rect 213294 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 213914 -7066
rect 213294 -7386 213914 -7302
rect 213294 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 213914 -7386
rect 213294 -7654 213914 -7622
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 222294 705798 222914 711590
rect 222294 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 222914 705798
rect 222294 705478 222914 705562
rect 222294 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 222914 705478
rect 222294 691954 222914 705242
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 655954 222914 691398
rect 222294 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 222914 655954
rect 222294 655634 222914 655718
rect 222294 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 222914 655634
rect 222294 619954 222914 655398
rect 222294 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 222914 619954
rect 222294 619634 222914 619718
rect 222294 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 222914 619634
rect 222294 583954 222914 619398
rect 222294 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 222914 583954
rect 222294 583634 222914 583718
rect 222294 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 222914 583634
rect 222294 547954 222914 583398
rect 222294 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 222914 547954
rect 222294 547634 222914 547718
rect 222294 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 222914 547634
rect 222294 511954 222914 547398
rect 222294 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 222914 511954
rect 222294 511634 222914 511718
rect 222294 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 222914 511634
rect 222294 475954 222914 511398
rect 222294 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 222914 475954
rect 222294 475634 222914 475718
rect 222294 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 222914 475634
rect 222294 439954 222914 475398
rect 222294 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 222914 439954
rect 222294 439634 222914 439718
rect 222294 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 222914 439634
rect 222294 403954 222914 439398
rect 222294 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 222914 403954
rect 222294 403634 222914 403718
rect 222294 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 222914 403634
rect 222294 367954 222914 403398
rect 222294 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 222914 367954
rect 222294 367634 222914 367718
rect 222294 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 222914 367634
rect 222294 331954 222914 367398
rect 222294 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 222914 331954
rect 222294 331634 222914 331718
rect 222294 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 222914 331634
rect 222294 295954 222914 331398
rect 222294 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 222914 295954
rect 222294 295634 222914 295718
rect 222294 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 222914 295634
rect 222294 259954 222914 295398
rect 222294 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 222914 259954
rect 222294 259634 222914 259718
rect 222294 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 222914 259634
rect 222294 223954 222914 259398
rect 222294 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 222914 223954
rect 222294 223634 222914 223718
rect 222294 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 222914 223634
rect 222294 187954 222914 223398
rect 222294 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 222914 187954
rect 222294 187634 222914 187718
rect 222294 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 222914 187634
rect 222294 151954 222914 187398
rect 222294 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 222914 151954
rect 222294 151634 222914 151718
rect 222294 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 222914 151634
rect 222294 115954 222914 151398
rect 222294 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 222914 115954
rect 222294 115634 222914 115718
rect 222294 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 222914 115634
rect 222294 79954 222914 115398
rect 222294 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 222914 79954
rect 222294 79634 222914 79718
rect 222294 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 222914 79634
rect 222294 43954 222914 79398
rect 222294 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 222914 43954
rect 222294 43634 222914 43718
rect 222294 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 222914 43634
rect 222294 7954 222914 43398
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 222294 -1306 222914 7398
rect 222294 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 222914 -1306
rect 222294 -1626 222914 -1542
rect 222294 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 222914 -1626
rect 222294 -7654 222914 -1862
rect 226794 706758 227414 711590
rect 226794 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 227414 706758
rect 226794 706438 227414 706522
rect 226794 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 227414 706438
rect 226794 696454 227414 706202
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 660454 227414 695898
rect 226794 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 227414 660454
rect 226794 660134 227414 660218
rect 226794 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 227414 660134
rect 226794 624454 227414 659898
rect 226794 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 227414 624454
rect 226794 624134 227414 624218
rect 226794 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 227414 624134
rect 226794 588454 227414 623898
rect 226794 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 227414 588454
rect 226794 588134 227414 588218
rect 226794 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 227414 588134
rect 226794 552454 227414 587898
rect 226794 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 227414 552454
rect 226794 552134 227414 552218
rect 226794 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 227414 552134
rect 226794 516454 227414 551898
rect 226794 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 227414 516454
rect 226794 516134 227414 516218
rect 226794 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 227414 516134
rect 226794 480454 227414 515898
rect 226794 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 227414 480454
rect 226794 480134 227414 480218
rect 226794 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 227414 480134
rect 226794 444454 227414 479898
rect 226794 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 227414 444454
rect 226794 444134 227414 444218
rect 226794 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 227414 444134
rect 226794 408454 227414 443898
rect 226794 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 227414 408454
rect 226794 408134 227414 408218
rect 226794 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 227414 408134
rect 226794 372454 227414 407898
rect 226794 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 227414 372454
rect 226794 372134 227414 372218
rect 226794 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 227414 372134
rect 226794 336454 227414 371898
rect 226794 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 227414 336454
rect 226794 336134 227414 336218
rect 226794 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 227414 336134
rect 226794 300454 227414 335898
rect 226794 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 227414 300454
rect 226794 300134 227414 300218
rect 226794 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 227414 300134
rect 226794 264454 227414 299898
rect 226794 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 227414 264454
rect 226794 264134 227414 264218
rect 226794 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 227414 264134
rect 226794 228454 227414 263898
rect 226794 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 227414 228454
rect 226794 228134 227414 228218
rect 226794 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 227414 228134
rect 226794 192454 227414 227898
rect 226794 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 227414 192454
rect 226794 192134 227414 192218
rect 226794 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 227414 192134
rect 226794 156454 227414 191898
rect 226794 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 227414 156454
rect 226794 156134 227414 156218
rect 226794 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 227414 156134
rect 226794 120454 227414 155898
rect 226794 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 227414 120454
rect 226794 120134 227414 120218
rect 226794 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 227414 120134
rect 226794 84454 227414 119898
rect 226794 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 227414 84454
rect 226794 84134 227414 84218
rect 226794 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 227414 84134
rect 226794 48454 227414 83898
rect 226794 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 227414 48454
rect 226794 48134 227414 48218
rect 226794 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 227414 48134
rect 226794 12454 227414 47898
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2266 227414 11898
rect 226794 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 227414 -2266
rect 226794 -2586 227414 -2502
rect 226794 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 227414 -2586
rect 226794 -7654 227414 -2822
rect 231294 707718 231914 711590
rect 231294 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 231914 707718
rect 231294 707398 231914 707482
rect 231294 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 231914 707398
rect 231294 700954 231914 707162
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 664954 231914 700398
rect 231294 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 231914 664954
rect 231294 664634 231914 664718
rect 231294 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 231914 664634
rect 231294 628954 231914 664398
rect 231294 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 231914 628954
rect 231294 628634 231914 628718
rect 231294 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 231914 628634
rect 231294 592954 231914 628398
rect 231294 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 231914 592954
rect 231294 592634 231914 592718
rect 231294 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 231914 592634
rect 231294 556954 231914 592398
rect 231294 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 231914 556954
rect 231294 556634 231914 556718
rect 231294 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 231914 556634
rect 231294 520954 231914 556398
rect 231294 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 231914 520954
rect 231294 520634 231914 520718
rect 231294 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 231914 520634
rect 231294 484954 231914 520398
rect 231294 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 231914 484954
rect 231294 484634 231914 484718
rect 231294 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 231914 484634
rect 231294 448954 231914 484398
rect 231294 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 231914 448954
rect 231294 448634 231914 448718
rect 231294 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 231914 448634
rect 231294 412954 231914 448398
rect 231294 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 231914 412954
rect 231294 412634 231914 412718
rect 231294 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 231914 412634
rect 231294 376954 231914 412398
rect 231294 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 231914 376954
rect 231294 376634 231914 376718
rect 231294 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 231914 376634
rect 231294 340954 231914 376398
rect 231294 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 231914 340954
rect 231294 340634 231914 340718
rect 231294 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 231914 340634
rect 231294 304954 231914 340398
rect 231294 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 231914 304954
rect 231294 304634 231914 304718
rect 231294 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 231914 304634
rect 231294 268954 231914 304398
rect 231294 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 231914 268954
rect 231294 268634 231914 268718
rect 231294 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 231914 268634
rect 231294 232954 231914 268398
rect 231294 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 231914 232954
rect 231294 232634 231914 232718
rect 231294 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 231914 232634
rect 231294 196954 231914 232398
rect 231294 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 231914 196954
rect 231294 196634 231914 196718
rect 231294 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 231914 196634
rect 231294 160954 231914 196398
rect 231294 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 231914 160954
rect 231294 160634 231914 160718
rect 231294 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 231914 160634
rect 231294 124954 231914 160398
rect 231294 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 231914 124954
rect 231294 124634 231914 124718
rect 231294 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 231914 124634
rect 231294 88954 231914 124398
rect 231294 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 231914 88954
rect 231294 88634 231914 88718
rect 231294 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 231914 88634
rect 231294 52954 231914 88398
rect 231294 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 231914 52954
rect 231294 52634 231914 52718
rect 231294 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 231914 52634
rect 231294 16954 231914 52398
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3226 231914 16398
rect 231294 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 231914 -3226
rect 231294 -3546 231914 -3462
rect 231294 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 231914 -3546
rect 231294 -7654 231914 -3782
rect 235794 708678 236414 711590
rect 235794 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 236414 708678
rect 235794 708358 236414 708442
rect 235794 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 236414 708358
rect 235794 669454 236414 708122
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 237454 236414 272898
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4186 236414 20898
rect 235794 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 236414 -4186
rect 235794 -4506 236414 -4422
rect 235794 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 236414 -4506
rect 235794 -7654 236414 -4742
rect 240294 709638 240914 711590
rect 240294 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 240914 709638
rect 240294 709318 240914 709402
rect 240294 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 240914 709318
rect 240294 673954 240914 709082
rect 240294 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 240914 673954
rect 240294 673634 240914 673718
rect 240294 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 240914 673634
rect 240294 637954 240914 673398
rect 240294 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 240914 637954
rect 240294 637634 240914 637718
rect 240294 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 240914 637634
rect 240294 601954 240914 637398
rect 240294 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 240914 601954
rect 240294 601634 240914 601718
rect 240294 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 240914 601634
rect 240294 565954 240914 601398
rect 240294 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 240914 565954
rect 240294 565634 240914 565718
rect 240294 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 240914 565634
rect 240294 529954 240914 565398
rect 240294 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 240914 529954
rect 240294 529634 240914 529718
rect 240294 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 240914 529634
rect 240294 493954 240914 529398
rect 240294 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 240914 493954
rect 240294 493634 240914 493718
rect 240294 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 240914 493634
rect 240294 457954 240914 493398
rect 240294 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 240914 457954
rect 240294 457634 240914 457718
rect 240294 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 240914 457634
rect 240294 421954 240914 457398
rect 240294 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 240914 421954
rect 240294 421634 240914 421718
rect 240294 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 240914 421634
rect 240294 385954 240914 421398
rect 240294 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 240914 385954
rect 240294 385634 240914 385718
rect 240294 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 240914 385634
rect 240294 349954 240914 385398
rect 240294 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 240914 349954
rect 240294 349634 240914 349718
rect 240294 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 240914 349634
rect 240294 313954 240914 349398
rect 240294 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 240914 313954
rect 240294 313634 240914 313718
rect 240294 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 240914 313634
rect 240294 277954 240914 313398
rect 240294 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 240914 277954
rect 240294 277634 240914 277718
rect 240294 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 240914 277634
rect 240294 241954 240914 277398
rect 240294 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 240914 241954
rect 240294 241634 240914 241718
rect 240294 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 240914 241634
rect 240294 205954 240914 241398
rect 240294 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 240914 205954
rect 240294 205634 240914 205718
rect 240294 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 240914 205634
rect 240294 169954 240914 205398
rect 240294 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 240914 169954
rect 240294 169634 240914 169718
rect 240294 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 240914 169634
rect 240294 133954 240914 169398
rect 240294 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 240914 133954
rect 240294 133634 240914 133718
rect 240294 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 240914 133634
rect 240294 97954 240914 133398
rect 240294 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 240914 97954
rect 240294 97634 240914 97718
rect 240294 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 240914 97634
rect 240294 61954 240914 97398
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 25954 240914 61398
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 240294 -5146 240914 25398
rect 240294 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 240914 -5146
rect 240294 -5466 240914 -5382
rect 240294 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 240914 -5466
rect 240294 -7654 240914 -5702
rect 244794 710598 245414 711590
rect 244794 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 245414 710598
rect 244794 710278 245414 710362
rect 244794 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 245414 710278
rect 244794 678454 245414 710042
rect 244794 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 245414 678454
rect 244794 678134 245414 678218
rect 244794 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 245414 678134
rect 244794 642454 245414 677898
rect 244794 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 245414 642454
rect 244794 642134 245414 642218
rect 244794 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 245414 642134
rect 244794 606454 245414 641898
rect 244794 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 245414 606454
rect 244794 606134 245414 606218
rect 244794 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 245414 606134
rect 244794 570454 245414 605898
rect 244794 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 245414 570454
rect 244794 570134 245414 570218
rect 244794 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 245414 570134
rect 244794 534454 245414 569898
rect 244794 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 245414 534454
rect 244794 534134 245414 534218
rect 244794 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 245414 534134
rect 244794 498454 245414 533898
rect 244794 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 245414 498454
rect 244794 498134 245414 498218
rect 244794 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 245414 498134
rect 244794 462454 245414 497898
rect 244794 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 245414 462454
rect 244794 462134 245414 462218
rect 244794 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 245414 462134
rect 244794 426454 245414 461898
rect 244794 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 245414 426454
rect 244794 426134 245414 426218
rect 244794 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 245414 426134
rect 244794 390454 245414 425898
rect 244794 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 245414 390454
rect 244794 390134 245414 390218
rect 244794 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 245414 390134
rect 244794 354454 245414 389898
rect 244794 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 245414 354454
rect 244794 354134 245414 354218
rect 244794 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 245414 354134
rect 244794 318454 245414 353898
rect 244794 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 245414 318454
rect 244794 318134 245414 318218
rect 244794 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 245414 318134
rect 244794 282454 245414 317898
rect 244794 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 245414 282454
rect 244794 282134 245414 282218
rect 244794 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 245414 282134
rect 244794 246454 245414 281898
rect 244794 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 245414 246454
rect 244794 246134 245414 246218
rect 244794 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 245414 246134
rect 244794 210454 245414 245898
rect 244794 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 245414 210454
rect 244794 210134 245414 210218
rect 244794 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 245414 210134
rect 244794 174454 245414 209898
rect 244794 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 245414 174454
rect 244794 174134 245414 174218
rect 244794 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 245414 174134
rect 244794 138454 245414 173898
rect 244794 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 245414 138454
rect 244794 138134 245414 138218
rect 244794 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 245414 138134
rect 244794 102454 245414 137898
rect 244794 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 245414 102454
rect 244794 102134 245414 102218
rect 244794 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 245414 102134
rect 244794 66454 245414 101898
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 30454 245414 65898
rect 244794 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 245414 30454
rect 244794 30134 245414 30218
rect 244794 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 245414 30134
rect 244794 -6106 245414 29898
rect 244794 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 245414 -6106
rect 244794 -6426 245414 -6342
rect 244794 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 245414 -6426
rect 244794 -7654 245414 -6662
rect 249294 711558 249914 711590
rect 249294 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 249914 711558
rect 249294 711238 249914 711322
rect 249294 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 249914 711238
rect 249294 682954 249914 711002
rect 249294 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 249914 682954
rect 249294 682634 249914 682718
rect 249294 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 249914 682634
rect 249294 646954 249914 682398
rect 249294 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 249914 646954
rect 249294 646634 249914 646718
rect 249294 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 249914 646634
rect 249294 610954 249914 646398
rect 249294 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 249914 610954
rect 249294 610634 249914 610718
rect 249294 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 249914 610634
rect 249294 574954 249914 610398
rect 249294 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 249914 574954
rect 249294 574634 249914 574718
rect 249294 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 249914 574634
rect 249294 538954 249914 574398
rect 249294 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 249914 538954
rect 249294 538634 249914 538718
rect 249294 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 249914 538634
rect 249294 502954 249914 538398
rect 249294 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 249914 502954
rect 249294 502634 249914 502718
rect 249294 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 249914 502634
rect 249294 466954 249914 502398
rect 249294 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 249914 466954
rect 249294 466634 249914 466718
rect 249294 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 249914 466634
rect 249294 430954 249914 466398
rect 249294 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 249914 430954
rect 249294 430634 249914 430718
rect 249294 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 249914 430634
rect 249294 394954 249914 430398
rect 249294 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 249914 394954
rect 249294 394634 249914 394718
rect 249294 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 249914 394634
rect 249294 358954 249914 394398
rect 249294 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 249914 358954
rect 249294 358634 249914 358718
rect 249294 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 249914 358634
rect 249294 322954 249914 358398
rect 249294 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 249914 322954
rect 249294 322634 249914 322718
rect 249294 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 249914 322634
rect 249294 286954 249914 322398
rect 249294 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 249914 286954
rect 249294 286634 249914 286718
rect 249294 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 249914 286634
rect 249294 250954 249914 286398
rect 249294 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 249914 250954
rect 249294 250634 249914 250718
rect 249294 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 249914 250634
rect 249294 214954 249914 250398
rect 249294 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 249914 214954
rect 249294 214634 249914 214718
rect 249294 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 249914 214634
rect 249294 178954 249914 214398
rect 249294 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 249914 178954
rect 249294 178634 249914 178718
rect 249294 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 249914 178634
rect 249294 142954 249914 178398
rect 249294 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 249914 142954
rect 249294 142634 249914 142718
rect 249294 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 249914 142634
rect 249294 106954 249914 142398
rect 249294 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 249914 106954
rect 249294 106634 249914 106718
rect 249294 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 249914 106634
rect 249294 70954 249914 106398
rect 249294 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 249914 70954
rect 249294 70634 249914 70718
rect 249294 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 249914 70634
rect 249294 34954 249914 70398
rect 249294 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 249914 34954
rect 249294 34634 249914 34718
rect 249294 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 249914 34634
rect 249294 -7066 249914 34398
rect 249294 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 249914 -7066
rect 249294 -7386 249914 -7302
rect 249294 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 249914 -7386
rect 249294 -7654 249914 -7622
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 258294 705798 258914 711590
rect 258294 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 258914 705798
rect 258294 705478 258914 705562
rect 258294 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 258914 705478
rect 258294 691954 258914 705242
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 655954 258914 691398
rect 258294 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 258914 655954
rect 258294 655634 258914 655718
rect 258294 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 258914 655634
rect 258294 619954 258914 655398
rect 258294 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 258914 619954
rect 258294 619634 258914 619718
rect 258294 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 258914 619634
rect 258294 583954 258914 619398
rect 258294 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 258914 583954
rect 258294 583634 258914 583718
rect 258294 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 258914 583634
rect 258294 547954 258914 583398
rect 258294 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 258914 547954
rect 258294 547634 258914 547718
rect 258294 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 258914 547634
rect 258294 511954 258914 547398
rect 258294 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 258914 511954
rect 258294 511634 258914 511718
rect 258294 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 258914 511634
rect 258294 475954 258914 511398
rect 258294 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 258914 475954
rect 258294 475634 258914 475718
rect 258294 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 258914 475634
rect 258294 439954 258914 475398
rect 258294 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 258914 439954
rect 258294 439634 258914 439718
rect 258294 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 258914 439634
rect 258294 403954 258914 439398
rect 258294 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 258914 403954
rect 258294 403634 258914 403718
rect 258294 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 258914 403634
rect 258294 367954 258914 403398
rect 258294 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 258914 367954
rect 258294 367634 258914 367718
rect 258294 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 258914 367634
rect 258294 331954 258914 367398
rect 258294 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 258914 331954
rect 258294 331634 258914 331718
rect 258294 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 258914 331634
rect 258294 295954 258914 331398
rect 258294 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 258914 295954
rect 258294 295634 258914 295718
rect 258294 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 258914 295634
rect 258294 259954 258914 295398
rect 258294 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 258914 259954
rect 258294 259634 258914 259718
rect 258294 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 258914 259634
rect 258294 223954 258914 259398
rect 258294 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 258914 223954
rect 258294 223634 258914 223718
rect 258294 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 258914 223634
rect 258294 187954 258914 223398
rect 258294 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 258914 187954
rect 258294 187634 258914 187718
rect 258294 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 258914 187634
rect 258294 151954 258914 187398
rect 258294 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 258914 151954
rect 258294 151634 258914 151718
rect 258294 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 258914 151634
rect 258294 115954 258914 151398
rect 258294 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 258914 115954
rect 258294 115634 258914 115718
rect 258294 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 258914 115634
rect 258294 79954 258914 115398
rect 258294 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 258914 79954
rect 258294 79634 258914 79718
rect 258294 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 258914 79634
rect 258294 43954 258914 79398
rect 258294 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 258914 43954
rect 258294 43634 258914 43718
rect 258294 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 258914 43634
rect 258294 7954 258914 43398
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258294 -1306 258914 7398
rect 258294 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 258914 -1306
rect 258294 -1626 258914 -1542
rect 258294 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 258914 -1626
rect 258294 -7654 258914 -1862
rect 262794 706758 263414 711590
rect 262794 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 263414 706758
rect 262794 706438 263414 706522
rect 262794 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 263414 706438
rect 262794 696454 263414 706202
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 660454 263414 695898
rect 262794 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 263414 660454
rect 262794 660134 263414 660218
rect 262794 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 263414 660134
rect 262794 624454 263414 659898
rect 262794 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 263414 624454
rect 262794 624134 263414 624218
rect 262794 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 263414 624134
rect 262794 588454 263414 623898
rect 262794 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 263414 588454
rect 262794 588134 263414 588218
rect 262794 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 263414 588134
rect 262794 552454 263414 587898
rect 262794 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 263414 552454
rect 262794 552134 263414 552218
rect 262794 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 263414 552134
rect 262794 516454 263414 551898
rect 262794 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 263414 516454
rect 262794 516134 263414 516218
rect 262794 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 263414 516134
rect 262794 480454 263414 515898
rect 262794 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 263414 480454
rect 262794 480134 263414 480218
rect 262794 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 263414 480134
rect 262794 444454 263414 479898
rect 262794 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 263414 444454
rect 262794 444134 263414 444218
rect 262794 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 263414 444134
rect 262794 408454 263414 443898
rect 262794 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 263414 408454
rect 262794 408134 263414 408218
rect 262794 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 263414 408134
rect 262794 372454 263414 407898
rect 262794 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 263414 372454
rect 262794 372134 263414 372218
rect 262794 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 263414 372134
rect 262794 336454 263414 371898
rect 262794 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 263414 336454
rect 262794 336134 263414 336218
rect 262794 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 263414 336134
rect 262794 300454 263414 335898
rect 262794 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 263414 300454
rect 262794 300134 263414 300218
rect 262794 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 263414 300134
rect 262794 264454 263414 299898
rect 262794 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 263414 264454
rect 262794 264134 263414 264218
rect 262794 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 263414 264134
rect 262794 228454 263414 263898
rect 262794 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 263414 228454
rect 262794 228134 263414 228218
rect 262794 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 263414 228134
rect 262794 192454 263414 227898
rect 262794 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 263414 192454
rect 262794 192134 263414 192218
rect 262794 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 263414 192134
rect 262794 156454 263414 191898
rect 262794 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 263414 156454
rect 262794 156134 263414 156218
rect 262794 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 263414 156134
rect 262794 120454 263414 155898
rect 262794 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 263414 120454
rect 262794 120134 263414 120218
rect 262794 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 263414 120134
rect 262794 84454 263414 119898
rect 262794 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 263414 84454
rect 262794 84134 263414 84218
rect 262794 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 263414 84134
rect 262794 48454 263414 83898
rect 262794 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 263414 48454
rect 262794 48134 263414 48218
rect 262794 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 263414 48134
rect 262794 12454 263414 47898
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2266 263414 11898
rect 262794 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 263414 -2266
rect 262794 -2586 263414 -2502
rect 262794 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 263414 -2586
rect 262794 -7654 263414 -2822
rect 267294 707718 267914 711590
rect 267294 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 267914 707718
rect 267294 707398 267914 707482
rect 267294 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 267914 707398
rect 267294 700954 267914 707162
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 664954 267914 700398
rect 267294 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 267914 664954
rect 267294 664634 267914 664718
rect 267294 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 267914 664634
rect 267294 628954 267914 664398
rect 267294 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 267914 628954
rect 267294 628634 267914 628718
rect 267294 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 267914 628634
rect 267294 592954 267914 628398
rect 267294 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 267914 592954
rect 267294 592634 267914 592718
rect 267294 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 267914 592634
rect 267294 556954 267914 592398
rect 267294 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 267914 556954
rect 267294 556634 267914 556718
rect 267294 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 267914 556634
rect 267294 520954 267914 556398
rect 267294 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 267914 520954
rect 267294 520634 267914 520718
rect 267294 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 267914 520634
rect 267294 484954 267914 520398
rect 267294 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 267914 484954
rect 267294 484634 267914 484718
rect 267294 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 267914 484634
rect 267294 448954 267914 484398
rect 267294 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 267914 448954
rect 267294 448634 267914 448718
rect 267294 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 267914 448634
rect 267294 412954 267914 448398
rect 267294 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 267914 412954
rect 267294 412634 267914 412718
rect 267294 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 267914 412634
rect 267294 376954 267914 412398
rect 267294 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 267914 376954
rect 267294 376634 267914 376718
rect 267294 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 267914 376634
rect 267294 340954 267914 376398
rect 267294 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 267914 340954
rect 267294 340634 267914 340718
rect 267294 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 267914 340634
rect 267294 304954 267914 340398
rect 267294 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 267914 304954
rect 267294 304634 267914 304718
rect 267294 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 267914 304634
rect 267294 268954 267914 304398
rect 267294 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 267914 268954
rect 267294 268634 267914 268718
rect 267294 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 267914 268634
rect 267294 232954 267914 268398
rect 267294 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 267914 232954
rect 267294 232634 267914 232718
rect 267294 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 267914 232634
rect 267294 196954 267914 232398
rect 267294 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 267914 196954
rect 267294 196634 267914 196718
rect 267294 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 267914 196634
rect 267294 160954 267914 196398
rect 267294 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 267914 160954
rect 267294 160634 267914 160718
rect 267294 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 267914 160634
rect 267294 124954 267914 160398
rect 267294 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 267914 124954
rect 267294 124634 267914 124718
rect 267294 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 267914 124634
rect 267294 88954 267914 124398
rect 267294 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 267914 88954
rect 267294 88634 267914 88718
rect 267294 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 267914 88634
rect 267294 52954 267914 88398
rect 267294 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 267914 52954
rect 267294 52634 267914 52718
rect 267294 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 267914 52634
rect 267294 16954 267914 52398
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3226 267914 16398
rect 267294 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 267914 -3226
rect 267294 -3546 267914 -3462
rect 267294 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 267914 -3546
rect 267294 -7654 267914 -3782
rect 271794 708678 272414 711590
rect 271794 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 272414 708678
rect 271794 708358 272414 708442
rect 271794 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 272414 708358
rect 271794 669454 272414 708122
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4186 272414 20898
rect 271794 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 272414 -4186
rect 271794 -4506 272414 -4422
rect 271794 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 272414 -4506
rect 271794 -7654 272414 -4742
rect 276294 709638 276914 711590
rect 276294 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 276914 709638
rect 276294 709318 276914 709402
rect 276294 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 276914 709318
rect 276294 673954 276914 709082
rect 276294 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 276914 673954
rect 276294 673634 276914 673718
rect 276294 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 276914 673634
rect 276294 637954 276914 673398
rect 276294 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 276914 637954
rect 276294 637634 276914 637718
rect 276294 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 276914 637634
rect 276294 601954 276914 637398
rect 276294 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 276914 601954
rect 276294 601634 276914 601718
rect 276294 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 276914 601634
rect 276294 565954 276914 601398
rect 276294 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 276914 565954
rect 276294 565634 276914 565718
rect 276294 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 276914 565634
rect 276294 529954 276914 565398
rect 276294 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 276914 529954
rect 276294 529634 276914 529718
rect 276294 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 276914 529634
rect 276294 493954 276914 529398
rect 276294 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 276914 493954
rect 276294 493634 276914 493718
rect 276294 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 276914 493634
rect 276294 457954 276914 493398
rect 276294 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 276914 457954
rect 276294 457634 276914 457718
rect 276294 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 276914 457634
rect 276294 421954 276914 457398
rect 276294 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 276914 421954
rect 276294 421634 276914 421718
rect 276294 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 276914 421634
rect 276294 385954 276914 421398
rect 276294 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 276914 385954
rect 276294 385634 276914 385718
rect 276294 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 276914 385634
rect 276294 349954 276914 385398
rect 276294 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 276914 349954
rect 276294 349634 276914 349718
rect 276294 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 276914 349634
rect 276294 313954 276914 349398
rect 276294 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 276914 313954
rect 276294 313634 276914 313718
rect 276294 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 276914 313634
rect 276294 277954 276914 313398
rect 276294 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 276914 277954
rect 276294 277634 276914 277718
rect 276294 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 276914 277634
rect 276294 241954 276914 277398
rect 276294 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 276914 241954
rect 276294 241634 276914 241718
rect 276294 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 276914 241634
rect 276294 205954 276914 241398
rect 276294 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 276914 205954
rect 276294 205634 276914 205718
rect 276294 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 276914 205634
rect 276294 169954 276914 205398
rect 276294 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 276914 169954
rect 276294 169634 276914 169718
rect 276294 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 276914 169634
rect 276294 133954 276914 169398
rect 276294 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 276914 133954
rect 276294 133634 276914 133718
rect 276294 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 276914 133634
rect 276294 97954 276914 133398
rect 276294 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 276914 97954
rect 276294 97634 276914 97718
rect 276294 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 276914 97634
rect 276294 61954 276914 97398
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 25954 276914 61398
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 276294 -5146 276914 25398
rect 276294 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 276914 -5146
rect 276294 -5466 276914 -5382
rect 276294 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 276914 -5466
rect 276294 -7654 276914 -5702
rect 280794 710598 281414 711590
rect 280794 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 281414 710598
rect 280794 710278 281414 710362
rect 280794 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 281414 710278
rect 280794 678454 281414 710042
rect 280794 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 281414 678454
rect 280794 678134 281414 678218
rect 280794 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 281414 678134
rect 280794 642454 281414 677898
rect 280794 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 281414 642454
rect 280794 642134 281414 642218
rect 280794 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 281414 642134
rect 280794 606454 281414 641898
rect 280794 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 281414 606454
rect 280794 606134 281414 606218
rect 280794 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 281414 606134
rect 280794 570454 281414 605898
rect 280794 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 281414 570454
rect 280794 570134 281414 570218
rect 280794 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 281414 570134
rect 280794 534454 281414 569898
rect 280794 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 281414 534454
rect 280794 534134 281414 534218
rect 280794 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 281414 534134
rect 280794 498454 281414 533898
rect 280794 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 281414 498454
rect 280794 498134 281414 498218
rect 280794 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 281414 498134
rect 280794 462454 281414 497898
rect 280794 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 281414 462454
rect 280794 462134 281414 462218
rect 280794 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 281414 462134
rect 280794 426454 281414 461898
rect 280794 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 281414 426454
rect 280794 426134 281414 426218
rect 280794 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 281414 426134
rect 280794 390454 281414 425898
rect 280794 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 281414 390454
rect 280794 390134 281414 390218
rect 280794 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 281414 390134
rect 280794 354454 281414 389898
rect 280794 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 281414 354454
rect 280794 354134 281414 354218
rect 280794 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 281414 354134
rect 280794 318454 281414 353898
rect 280794 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 281414 318454
rect 280794 318134 281414 318218
rect 280794 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 281414 318134
rect 280794 282454 281414 317898
rect 280794 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 281414 282454
rect 280794 282134 281414 282218
rect 280794 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 281414 282134
rect 280794 246454 281414 281898
rect 280794 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 281414 246454
rect 280794 246134 281414 246218
rect 280794 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 281414 246134
rect 280794 210454 281414 245898
rect 280794 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 281414 210454
rect 280794 210134 281414 210218
rect 280794 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 281414 210134
rect 280794 174454 281414 209898
rect 280794 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 281414 174454
rect 280794 174134 281414 174218
rect 280794 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 281414 174134
rect 280794 138454 281414 173898
rect 280794 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 281414 138454
rect 280794 138134 281414 138218
rect 280794 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 281414 138134
rect 280794 102454 281414 137898
rect 280794 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 281414 102454
rect 280794 102134 281414 102218
rect 280794 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 281414 102134
rect 280794 66454 281414 101898
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 30454 281414 65898
rect 280794 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 281414 30454
rect 280794 30134 281414 30218
rect 280794 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 281414 30134
rect 280794 -6106 281414 29898
rect 280794 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 281414 -6106
rect 280794 -6426 281414 -6342
rect 280794 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 281414 -6426
rect 280794 -7654 281414 -6662
rect 285294 711558 285914 711590
rect 285294 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 285914 711558
rect 285294 711238 285914 711322
rect 285294 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 285914 711238
rect 285294 682954 285914 711002
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 285294 646954 285914 682398
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 285294 610954 285914 646398
rect 285294 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 285914 610954
rect 285294 610634 285914 610718
rect 285294 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 285914 610634
rect 285294 574954 285914 610398
rect 285294 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 285914 574954
rect 285294 574634 285914 574718
rect 285294 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 285914 574634
rect 285294 538954 285914 574398
rect 285294 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 285914 538954
rect 285294 538634 285914 538718
rect 285294 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 285914 538634
rect 285294 502954 285914 538398
rect 285294 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 285914 502954
rect 285294 502634 285914 502718
rect 285294 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 285914 502634
rect 285294 466954 285914 502398
rect 285294 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 285914 466954
rect 285294 466634 285914 466718
rect 285294 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 285914 466634
rect 285294 430954 285914 466398
rect 285294 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 285914 430954
rect 285294 430634 285914 430718
rect 285294 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 285914 430634
rect 285294 394954 285914 430398
rect 285294 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 285914 394954
rect 285294 394634 285914 394718
rect 285294 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 285914 394634
rect 285294 358954 285914 394398
rect 285294 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 285914 358954
rect 285294 358634 285914 358718
rect 285294 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 285914 358634
rect 285294 322954 285914 358398
rect 285294 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 285914 322954
rect 285294 322634 285914 322718
rect 285294 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 285914 322634
rect 285294 286954 285914 322398
rect 285294 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 285914 286954
rect 285294 286634 285914 286718
rect 285294 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 285914 286634
rect 285294 250954 285914 286398
rect 285294 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 285914 250954
rect 285294 250634 285914 250718
rect 285294 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 285914 250634
rect 285294 214954 285914 250398
rect 285294 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 285914 214954
rect 285294 214634 285914 214718
rect 285294 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 285914 214634
rect 285294 178954 285914 214398
rect 285294 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 285914 178954
rect 285294 178634 285914 178718
rect 285294 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 285914 178634
rect 285294 142954 285914 178398
rect 285294 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 285914 142954
rect 285294 142634 285914 142718
rect 285294 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 285914 142634
rect 285294 106954 285914 142398
rect 285294 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 285914 106954
rect 285294 106634 285914 106718
rect 285294 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 285914 106634
rect 285294 70954 285914 106398
rect 285294 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 285914 70954
rect 285294 70634 285914 70718
rect 285294 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 285914 70634
rect 285294 34954 285914 70398
rect 285294 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 285914 34954
rect 285294 34634 285914 34718
rect 285294 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 285914 34634
rect 285294 -7066 285914 34398
rect 285294 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 285914 -7066
rect 285294 -7386 285914 -7302
rect 285294 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 285914 -7386
rect 285294 -7654 285914 -7622
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 294294 705798 294914 711590
rect 294294 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 294914 705798
rect 294294 705478 294914 705562
rect 294294 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 294914 705478
rect 294294 691954 294914 705242
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 619954 294914 655398
rect 294294 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 294914 619954
rect 294294 619634 294914 619718
rect 294294 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 294914 619634
rect 294294 583954 294914 619398
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 294294 547954 294914 583398
rect 294294 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 294914 547954
rect 294294 547634 294914 547718
rect 294294 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 294914 547634
rect 294294 511954 294914 547398
rect 294294 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 294914 511954
rect 294294 511634 294914 511718
rect 294294 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 294914 511634
rect 294294 475954 294914 511398
rect 294294 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 294914 475954
rect 294294 475634 294914 475718
rect 294294 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 294914 475634
rect 294294 439954 294914 475398
rect 294294 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 294914 439954
rect 294294 439634 294914 439718
rect 294294 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 294914 439634
rect 294294 403954 294914 439398
rect 294294 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 294914 403954
rect 294294 403634 294914 403718
rect 294294 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 294914 403634
rect 294294 367954 294914 403398
rect 294294 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 294914 367954
rect 294294 367634 294914 367718
rect 294294 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 294914 367634
rect 294294 331954 294914 367398
rect 294294 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 294914 331954
rect 294294 331634 294914 331718
rect 294294 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 294914 331634
rect 294294 295954 294914 331398
rect 294294 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 294914 295954
rect 294294 295634 294914 295718
rect 294294 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 294914 295634
rect 294294 259954 294914 295398
rect 294294 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 294914 259954
rect 294294 259634 294914 259718
rect 294294 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 294914 259634
rect 294294 223954 294914 259398
rect 294294 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 294914 223954
rect 294294 223634 294914 223718
rect 294294 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 294914 223634
rect 294294 187954 294914 223398
rect 294294 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 294914 187954
rect 294294 187634 294914 187718
rect 294294 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 294914 187634
rect 294294 151954 294914 187398
rect 294294 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 294914 151954
rect 294294 151634 294914 151718
rect 294294 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 294914 151634
rect 294294 115954 294914 151398
rect 294294 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 294914 115954
rect 294294 115634 294914 115718
rect 294294 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 294914 115634
rect 294294 79954 294914 115398
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 294294 43954 294914 79398
rect 294294 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 294914 43954
rect 294294 43634 294914 43718
rect 294294 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 294914 43634
rect 294294 7954 294914 43398
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1306 294914 7398
rect 294294 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 294914 -1306
rect 294294 -1626 294914 -1542
rect 294294 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 294914 -1626
rect 294294 -7654 294914 -1862
rect 298794 706758 299414 711590
rect 298794 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 299414 706758
rect 298794 706438 299414 706522
rect 298794 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 299414 706438
rect 298794 696454 299414 706202
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 660454 299414 695898
rect 298794 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 299414 660454
rect 298794 660134 299414 660218
rect 298794 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 299414 660134
rect 298794 624454 299414 659898
rect 298794 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 299414 624454
rect 298794 624134 299414 624218
rect 298794 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 299414 624134
rect 298794 588454 299414 623898
rect 298794 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 299414 588454
rect 298794 588134 299414 588218
rect 298794 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 299414 588134
rect 298794 552454 299414 587898
rect 298794 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 299414 552454
rect 298794 552134 299414 552218
rect 298794 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 299414 552134
rect 298794 516454 299414 551898
rect 298794 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 299414 516454
rect 298794 516134 299414 516218
rect 298794 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 299414 516134
rect 298794 480454 299414 515898
rect 298794 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 299414 480454
rect 298794 480134 299414 480218
rect 298794 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 299414 480134
rect 298794 444454 299414 479898
rect 298794 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 299414 444454
rect 298794 444134 299414 444218
rect 298794 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 299414 444134
rect 298794 408454 299414 443898
rect 298794 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 299414 408454
rect 298794 408134 299414 408218
rect 298794 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 299414 408134
rect 298794 372454 299414 407898
rect 298794 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 299414 372454
rect 298794 372134 299414 372218
rect 298794 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 299414 372134
rect 298794 336454 299414 371898
rect 298794 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 299414 336454
rect 298794 336134 299414 336218
rect 298794 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 299414 336134
rect 298794 300454 299414 335898
rect 298794 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 299414 300454
rect 298794 300134 299414 300218
rect 298794 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 299414 300134
rect 298794 264454 299414 299898
rect 298794 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 299414 264454
rect 298794 264134 299414 264218
rect 298794 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 299414 264134
rect 298794 228454 299414 263898
rect 298794 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 299414 228454
rect 298794 228134 299414 228218
rect 298794 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 299414 228134
rect 298794 192454 299414 227898
rect 298794 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 299414 192454
rect 298794 192134 299414 192218
rect 298794 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 299414 192134
rect 298794 156454 299414 191898
rect 298794 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 299414 156454
rect 298794 156134 299414 156218
rect 298794 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 299414 156134
rect 298794 120454 299414 155898
rect 298794 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 299414 120454
rect 298794 120134 299414 120218
rect 298794 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 299414 120134
rect 298794 84454 299414 119898
rect 298794 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 299414 84454
rect 298794 84134 299414 84218
rect 298794 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 299414 84134
rect 298794 48454 299414 83898
rect 298794 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 299414 48454
rect 298794 48134 299414 48218
rect 298794 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 299414 48134
rect 298794 12454 299414 47898
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298794 -2266 299414 11898
rect 298794 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 299414 -2266
rect 298794 -2586 299414 -2502
rect 298794 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 299414 -2586
rect 298794 -7654 299414 -2822
rect 303294 707718 303914 711590
rect 303294 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 303914 707718
rect 303294 707398 303914 707482
rect 303294 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 303914 707398
rect 303294 700954 303914 707162
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 664954 303914 700398
rect 303294 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 303914 664954
rect 303294 664634 303914 664718
rect 303294 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 303914 664634
rect 303294 628954 303914 664398
rect 303294 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 303914 628954
rect 303294 628634 303914 628718
rect 303294 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 303914 628634
rect 303294 592954 303914 628398
rect 303294 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 303914 592954
rect 303294 592634 303914 592718
rect 303294 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 303914 592634
rect 303294 556954 303914 592398
rect 303294 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 303914 556954
rect 303294 556634 303914 556718
rect 303294 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 303914 556634
rect 303294 520954 303914 556398
rect 303294 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 303914 520954
rect 303294 520634 303914 520718
rect 303294 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 303914 520634
rect 303294 484954 303914 520398
rect 303294 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 303914 484954
rect 303294 484634 303914 484718
rect 303294 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 303914 484634
rect 303294 448954 303914 484398
rect 303294 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 303914 448954
rect 303294 448634 303914 448718
rect 303294 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 303914 448634
rect 303294 412954 303914 448398
rect 303294 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 303914 412954
rect 303294 412634 303914 412718
rect 303294 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 303914 412634
rect 303294 376954 303914 412398
rect 303294 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 303914 376954
rect 303294 376634 303914 376718
rect 303294 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 303914 376634
rect 303294 340954 303914 376398
rect 303294 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 303914 340954
rect 303294 340634 303914 340718
rect 303294 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 303914 340634
rect 303294 304954 303914 340398
rect 303294 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 303914 304954
rect 303294 304634 303914 304718
rect 303294 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 303914 304634
rect 303294 268954 303914 304398
rect 303294 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 303914 268954
rect 303294 268634 303914 268718
rect 303294 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 303914 268634
rect 303294 232954 303914 268398
rect 303294 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 303914 232954
rect 303294 232634 303914 232718
rect 303294 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 303914 232634
rect 303294 196954 303914 232398
rect 303294 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 303914 196954
rect 303294 196634 303914 196718
rect 303294 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 303914 196634
rect 303294 160954 303914 196398
rect 303294 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 303914 160954
rect 303294 160634 303914 160718
rect 303294 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 303914 160634
rect 303294 124954 303914 160398
rect 303294 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 303914 124954
rect 303294 124634 303914 124718
rect 303294 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 303914 124634
rect 303294 88954 303914 124398
rect 303294 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 303914 88954
rect 303294 88634 303914 88718
rect 303294 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 303914 88634
rect 303294 52954 303914 88398
rect 303294 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 303914 52954
rect 303294 52634 303914 52718
rect 303294 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 303914 52634
rect 303294 16954 303914 52398
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 303294 -3226 303914 16398
rect 303294 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 303914 -3226
rect 303294 -3546 303914 -3462
rect 303294 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 303914 -3546
rect 303294 -7654 303914 -3782
rect 307794 708678 308414 711590
rect 307794 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 308414 708678
rect 307794 708358 308414 708442
rect 307794 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 308414 708358
rect 307794 669454 308414 708122
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4186 308414 20898
rect 307794 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 308414 -4186
rect 307794 -4506 308414 -4422
rect 307794 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 308414 -4506
rect 307794 -7654 308414 -4742
rect 312294 709638 312914 711590
rect 312294 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 312914 709638
rect 312294 709318 312914 709402
rect 312294 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 312914 709318
rect 312294 673954 312914 709082
rect 312294 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 312914 673954
rect 312294 673634 312914 673718
rect 312294 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 312914 673634
rect 312294 637954 312914 673398
rect 312294 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 312914 637954
rect 312294 637634 312914 637718
rect 312294 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 312914 637634
rect 312294 601954 312914 637398
rect 312294 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 312914 601954
rect 312294 601634 312914 601718
rect 312294 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 312914 601634
rect 312294 565954 312914 601398
rect 312294 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 312914 565954
rect 312294 565634 312914 565718
rect 312294 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 312914 565634
rect 312294 529954 312914 565398
rect 312294 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 312914 529954
rect 312294 529634 312914 529718
rect 312294 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 312914 529634
rect 312294 493954 312914 529398
rect 312294 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 312914 493954
rect 312294 493634 312914 493718
rect 312294 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 312914 493634
rect 312294 457954 312914 493398
rect 312294 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 312914 457954
rect 312294 457634 312914 457718
rect 312294 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 312914 457634
rect 312294 421954 312914 457398
rect 312294 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 312914 421954
rect 312294 421634 312914 421718
rect 312294 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 312914 421634
rect 312294 385954 312914 421398
rect 312294 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 312914 385954
rect 312294 385634 312914 385718
rect 312294 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 312914 385634
rect 312294 349954 312914 385398
rect 312294 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 312914 349954
rect 312294 349634 312914 349718
rect 312294 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 312914 349634
rect 312294 313954 312914 349398
rect 312294 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 312914 313954
rect 312294 313634 312914 313718
rect 312294 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 312914 313634
rect 312294 277954 312914 313398
rect 312294 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 312914 277954
rect 312294 277634 312914 277718
rect 312294 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 312914 277634
rect 312294 241954 312914 277398
rect 312294 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 312914 241954
rect 312294 241634 312914 241718
rect 312294 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 312914 241634
rect 312294 205954 312914 241398
rect 312294 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 312914 205954
rect 312294 205634 312914 205718
rect 312294 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 312914 205634
rect 312294 169954 312914 205398
rect 312294 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 312914 169954
rect 312294 169634 312914 169718
rect 312294 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 312914 169634
rect 312294 133954 312914 169398
rect 312294 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 312914 133954
rect 312294 133634 312914 133718
rect 312294 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 312914 133634
rect 312294 97954 312914 133398
rect 312294 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 312914 97954
rect 312294 97634 312914 97718
rect 312294 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 312914 97634
rect 312294 61954 312914 97398
rect 312294 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 312914 61954
rect 312294 61634 312914 61718
rect 312294 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 312914 61634
rect 312294 25954 312914 61398
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 312294 -5146 312914 25398
rect 312294 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 312914 -5146
rect 312294 -5466 312914 -5382
rect 312294 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 312914 -5466
rect 312294 -7654 312914 -5702
rect 316794 710598 317414 711590
rect 316794 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 317414 710598
rect 316794 710278 317414 710362
rect 316794 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 317414 710278
rect 316794 678454 317414 710042
rect 316794 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 317414 678454
rect 316794 678134 317414 678218
rect 316794 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 317414 678134
rect 316794 642454 317414 677898
rect 316794 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 317414 642454
rect 316794 642134 317414 642218
rect 316794 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 317414 642134
rect 316794 606454 317414 641898
rect 316794 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 317414 606454
rect 316794 606134 317414 606218
rect 316794 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 317414 606134
rect 316794 570454 317414 605898
rect 316794 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 317414 570454
rect 316794 570134 317414 570218
rect 316794 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 317414 570134
rect 316794 534454 317414 569898
rect 316794 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 317414 534454
rect 316794 534134 317414 534218
rect 316794 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 317414 534134
rect 316794 498454 317414 533898
rect 316794 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 317414 498454
rect 316794 498134 317414 498218
rect 316794 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 317414 498134
rect 316794 462454 317414 497898
rect 316794 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 317414 462454
rect 316794 462134 317414 462218
rect 316794 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 317414 462134
rect 316794 426454 317414 461898
rect 316794 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 317414 426454
rect 316794 426134 317414 426218
rect 316794 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 317414 426134
rect 316794 390454 317414 425898
rect 316794 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 317414 390454
rect 316794 390134 317414 390218
rect 316794 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 317414 390134
rect 316794 354454 317414 389898
rect 316794 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 317414 354454
rect 316794 354134 317414 354218
rect 316794 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 317414 354134
rect 316794 318454 317414 353898
rect 316794 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 317414 318454
rect 316794 318134 317414 318218
rect 316794 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 317414 318134
rect 316794 282454 317414 317898
rect 316794 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 317414 282454
rect 316794 282134 317414 282218
rect 316794 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 317414 282134
rect 316794 246454 317414 281898
rect 316794 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 317414 246454
rect 316794 246134 317414 246218
rect 316794 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 317414 246134
rect 316794 210454 317414 245898
rect 316794 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 317414 210454
rect 316794 210134 317414 210218
rect 316794 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 317414 210134
rect 316794 174454 317414 209898
rect 316794 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 317414 174454
rect 316794 174134 317414 174218
rect 316794 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 317414 174134
rect 316794 138454 317414 173898
rect 316794 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 317414 138454
rect 316794 138134 317414 138218
rect 316794 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 317414 138134
rect 316794 102454 317414 137898
rect 316794 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 317414 102454
rect 316794 102134 317414 102218
rect 316794 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 317414 102134
rect 316794 66454 317414 101898
rect 316794 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 317414 66454
rect 316794 66134 317414 66218
rect 316794 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 317414 66134
rect 316794 30454 317414 65898
rect 316794 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 317414 30454
rect 316794 30134 317414 30218
rect 316794 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 317414 30134
rect 316794 -6106 317414 29898
rect 316794 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 317414 -6106
rect 316794 -6426 317414 -6342
rect 316794 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 317414 -6426
rect 316794 -7654 317414 -6662
rect 321294 711558 321914 711590
rect 321294 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 321914 711558
rect 321294 711238 321914 711322
rect 321294 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 321914 711238
rect 321294 682954 321914 711002
rect 321294 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 321914 682954
rect 321294 682634 321914 682718
rect 321294 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 321914 682634
rect 321294 646954 321914 682398
rect 321294 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 321914 646954
rect 321294 646634 321914 646718
rect 321294 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 321914 646634
rect 321294 610954 321914 646398
rect 321294 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 321914 610954
rect 321294 610634 321914 610718
rect 321294 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 321914 610634
rect 321294 574954 321914 610398
rect 321294 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 321914 574954
rect 321294 574634 321914 574718
rect 321294 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 321914 574634
rect 321294 538954 321914 574398
rect 321294 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 321914 538954
rect 321294 538634 321914 538718
rect 321294 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 321914 538634
rect 321294 502954 321914 538398
rect 321294 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 321914 502954
rect 321294 502634 321914 502718
rect 321294 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 321914 502634
rect 321294 466954 321914 502398
rect 321294 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 321914 466954
rect 321294 466634 321914 466718
rect 321294 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 321914 466634
rect 321294 430954 321914 466398
rect 321294 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 321914 430954
rect 321294 430634 321914 430718
rect 321294 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 321914 430634
rect 321294 394954 321914 430398
rect 321294 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 321914 394954
rect 321294 394634 321914 394718
rect 321294 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 321914 394634
rect 321294 358954 321914 394398
rect 321294 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 321914 358954
rect 321294 358634 321914 358718
rect 321294 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 321914 358634
rect 321294 322954 321914 358398
rect 321294 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 321914 322954
rect 321294 322634 321914 322718
rect 321294 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 321914 322634
rect 321294 286954 321914 322398
rect 321294 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 321914 286954
rect 321294 286634 321914 286718
rect 321294 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 321914 286634
rect 321294 250954 321914 286398
rect 321294 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 321914 250954
rect 321294 250634 321914 250718
rect 321294 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 321914 250634
rect 321294 214954 321914 250398
rect 321294 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 321914 214954
rect 321294 214634 321914 214718
rect 321294 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 321914 214634
rect 321294 178954 321914 214398
rect 321294 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 321914 178954
rect 321294 178634 321914 178718
rect 321294 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 321914 178634
rect 321294 142954 321914 178398
rect 321294 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 321914 142954
rect 321294 142634 321914 142718
rect 321294 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 321914 142634
rect 321294 106954 321914 142398
rect 321294 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 321914 106954
rect 321294 106634 321914 106718
rect 321294 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 321914 106634
rect 321294 70954 321914 106398
rect 321294 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 321914 70954
rect 321294 70634 321914 70718
rect 321294 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 321914 70634
rect 321294 34954 321914 70398
rect 321294 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 321914 34954
rect 321294 34634 321914 34718
rect 321294 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 321914 34634
rect 321294 -7066 321914 34398
rect 321294 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 321914 -7066
rect 321294 -7386 321914 -7302
rect 321294 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 321914 -7386
rect 321294 -7654 321914 -7622
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 330294 705798 330914 711590
rect 330294 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 330914 705798
rect 330294 705478 330914 705562
rect 330294 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 330914 705478
rect 330294 691954 330914 705242
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 655954 330914 691398
rect 330294 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 330914 655954
rect 330294 655634 330914 655718
rect 330294 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 330914 655634
rect 330294 619954 330914 655398
rect 330294 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 330914 619954
rect 330294 619634 330914 619718
rect 330294 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 330914 619634
rect 330294 583954 330914 619398
rect 330294 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 330914 583954
rect 330294 583634 330914 583718
rect 330294 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 330914 583634
rect 330294 547954 330914 583398
rect 330294 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 330914 547954
rect 330294 547634 330914 547718
rect 330294 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 330914 547634
rect 330294 511954 330914 547398
rect 330294 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 330914 511954
rect 330294 511634 330914 511718
rect 330294 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 330914 511634
rect 330294 475954 330914 511398
rect 330294 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 330914 475954
rect 330294 475634 330914 475718
rect 330294 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 330914 475634
rect 330294 439954 330914 475398
rect 330294 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 330914 439954
rect 330294 439634 330914 439718
rect 330294 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 330914 439634
rect 330294 403954 330914 439398
rect 330294 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 330914 403954
rect 330294 403634 330914 403718
rect 330294 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 330914 403634
rect 330294 367954 330914 403398
rect 330294 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 330914 367954
rect 330294 367634 330914 367718
rect 330294 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 330914 367634
rect 330294 331954 330914 367398
rect 330294 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 330914 331954
rect 330294 331634 330914 331718
rect 330294 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 330914 331634
rect 330294 295954 330914 331398
rect 330294 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 330914 295954
rect 330294 295634 330914 295718
rect 330294 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 330914 295634
rect 330294 259954 330914 295398
rect 330294 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 330914 259954
rect 330294 259634 330914 259718
rect 330294 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 330914 259634
rect 330294 223954 330914 259398
rect 330294 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 330914 223954
rect 330294 223634 330914 223718
rect 330294 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 330914 223634
rect 330294 187954 330914 223398
rect 330294 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 330914 187954
rect 330294 187634 330914 187718
rect 330294 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 330914 187634
rect 330294 151954 330914 187398
rect 330294 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 330914 151954
rect 330294 151634 330914 151718
rect 330294 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 330914 151634
rect 330294 115954 330914 151398
rect 330294 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 330914 115954
rect 330294 115634 330914 115718
rect 330294 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 330914 115634
rect 330294 79954 330914 115398
rect 330294 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 330914 79954
rect 330294 79634 330914 79718
rect 330294 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 330914 79634
rect 330294 43954 330914 79398
rect 330294 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 330914 43954
rect 330294 43634 330914 43718
rect 330294 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 330914 43634
rect 330294 7954 330914 43398
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1306 330914 7398
rect 330294 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 330914 -1306
rect 330294 -1626 330914 -1542
rect 330294 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 330914 -1626
rect 330294 -7654 330914 -1862
rect 334794 706758 335414 711590
rect 334794 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 335414 706758
rect 334794 706438 335414 706522
rect 334794 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 335414 706438
rect 334794 696454 335414 706202
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 660454 335414 695898
rect 334794 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 335414 660454
rect 334794 660134 335414 660218
rect 334794 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 335414 660134
rect 334794 624454 335414 659898
rect 334794 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 335414 624454
rect 334794 624134 335414 624218
rect 334794 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 335414 624134
rect 334794 588454 335414 623898
rect 334794 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 335414 588454
rect 334794 588134 335414 588218
rect 334794 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 335414 588134
rect 334794 552454 335414 587898
rect 334794 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 335414 552454
rect 334794 552134 335414 552218
rect 334794 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 335414 552134
rect 334794 516454 335414 551898
rect 334794 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 335414 516454
rect 334794 516134 335414 516218
rect 334794 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 335414 516134
rect 334794 480454 335414 515898
rect 334794 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 335414 480454
rect 334794 480134 335414 480218
rect 334794 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 335414 480134
rect 334794 444454 335414 479898
rect 334794 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 335414 444454
rect 334794 444134 335414 444218
rect 334794 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 335414 444134
rect 334794 408454 335414 443898
rect 334794 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 335414 408454
rect 334794 408134 335414 408218
rect 334794 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 335414 408134
rect 334794 372454 335414 407898
rect 334794 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 335414 372454
rect 334794 372134 335414 372218
rect 334794 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 335414 372134
rect 334794 336454 335414 371898
rect 334794 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 335414 336454
rect 334794 336134 335414 336218
rect 334794 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 335414 336134
rect 334794 300454 335414 335898
rect 334794 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 335414 300454
rect 334794 300134 335414 300218
rect 334794 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 335414 300134
rect 334794 264454 335414 299898
rect 334794 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 335414 264454
rect 334794 264134 335414 264218
rect 334794 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 335414 264134
rect 334794 228454 335414 263898
rect 334794 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 335414 228454
rect 334794 228134 335414 228218
rect 334794 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 335414 228134
rect 334794 192454 335414 227898
rect 334794 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 335414 192454
rect 334794 192134 335414 192218
rect 334794 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 335414 192134
rect 334794 156454 335414 191898
rect 334794 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 335414 156454
rect 334794 156134 335414 156218
rect 334794 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 335414 156134
rect 334794 120454 335414 155898
rect 334794 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 335414 120454
rect 334794 120134 335414 120218
rect 334794 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 335414 120134
rect 334794 84454 335414 119898
rect 334794 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 335414 84454
rect 334794 84134 335414 84218
rect 334794 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 335414 84134
rect 334794 48454 335414 83898
rect 334794 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 335414 48454
rect 334794 48134 335414 48218
rect 334794 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 335414 48134
rect 334794 12454 335414 47898
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2266 335414 11898
rect 334794 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 335414 -2266
rect 334794 -2586 335414 -2502
rect 334794 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 335414 -2586
rect 334794 -7654 335414 -2822
rect 339294 707718 339914 711590
rect 339294 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 339914 707718
rect 339294 707398 339914 707482
rect 339294 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 339914 707398
rect 339294 700954 339914 707162
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 664954 339914 700398
rect 339294 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 339914 664954
rect 339294 664634 339914 664718
rect 339294 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 339914 664634
rect 339294 628954 339914 664398
rect 339294 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 339914 628954
rect 339294 628634 339914 628718
rect 339294 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 339914 628634
rect 339294 592954 339914 628398
rect 339294 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 339914 592954
rect 339294 592634 339914 592718
rect 339294 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 339914 592634
rect 339294 556954 339914 592398
rect 339294 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 339914 556954
rect 339294 556634 339914 556718
rect 339294 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 339914 556634
rect 339294 520954 339914 556398
rect 339294 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 339914 520954
rect 339294 520634 339914 520718
rect 339294 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 339914 520634
rect 339294 484954 339914 520398
rect 339294 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 339914 484954
rect 339294 484634 339914 484718
rect 339294 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 339914 484634
rect 339294 448954 339914 484398
rect 339294 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 339914 448954
rect 339294 448634 339914 448718
rect 339294 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 339914 448634
rect 339294 412954 339914 448398
rect 339294 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 339914 412954
rect 339294 412634 339914 412718
rect 339294 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 339914 412634
rect 339294 376954 339914 412398
rect 339294 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 339914 376954
rect 339294 376634 339914 376718
rect 339294 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 339914 376634
rect 339294 340954 339914 376398
rect 339294 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 339914 340954
rect 339294 340634 339914 340718
rect 339294 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 339914 340634
rect 339294 304954 339914 340398
rect 339294 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 339914 304954
rect 339294 304634 339914 304718
rect 339294 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 339914 304634
rect 339294 268954 339914 304398
rect 339294 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 339914 268954
rect 339294 268634 339914 268718
rect 339294 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 339914 268634
rect 339294 232954 339914 268398
rect 339294 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 339914 232954
rect 339294 232634 339914 232718
rect 339294 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 339914 232634
rect 339294 196954 339914 232398
rect 339294 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 339914 196954
rect 339294 196634 339914 196718
rect 339294 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 339914 196634
rect 339294 160954 339914 196398
rect 339294 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 339914 160954
rect 339294 160634 339914 160718
rect 339294 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 339914 160634
rect 339294 124954 339914 160398
rect 339294 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 339914 124954
rect 339294 124634 339914 124718
rect 339294 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 339914 124634
rect 339294 88954 339914 124398
rect 339294 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 339914 88954
rect 339294 88634 339914 88718
rect 339294 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 339914 88634
rect 339294 52954 339914 88398
rect 339294 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 339914 52954
rect 339294 52634 339914 52718
rect 339294 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 339914 52634
rect 339294 16954 339914 52398
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3226 339914 16398
rect 339294 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 339914 -3226
rect 339294 -3546 339914 -3462
rect 339294 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 339914 -3546
rect 339294 -7654 339914 -3782
rect 343794 708678 344414 711590
rect 343794 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 344414 708678
rect 343794 708358 344414 708442
rect 343794 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 344414 708358
rect 343794 669454 344414 708122
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -4186 344414 20898
rect 343794 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 344414 -4186
rect 343794 -4506 344414 -4422
rect 343794 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 344414 -4506
rect 343794 -7654 344414 -4742
rect 348294 709638 348914 711590
rect 348294 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 348914 709638
rect 348294 709318 348914 709402
rect 348294 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 348914 709318
rect 348294 673954 348914 709082
rect 348294 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 348914 673954
rect 348294 673634 348914 673718
rect 348294 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 348914 673634
rect 348294 637954 348914 673398
rect 348294 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 348914 637954
rect 348294 637634 348914 637718
rect 348294 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 348914 637634
rect 348294 601954 348914 637398
rect 348294 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 348914 601954
rect 348294 601634 348914 601718
rect 348294 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 348914 601634
rect 348294 565954 348914 601398
rect 348294 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 348914 565954
rect 348294 565634 348914 565718
rect 348294 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 348914 565634
rect 348294 529954 348914 565398
rect 348294 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 348914 529954
rect 348294 529634 348914 529718
rect 348294 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 348914 529634
rect 348294 493954 348914 529398
rect 348294 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 348914 493954
rect 348294 493634 348914 493718
rect 348294 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 348914 493634
rect 348294 457954 348914 493398
rect 348294 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 348914 457954
rect 348294 457634 348914 457718
rect 348294 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 348914 457634
rect 348294 421954 348914 457398
rect 348294 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 348914 421954
rect 348294 421634 348914 421718
rect 348294 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 348914 421634
rect 348294 385954 348914 421398
rect 348294 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 348914 385954
rect 348294 385634 348914 385718
rect 348294 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 348914 385634
rect 348294 349954 348914 385398
rect 348294 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 348914 349954
rect 348294 349634 348914 349718
rect 348294 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 348914 349634
rect 348294 313954 348914 349398
rect 348294 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 348914 313954
rect 348294 313634 348914 313718
rect 348294 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 348914 313634
rect 348294 277954 348914 313398
rect 348294 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 348914 277954
rect 348294 277634 348914 277718
rect 348294 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 348914 277634
rect 348294 241954 348914 277398
rect 348294 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 348914 241954
rect 348294 241634 348914 241718
rect 348294 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 348914 241634
rect 348294 205954 348914 241398
rect 348294 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 348914 205954
rect 348294 205634 348914 205718
rect 348294 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 348914 205634
rect 348294 169954 348914 205398
rect 348294 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 348914 169954
rect 348294 169634 348914 169718
rect 348294 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 348914 169634
rect 348294 133954 348914 169398
rect 348294 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 348914 133954
rect 348294 133634 348914 133718
rect 348294 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 348914 133634
rect 348294 97954 348914 133398
rect 348294 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 348914 97954
rect 348294 97634 348914 97718
rect 348294 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 348914 97634
rect 348294 61954 348914 97398
rect 348294 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 348914 61954
rect 348294 61634 348914 61718
rect 348294 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 348914 61634
rect 348294 25954 348914 61398
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 348294 -5146 348914 25398
rect 348294 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 348914 -5146
rect 348294 -5466 348914 -5382
rect 348294 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 348914 -5466
rect 348294 -7654 348914 -5702
rect 352794 710598 353414 711590
rect 352794 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 353414 710598
rect 352794 710278 353414 710362
rect 352794 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 353414 710278
rect 352794 678454 353414 710042
rect 352794 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 353414 678454
rect 352794 678134 353414 678218
rect 352794 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 353414 678134
rect 352794 642454 353414 677898
rect 352794 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 353414 642454
rect 352794 642134 353414 642218
rect 352794 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 353414 642134
rect 352794 606454 353414 641898
rect 352794 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 353414 606454
rect 352794 606134 353414 606218
rect 352794 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 353414 606134
rect 352794 570454 353414 605898
rect 352794 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 353414 570454
rect 352794 570134 353414 570218
rect 352794 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 353414 570134
rect 352794 534454 353414 569898
rect 352794 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 353414 534454
rect 352794 534134 353414 534218
rect 352794 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 353414 534134
rect 352794 498454 353414 533898
rect 352794 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 353414 498454
rect 352794 498134 353414 498218
rect 352794 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 353414 498134
rect 352794 462454 353414 497898
rect 352794 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 353414 462454
rect 352794 462134 353414 462218
rect 352794 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 353414 462134
rect 352794 426454 353414 461898
rect 352794 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 353414 426454
rect 352794 426134 353414 426218
rect 352794 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 353414 426134
rect 352794 390454 353414 425898
rect 352794 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 353414 390454
rect 352794 390134 353414 390218
rect 352794 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 353414 390134
rect 352794 354454 353414 389898
rect 352794 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 353414 354454
rect 352794 354134 353414 354218
rect 352794 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 353414 354134
rect 352794 318454 353414 353898
rect 352794 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 353414 318454
rect 352794 318134 353414 318218
rect 352794 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 353414 318134
rect 352794 282454 353414 317898
rect 352794 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 353414 282454
rect 352794 282134 353414 282218
rect 352794 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 353414 282134
rect 352794 246454 353414 281898
rect 352794 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 353414 246454
rect 352794 246134 353414 246218
rect 352794 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 353414 246134
rect 352794 210454 353414 245898
rect 352794 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 353414 210454
rect 352794 210134 353414 210218
rect 352794 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 353414 210134
rect 352794 174454 353414 209898
rect 352794 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 353414 174454
rect 352794 174134 353414 174218
rect 352794 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 353414 174134
rect 352794 138454 353414 173898
rect 352794 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 353414 138454
rect 352794 138134 353414 138218
rect 352794 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 353414 138134
rect 352794 102454 353414 137898
rect 352794 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 353414 102454
rect 352794 102134 353414 102218
rect 352794 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 353414 102134
rect 352794 66454 353414 101898
rect 352794 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 353414 66454
rect 352794 66134 353414 66218
rect 352794 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 353414 66134
rect 352794 30454 353414 65898
rect 352794 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 353414 30454
rect 352794 30134 353414 30218
rect 352794 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 353414 30134
rect 352794 -6106 353414 29898
rect 352794 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 353414 -6106
rect 352794 -6426 353414 -6342
rect 352794 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 353414 -6426
rect 352794 -7654 353414 -6662
rect 357294 711558 357914 711590
rect 357294 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 357914 711558
rect 357294 711238 357914 711322
rect 357294 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 357914 711238
rect 357294 682954 357914 711002
rect 357294 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 357914 682954
rect 357294 682634 357914 682718
rect 357294 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 357914 682634
rect 357294 646954 357914 682398
rect 357294 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 357914 646954
rect 357294 646634 357914 646718
rect 357294 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 357914 646634
rect 357294 610954 357914 646398
rect 357294 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 357914 610954
rect 357294 610634 357914 610718
rect 357294 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 357914 610634
rect 357294 574954 357914 610398
rect 357294 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 357914 574954
rect 357294 574634 357914 574718
rect 357294 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 357914 574634
rect 357294 538954 357914 574398
rect 357294 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 357914 538954
rect 357294 538634 357914 538718
rect 357294 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 357914 538634
rect 357294 502954 357914 538398
rect 357294 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 357914 502954
rect 357294 502634 357914 502718
rect 357294 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 357914 502634
rect 357294 466954 357914 502398
rect 357294 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 357914 466954
rect 357294 466634 357914 466718
rect 357294 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 357914 466634
rect 357294 430954 357914 466398
rect 357294 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 357914 430954
rect 357294 430634 357914 430718
rect 357294 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 357914 430634
rect 357294 394954 357914 430398
rect 357294 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 357914 394954
rect 357294 394634 357914 394718
rect 357294 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 357914 394634
rect 357294 358954 357914 394398
rect 357294 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 357914 358954
rect 357294 358634 357914 358718
rect 357294 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 357914 358634
rect 357294 322954 357914 358398
rect 357294 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 357914 322954
rect 357294 322634 357914 322718
rect 357294 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 357914 322634
rect 357294 286954 357914 322398
rect 357294 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 357914 286954
rect 357294 286634 357914 286718
rect 357294 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 357914 286634
rect 357294 250954 357914 286398
rect 357294 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 357914 250954
rect 357294 250634 357914 250718
rect 357294 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 357914 250634
rect 357294 214954 357914 250398
rect 357294 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 357914 214954
rect 357294 214634 357914 214718
rect 357294 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 357914 214634
rect 357294 178954 357914 214398
rect 357294 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 357914 178954
rect 357294 178634 357914 178718
rect 357294 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 357914 178634
rect 357294 142954 357914 178398
rect 357294 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 357914 142954
rect 357294 142634 357914 142718
rect 357294 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 357914 142634
rect 357294 106954 357914 142398
rect 357294 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 357914 106954
rect 357294 106634 357914 106718
rect 357294 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 357914 106634
rect 357294 70954 357914 106398
rect 357294 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 357914 70954
rect 357294 70634 357914 70718
rect 357294 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 357914 70634
rect 357294 34954 357914 70398
rect 357294 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 357914 34954
rect 357294 34634 357914 34718
rect 357294 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 357914 34634
rect 357294 -7066 357914 34398
rect 357294 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 357914 -7066
rect 357294 -7386 357914 -7302
rect 357294 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 357914 -7386
rect 357294 -7654 357914 -7622
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 366294 705798 366914 711590
rect 366294 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 366914 705798
rect 366294 705478 366914 705562
rect 366294 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 366914 705478
rect 366294 691954 366914 705242
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 655954 366914 691398
rect 366294 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 366914 655954
rect 366294 655634 366914 655718
rect 366294 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 366914 655634
rect 366294 619954 366914 655398
rect 366294 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 366914 619954
rect 366294 619634 366914 619718
rect 366294 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 366914 619634
rect 366294 583954 366914 619398
rect 366294 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 366914 583954
rect 366294 583634 366914 583718
rect 366294 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 366914 583634
rect 366294 547954 366914 583398
rect 366294 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 366914 547954
rect 366294 547634 366914 547718
rect 366294 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 366914 547634
rect 366294 511954 366914 547398
rect 366294 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 366914 511954
rect 366294 511634 366914 511718
rect 366294 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 366914 511634
rect 366294 475954 366914 511398
rect 366294 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 366914 475954
rect 366294 475634 366914 475718
rect 366294 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 366914 475634
rect 366294 439954 366914 475398
rect 366294 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 366914 439954
rect 366294 439634 366914 439718
rect 366294 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 366914 439634
rect 366294 403954 366914 439398
rect 366294 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 366914 403954
rect 366294 403634 366914 403718
rect 366294 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 366914 403634
rect 366294 367954 366914 403398
rect 366294 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 366914 367954
rect 366294 367634 366914 367718
rect 366294 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 366914 367634
rect 366294 331954 366914 367398
rect 366294 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 366914 331954
rect 366294 331634 366914 331718
rect 366294 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 366914 331634
rect 366294 295954 366914 331398
rect 366294 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 366914 295954
rect 366294 295634 366914 295718
rect 366294 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 366914 295634
rect 366294 259954 366914 295398
rect 366294 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 366914 259954
rect 366294 259634 366914 259718
rect 366294 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 366914 259634
rect 366294 223954 366914 259398
rect 366294 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 366914 223954
rect 366294 223634 366914 223718
rect 366294 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 366914 223634
rect 366294 187954 366914 223398
rect 366294 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 366914 187954
rect 366294 187634 366914 187718
rect 366294 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 366914 187634
rect 366294 151954 366914 187398
rect 366294 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 366914 151954
rect 366294 151634 366914 151718
rect 366294 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 366914 151634
rect 366294 115954 366914 151398
rect 366294 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 366914 115954
rect 366294 115634 366914 115718
rect 366294 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 366914 115634
rect 366294 79954 366914 115398
rect 366294 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 366914 79954
rect 366294 79634 366914 79718
rect 366294 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 366914 79634
rect 366294 43954 366914 79398
rect 366294 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 366914 43954
rect 366294 43634 366914 43718
rect 366294 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 366914 43634
rect 366294 7954 366914 43398
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 366294 -1306 366914 7398
rect 366294 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 366914 -1306
rect 366294 -1626 366914 -1542
rect 366294 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 366914 -1626
rect 366294 -7654 366914 -1862
rect 370794 706758 371414 711590
rect 370794 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 371414 706758
rect 370794 706438 371414 706522
rect 370794 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 371414 706438
rect 370794 696454 371414 706202
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 660454 371414 695898
rect 370794 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 371414 660454
rect 370794 660134 371414 660218
rect 370794 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 371414 660134
rect 370794 624454 371414 659898
rect 370794 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 371414 624454
rect 370794 624134 371414 624218
rect 370794 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 371414 624134
rect 370794 588454 371414 623898
rect 370794 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 371414 588454
rect 370794 588134 371414 588218
rect 370794 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 371414 588134
rect 370794 552454 371414 587898
rect 370794 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 371414 552454
rect 370794 552134 371414 552218
rect 370794 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 371414 552134
rect 370794 516454 371414 551898
rect 370794 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 371414 516454
rect 370794 516134 371414 516218
rect 370794 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 371414 516134
rect 370794 480454 371414 515898
rect 370794 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 371414 480454
rect 370794 480134 371414 480218
rect 370794 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 371414 480134
rect 370794 444454 371414 479898
rect 370794 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 371414 444454
rect 370794 444134 371414 444218
rect 370794 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 371414 444134
rect 370794 408454 371414 443898
rect 370794 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 371414 408454
rect 370794 408134 371414 408218
rect 370794 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 371414 408134
rect 370794 372454 371414 407898
rect 370794 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 371414 372454
rect 370794 372134 371414 372218
rect 370794 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 371414 372134
rect 370794 336454 371414 371898
rect 370794 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 371414 336454
rect 370794 336134 371414 336218
rect 370794 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 371414 336134
rect 370794 300454 371414 335898
rect 370794 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 371414 300454
rect 370794 300134 371414 300218
rect 370794 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 371414 300134
rect 370794 264454 371414 299898
rect 370794 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 371414 264454
rect 370794 264134 371414 264218
rect 370794 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 371414 264134
rect 370794 228454 371414 263898
rect 370794 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 371414 228454
rect 370794 228134 371414 228218
rect 370794 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 371414 228134
rect 370794 192454 371414 227898
rect 370794 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 371414 192454
rect 370794 192134 371414 192218
rect 370794 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 371414 192134
rect 370794 156454 371414 191898
rect 370794 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 371414 156454
rect 370794 156134 371414 156218
rect 370794 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 371414 156134
rect 370794 120454 371414 155898
rect 370794 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 371414 120454
rect 370794 120134 371414 120218
rect 370794 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 371414 120134
rect 370794 84454 371414 119898
rect 370794 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 371414 84454
rect 370794 84134 371414 84218
rect 370794 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 371414 84134
rect 370794 48454 371414 83898
rect 370794 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 371414 48454
rect 370794 48134 371414 48218
rect 370794 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 371414 48134
rect 370794 12454 371414 47898
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -2266 371414 11898
rect 370794 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 371414 -2266
rect 370794 -2586 371414 -2502
rect 370794 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 371414 -2586
rect 370794 -7654 371414 -2822
rect 375294 707718 375914 711590
rect 375294 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 375914 707718
rect 375294 707398 375914 707482
rect 375294 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 375914 707398
rect 375294 700954 375914 707162
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 664954 375914 700398
rect 375294 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 375914 664954
rect 375294 664634 375914 664718
rect 375294 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 375914 664634
rect 375294 628954 375914 664398
rect 375294 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 375914 628954
rect 375294 628634 375914 628718
rect 375294 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 375914 628634
rect 375294 592954 375914 628398
rect 375294 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 375914 592954
rect 375294 592634 375914 592718
rect 375294 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 375914 592634
rect 375294 556954 375914 592398
rect 375294 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 375914 556954
rect 375294 556634 375914 556718
rect 375294 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 375914 556634
rect 375294 520954 375914 556398
rect 375294 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 375914 520954
rect 375294 520634 375914 520718
rect 375294 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 375914 520634
rect 375294 484954 375914 520398
rect 375294 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 375914 484954
rect 375294 484634 375914 484718
rect 375294 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 375914 484634
rect 375294 448954 375914 484398
rect 375294 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 375914 448954
rect 375294 448634 375914 448718
rect 375294 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 375914 448634
rect 375294 412954 375914 448398
rect 375294 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 375914 412954
rect 375294 412634 375914 412718
rect 375294 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 375914 412634
rect 375294 376954 375914 412398
rect 375294 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 375914 376954
rect 375294 376634 375914 376718
rect 375294 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 375914 376634
rect 375294 340954 375914 376398
rect 375294 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 375914 340954
rect 375294 340634 375914 340718
rect 375294 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 375914 340634
rect 375294 304954 375914 340398
rect 375294 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 375914 304954
rect 375294 304634 375914 304718
rect 375294 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 375914 304634
rect 375294 268954 375914 304398
rect 375294 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 375914 268954
rect 375294 268634 375914 268718
rect 375294 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 375914 268634
rect 375294 232954 375914 268398
rect 375294 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 375914 232954
rect 375294 232634 375914 232718
rect 375294 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 375914 232634
rect 375294 196954 375914 232398
rect 375294 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 375914 196954
rect 375294 196634 375914 196718
rect 375294 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 375914 196634
rect 375294 160954 375914 196398
rect 375294 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 375914 160954
rect 375294 160634 375914 160718
rect 375294 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 375914 160634
rect 375294 124954 375914 160398
rect 375294 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 375914 124954
rect 375294 124634 375914 124718
rect 375294 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 375914 124634
rect 375294 88954 375914 124398
rect 375294 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 375914 88954
rect 375294 88634 375914 88718
rect 375294 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 375914 88634
rect 375294 52954 375914 88398
rect 375294 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 375914 52954
rect 375294 52634 375914 52718
rect 375294 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 375914 52634
rect 375294 16954 375914 52398
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3226 375914 16398
rect 375294 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 375914 -3226
rect 375294 -3546 375914 -3462
rect 375294 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 375914 -3546
rect 375294 -7654 375914 -3782
rect 379794 708678 380414 711590
rect 379794 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 380414 708678
rect 379794 708358 380414 708442
rect 379794 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 380414 708358
rect 379794 669454 380414 708122
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4186 380414 20898
rect 379794 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 380414 -4186
rect 379794 -4506 380414 -4422
rect 379794 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 380414 -4506
rect 379794 -7654 380414 -4742
rect 384294 709638 384914 711590
rect 384294 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 384914 709638
rect 384294 709318 384914 709402
rect 384294 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 384914 709318
rect 384294 673954 384914 709082
rect 384294 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 384914 673954
rect 384294 673634 384914 673718
rect 384294 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 384914 673634
rect 384294 637954 384914 673398
rect 384294 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 384914 637954
rect 384294 637634 384914 637718
rect 384294 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 384914 637634
rect 384294 601954 384914 637398
rect 384294 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 384914 601954
rect 384294 601634 384914 601718
rect 384294 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 384914 601634
rect 384294 565954 384914 601398
rect 384294 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 384914 565954
rect 384294 565634 384914 565718
rect 384294 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 384914 565634
rect 384294 529954 384914 565398
rect 384294 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 384914 529954
rect 384294 529634 384914 529718
rect 384294 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 384914 529634
rect 384294 493954 384914 529398
rect 384294 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 384914 493954
rect 384294 493634 384914 493718
rect 384294 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 384914 493634
rect 384294 457954 384914 493398
rect 384294 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 384914 457954
rect 384294 457634 384914 457718
rect 384294 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 384914 457634
rect 384294 421954 384914 457398
rect 384294 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 384914 421954
rect 384294 421634 384914 421718
rect 384294 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 384914 421634
rect 384294 385954 384914 421398
rect 384294 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 384914 385954
rect 384294 385634 384914 385718
rect 384294 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 384914 385634
rect 384294 349954 384914 385398
rect 384294 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 384914 349954
rect 384294 349634 384914 349718
rect 384294 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 384914 349634
rect 384294 313954 384914 349398
rect 384294 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 384914 313954
rect 384294 313634 384914 313718
rect 384294 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 384914 313634
rect 384294 277954 384914 313398
rect 384294 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 384914 277954
rect 384294 277634 384914 277718
rect 384294 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 384914 277634
rect 384294 241954 384914 277398
rect 384294 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 384914 241954
rect 384294 241634 384914 241718
rect 384294 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 384914 241634
rect 384294 205954 384914 241398
rect 384294 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 384914 205954
rect 384294 205634 384914 205718
rect 384294 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 384914 205634
rect 384294 169954 384914 205398
rect 384294 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 384914 169954
rect 384294 169634 384914 169718
rect 384294 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 384914 169634
rect 384294 133954 384914 169398
rect 384294 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 384914 133954
rect 384294 133634 384914 133718
rect 384294 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 384914 133634
rect 384294 97954 384914 133398
rect 384294 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 384914 97954
rect 384294 97634 384914 97718
rect 384294 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 384914 97634
rect 384294 61954 384914 97398
rect 384294 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 384914 61954
rect 384294 61634 384914 61718
rect 384294 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 384914 61634
rect 384294 25954 384914 61398
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5146 384914 25398
rect 384294 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 384914 -5146
rect 384294 -5466 384914 -5382
rect 384294 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 384914 -5466
rect 384294 -7654 384914 -5702
rect 388794 710598 389414 711590
rect 388794 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 389414 710598
rect 388794 710278 389414 710362
rect 388794 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 389414 710278
rect 388794 678454 389414 710042
rect 388794 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 389414 678454
rect 388794 678134 389414 678218
rect 388794 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 389414 678134
rect 388794 642454 389414 677898
rect 388794 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 389414 642454
rect 388794 642134 389414 642218
rect 388794 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 389414 642134
rect 388794 606454 389414 641898
rect 388794 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 389414 606454
rect 388794 606134 389414 606218
rect 388794 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 389414 606134
rect 388794 570454 389414 605898
rect 388794 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 389414 570454
rect 388794 570134 389414 570218
rect 388794 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 389414 570134
rect 388794 534454 389414 569898
rect 388794 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 389414 534454
rect 388794 534134 389414 534218
rect 388794 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 389414 534134
rect 388794 498454 389414 533898
rect 388794 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 389414 498454
rect 388794 498134 389414 498218
rect 388794 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 389414 498134
rect 388794 462454 389414 497898
rect 388794 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 389414 462454
rect 388794 462134 389414 462218
rect 388794 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 389414 462134
rect 388794 426454 389414 461898
rect 388794 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 389414 426454
rect 388794 426134 389414 426218
rect 388794 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 389414 426134
rect 388794 390454 389414 425898
rect 388794 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 389414 390454
rect 388794 390134 389414 390218
rect 388794 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 389414 390134
rect 388794 354454 389414 389898
rect 388794 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 389414 354454
rect 388794 354134 389414 354218
rect 388794 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 389414 354134
rect 388794 318454 389414 353898
rect 388794 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 389414 318454
rect 388794 318134 389414 318218
rect 388794 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 389414 318134
rect 388794 282454 389414 317898
rect 388794 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 389414 282454
rect 388794 282134 389414 282218
rect 388794 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 389414 282134
rect 388794 246454 389414 281898
rect 388794 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 389414 246454
rect 388794 246134 389414 246218
rect 388794 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 389414 246134
rect 388794 210454 389414 245898
rect 388794 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 389414 210454
rect 388794 210134 389414 210218
rect 388794 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 389414 210134
rect 388794 174454 389414 209898
rect 388794 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 389414 174454
rect 388794 174134 389414 174218
rect 388794 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 389414 174134
rect 388794 138454 389414 173898
rect 388794 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 389414 138454
rect 388794 138134 389414 138218
rect 388794 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 389414 138134
rect 388794 102454 389414 137898
rect 388794 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 389414 102454
rect 388794 102134 389414 102218
rect 388794 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 389414 102134
rect 388794 66454 389414 101898
rect 388794 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 389414 66454
rect 388794 66134 389414 66218
rect 388794 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 389414 66134
rect 388794 30454 389414 65898
rect 388794 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 389414 30454
rect 388794 30134 389414 30218
rect 388794 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 389414 30134
rect 388794 -6106 389414 29898
rect 388794 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 389414 -6106
rect 388794 -6426 389414 -6342
rect 388794 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 389414 -6426
rect 388794 -7654 389414 -6662
rect 393294 711558 393914 711590
rect 393294 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 393914 711558
rect 393294 711238 393914 711322
rect 393294 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 393914 711238
rect 393294 682954 393914 711002
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 393294 646954 393914 682398
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 393294 610954 393914 646398
rect 393294 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 393914 610954
rect 393294 610634 393914 610718
rect 393294 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 393914 610634
rect 393294 574954 393914 610398
rect 393294 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 393914 574954
rect 393294 574634 393914 574718
rect 393294 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 393914 574634
rect 393294 538954 393914 574398
rect 393294 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 393914 538954
rect 393294 538634 393914 538718
rect 393294 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 393914 538634
rect 393294 502954 393914 538398
rect 393294 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 393914 502954
rect 393294 502634 393914 502718
rect 393294 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 393914 502634
rect 393294 466954 393914 502398
rect 393294 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 393914 466954
rect 393294 466634 393914 466718
rect 393294 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 393914 466634
rect 393294 430954 393914 466398
rect 393294 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 393914 430954
rect 393294 430634 393914 430718
rect 393294 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 393914 430634
rect 393294 394954 393914 430398
rect 393294 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 393914 394954
rect 393294 394634 393914 394718
rect 393294 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 393914 394634
rect 393294 358954 393914 394398
rect 393294 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 393914 358954
rect 393294 358634 393914 358718
rect 393294 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 393914 358634
rect 393294 322954 393914 358398
rect 393294 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 393914 322954
rect 393294 322634 393914 322718
rect 393294 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 393914 322634
rect 393294 286954 393914 322398
rect 393294 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 393914 286954
rect 393294 286634 393914 286718
rect 393294 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 393914 286634
rect 393294 250954 393914 286398
rect 393294 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 393914 250954
rect 393294 250634 393914 250718
rect 393294 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 393914 250634
rect 393294 214954 393914 250398
rect 393294 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 393914 214954
rect 393294 214634 393914 214718
rect 393294 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 393914 214634
rect 393294 178954 393914 214398
rect 393294 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 393914 178954
rect 393294 178634 393914 178718
rect 393294 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 393914 178634
rect 393294 142954 393914 178398
rect 393294 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 393914 142954
rect 393294 142634 393914 142718
rect 393294 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 393914 142634
rect 393294 106954 393914 142398
rect 393294 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 393914 106954
rect 393294 106634 393914 106718
rect 393294 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 393914 106634
rect 393294 70954 393914 106398
rect 393294 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 393914 70954
rect 393294 70634 393914 70718
rect 393294 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 393914 70634
rect 393294 34954 393914 70398
rect 393294 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 393914 34954
rect 393294 34634 393914 34718
rect 393294 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 393914 34634
rect 393294 -7066 393914 34398
rect 393294 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 393914 -7066
rect 393294 -7386 393914 -7302
rect 393294 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 393914 -7386
rect 393294 -7654 393914 -7622
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 402294 705798 402914 711590
rect 402294 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 402914 705798
rect 402294 705478 402914 705562
rect 402294 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 402914 705478
rect 402294 691954 402914 705242
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 402294 655954 402914 691398
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402294 619954 402914 655398
rect 402294 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 402914 619954
rect 402294 619634 402914 619718
rect 402294 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 402914 619634
rect 402294 583954 402914 619398
rect 402294 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 402914 583954
rect 402294 583634 402914 583718
rect 402294 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 402914 583634
rect 402294 547954 402914 583398
rect 402294 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 402914 547954
rect 402294 547634 402914 547718
rect 402294 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 402914 547634
rect 402294 511954 402914 547398
rect 402294 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 402914 511954
rect 402294 511634 402914 511718
rect 402294 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 402914 511634
rect 402294 475954 402914 511398
rect 402294 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 402914 475954
rect 402294 475634 402914 475718
rect 402294 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 402914 475634
rect 402294 439954 402914 475398
rect 402294 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 402914 439954
rect 402294 439634 402914 439718
rect 402294 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 402914 439634
rect 402294 403954 402914 439398
rect 402294 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 402914 403954
rect 402294 403634 402914 403718
rect 402294 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 402914 403634
rect 402294 367954 402914 403398
rect 402294 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 402914 367954
rect 402294 367634 402914 367718
rect 402294 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 402914 367634
rect 402294 331954 402914 367398
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 295954 402914 331398
rect 402294 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 402914 295954
rect 402294 295634 402914 295718
rect 402294 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 402914 295634
rect 402294 259954 402914 295398
rect 402294 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 402914 259954
rect 402294 259634 402914 259718
rect 402294 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 402914 259634
rect 402294 223954 402914 259398
rect 402294 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 402914 223954
rect 402294 223634 402914 223718
rect 402294 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 402914 223634
rect 402294 187954 402914 223398
rect 402294 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 402914 187954
rect 402294 187634 402914 187718
rect 402294 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 402914 187634
rect 402294 151954 402914 187398
rect 402294 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 402914 151954
rect 402294 151634 402914 151718
rect 402294 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 402914 151634
rect 402294 115954 402914 151398
rect 402294 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 402914 115954
rect 402294 115634 402914 115718
rect 402294 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 402914 115634
rect 402294 79954 402914 115398
rect 402294 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 402914 79954
rect 402294 79634 402914 79718
rect 402294 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 402914 79634
rect 402294 43954 402914 79398
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1306 402914 7398
rect 402294 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 402914 -1306
rect 402294 -1626 402914 -1542
rect 402294 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 402914 -1626
rect 402294 -7654 402914 -1862
rect 406794 706758 407414 711590
rect 406794 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 407414 706758
rect 406794 706438 407414 706522
rect 406794 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 407414 706438
rect 406794 696454 407414 706202
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 406794 660454 407414 695898
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 624454 407414 659898
rect 406794 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 407414 624454
rect 406794 624134 407414 624218
rect 406794 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 407414 624134
rect 406794 588454 407414 623898
rect 406794 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 407414 588454
rect 406794 588134 407414 588218
rect 406794 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 407414 588134
rect 406794 552454 407414 587898
rect 406794 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 407414 552454
rect 406794 552134 407414 552218
rect 406794 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 407414 552134
rect 406794 516454 407414 551898
rect 406794 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 407414 516454
rect 406794 516134 407414 516218
rect 406794 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 407414 516134
rect 406794 480454 407414 515898
rect 406794 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 407414 480454
rect 406794 480134 407414 480218
rect 406794 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 407414 480134
rect 406794 444454 407414 479898
rect 406794 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 407414 444454
rect 406794 444134 407414 444218
rect 406794 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 407414 444134
rect 406794 408454 407414 443898
rect 406794 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 407414 408454
rect 406794 408134 407414 408218
rect 406794 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 407414 408134
rect 406794 372454 407414 407898
rect 406794 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 407414 372454
rect 406794 372134 407414 372218
rect 406794 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 407414 372134
rect 406794 336454 407414 371898
rect 406794 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 407414 336454
rect 406794 336134 407414 336218
rect 406794 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 407414 336134
rect 406794 300454 407414 335898
rect 406794 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 407414 300454
rect 406794 300134 407414 300218
rect 406794 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 407414 300134
rect 406794 264454 407414 299898
rect 406794 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 407414 264454
rect 406794 264134 407414 264218
rect 406794 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 407414 264134
rect 406794 228454 407414 263898
rect 406794 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 407414 228454
rect 406794 228134 407414 228218
rect 406794 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 407414 228134
rect 406794 192454 407414 227898
rect 406794 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 407414 192454
rect 406794 192134 407414 192218
rect 406794 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 407414 192134
rect 406794 156454 407414 191898
rect 406794 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 407414 156454
rect 406794 156134 407414 156218
rect 406794 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 407414 156134
rect 406794 120454 407414 155898
rect 406794 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 407414 120454
rect 406794 120134 407414 120218
rect 406794 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 407414 120134
rect 406794 84454 407414 119898
rect 406794 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 407414 84454
rect 406794 84134 407414 84218
rect 406794 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 407414 84134
rect 406794 48454 407414 83898
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2266 407414 11898
rect 406794 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 407414 -2266
rect 406794 -2586 407414 -2502
rect 406794 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 407414 -2586
rect 406794 -7654 407414 -2822
rect 411294 707718 411914 711590
rect 411294 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 411914 707718
rect 411294 707398 411914 707482
rect 411294 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 411914 707398
rect 411294 700954 411914 707162
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 664954 411914 700398
rect 411294 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 411914 664954
rect 411294 664634 411914 664718
rect 411294 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 411914 664634
rect 411294 628954 411914 664398
rect 411294 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 411914 628954
rect 411294 628634 411914 628718
rect 411294 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 411914 628634
rect 411294 592954 411914 628398
rect 411294 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 411914 592954
rect 411294 592634 411914 592718
rect 411294 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 411914 592634
rect 411294 556954 411914 592398
rect 411294 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 411914 556954
rect 411294 556634 411914 556718
rect 411294 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 411914 556634
rect 411294 520954 411914 556398
rect 411294 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 411914 520954
rect 411294 520634 411914 520718
rect 411294 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 411914 520634
rect 411294 484954 411914 520398
rect 411294 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 411914 484954
rect 411294 484634 411914 484718
rect 411294 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 411914 484634
rect 411294 448954 411914 484398
rect 411294 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 411914 448954
rect 411294 448634 411914 448718
rect 411294 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 411914 448634
rect 411294 412954 411914 448398
rect 411294 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 411914 412954
rect 411294 412634 411914 412718
rect 411294 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 411914 412634
rect 411294 376954 411914 412398
rect 411294 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 411914 376954
rect 411294 376634 411914 376718
rect 411294 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 411914 376634
rect 411294 340954 411914 376398
rect 411294 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 411914 340954
rect 411294 340634 411914 340718
rect 411294 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 411914 340634
rect 411294 304954 411914 340398
rect 411294 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 411914 304954
rect 411294 304634 411914 304718
rect 411294 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 411914 304634
rect 411294 268954 411914 304398
rect 411294 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 411914 268954
rect 411294 268634 411914 268718
rect 411294 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 411914 268634
rect 411294 232954 411914 268398
rect 411294 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 411914 232954
rect 411294 232634 411914 232718
rect 411294 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 411914 232634
rect 411294 196954 411914 232398
rect 411294 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 411914 196954
rect 411294 196634 411914 196718
rect 411294 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 411914 196634
rect 411294 160954 411914 196398
rect 411294 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 411914 160954
rect 411294 160634 411914 160718
rect 411294 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 411914 160634
rect 411294 124954 411914 160398
rect 411294 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 411914 124954
rect 411294 124634 411914 124718
rect 411294 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 411914 124634
rect 411294 88954 411914 124398
rect 411294 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 411914 88954
rect 411294 88634 411914 88718
rect 411294 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 411914 88634
rect 411294 52954 411914 88398
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3226 411914 16398
rect 411294 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 411914 -3226
rect 411294 -3546 411914 -3462
rect 411294 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 411914 -3546
rect 411294 -7654 411914 -3782
rect 415794 708678 416414 711590
rect 415794 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 416414 708678
rect 415794 708358 416414 708442
rect 415794 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 416414 708358
rect 415794 669454 416414 708122
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4186 416414 20898
rect 415794 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 416414 -4186
rect 415794 -4506 416414 -4422
rect 415794 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 416414 -4506
rect 415794 -7654 416414 -4742
rect 420294 709638 420914 711590
rect 420294 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 420914 709638
rect 420294 709318 420914 709402
rect 420294 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 420914 709318
rect 420294 673954 420914 709082
rect 420294 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 420914 673954
rect 420294 673634 420914 673718
rect 420294 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 420914 673634
rect 420294 637954 420914 673398
rect 420294 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 420914 637954
rect 420294 637634 420914 637718
rect 420294 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 420914 637634
rect 420294 601954 420914 637398
rect 420294 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 420914 601954
rect 420294 601634 420914 601718
rect 420294 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 420914 601634
rect 420294 565954 420914 601398
rect 420294 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 420914 565954
rect 420294 565634 420914 565718
rect 420294 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 420914 565634
rect 420294 529954 420914 565398
rect 420294 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 420914 529954
rect 420294 529634 420914 529718
rect 420294 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 420914 529634
rect 420294 493954 420914 529398
rect 420294 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 420914 493954
rect 420294 493634 420914 493718
rect 420294 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 420914 493634
rect 420294 457954 420914 493398
rect 420294 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 420914 457954
rect 420294 457634 420914 457718
rect 420294 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 420914 457634
rect 420294 421954 420914 457398
rect 420294 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 420914 421954
rect 420294 421634 420914 421718
rect 420294 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 420914 421634
rect 420294 385954 420914 421398
rect 420294 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 420914 385954
rect 420294 385634 420914 385718
rect 420294 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 420914 385634
rect 420294 349954 420914 385398
rect 420294 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 420914 349954
rect 420294 349634 420914 349718
rect 420294 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 420914 349634
rect 420294 313954 420914 349398
rect 420294 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 420914 313954
rect 420294 313634 420914 313718
rect 420294 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 420914 313634
rect 420294 277954 420914 313398
rect 420294 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 420914 277954
rect 420294 277634 420914 277718
rect 420294 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 420914 277634
rect 420294 241954 420914 277398
rect 420294 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 420914 241954
rect 420294 241634 420914 241718
rect 420294 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 420914 241634
rect 420294 205954 420914 241398
rect 420294 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 420914 205954
rect 420294 205634 420914 205718
rect 420294 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 420914 205634
rect 420294 169954 420914 205398
rect 420294 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 420914 169954
rect 420294 169634 420914 169718
rect 420294 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 420914 169634
rect 420294 133954 420914 169398
rect 420294 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 420914 133954
rect 420294 133634 420914 133718
rect 420294 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 420914 133634
rect 420294 97954 420914 133398
rect 420294 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 420914 97954
rect 420294 97634 420914 97718
rect 420294 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 420914 97634
rect 420294 61954 420914 97398
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5146 420914 25398
rect 420294 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 420914 -5146
rect 420294 -5466 420914 -5382
rect 420294 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 420914 -5466
rect 420294 -7654 420914 -5702
rect 424794 710598 425414 711590
rect 424794 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 425414 710598
rect 424794 710278 425414 710362
rect 424794 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 425414 710278
rect 424794 678454 425414 710042
rect 424794 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 425414 678454
rect 424794 678134 425414 678218
rect 424794 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 425414 678134
rect 424794 642454 425414 677898
rect 424794 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 425414 642454
rect 424794 642134 425414 642218
rect 424794 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 425414 642134
rect 424794 606454 425414 641898
rect 424794 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 425414 606454
rect 424794 606134 425414 606218
rect 424794 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 425414 606134
rect 424794 570454 425414 605898
rect 424794 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 425414 570454
rect 424794 570134 425414 570218
rect 424794 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 425414 570134
rect 424794 534454 425414 569898
rect 424794 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 425414 534454
rect 424794 534134 425414 534218
rect 424794 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 425414 534134
rect 424794 498454 425414 533898
rect 424794 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 425414 498454
rect 424794 498134 425414 498218
rect 424794 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 425414 498134
rect 424794 462454 425414 497898
rect 424794 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 425414 462454
rect 424794 462134 425414 462218
rect 424794 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 425414 462134
rect 424794 426454 425414 461898
rect 424794 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 425414 426454
rect 424794 426134 425414 426218
rect 424794 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 425414 426134
rect 424794 390454 425414 425898
rect 424794 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 425414 390454
rect 424794 390134 425414 390218
rect 424794 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 425414 390134
rect 424794 354454 425414 389898
rect 424794 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 425414 354454
rect 424794 354134 425414 354218
rect 424794 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 425414 354134
rect 424794 318454 425414 353898
rect 424794 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 425414 318454
rect 424794 318134 425414 318218
rect 424794 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 425414 318134
rect 424794 282454 425414 317898
rect 424794 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 425414 282454
rect 424794 282134 425414 282218
rect 424794 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 425414 282134
rect 424794 246454 425414 281898
rect 424794 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 425414 246454
rect 424794 246134 425414 246218
rect 424794 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 425414 246134
rect 424794 210454 425414 245898
rect 424794 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 425414 210454
rect 424794 210134 425414 210218
rect 424794 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 425414 210134
rect 424794 174454 425414 209898
rect 424794 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 425414 174454
rect 424794 174134 425414 174218
rect 424794 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 425414 174134
rect 424794 138454 425414 173898
rect 424794 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 425414 138454
rect 424794 138134 425414 138218
rect 424794 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 425414 138134
rect 424794 102454 425414 137898
rect 424794 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 425414 102454
rect 424794 102134 425414 102218
rect 424794 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 425414 102134
rect 424794 66454 425414 101898
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6106 425414 29898
rect 424794 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 425414 -6106
rect 424794 -6426 425414 -6342
rect 424794 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 425414 -6426
rect 424794 -7654 425414 -6662
rect 429294 711558 429914 711590
rect 429294 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 429914 711558
rect 429294 711238 429914 711322
rect 429294 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 429914 711238
rect 429294 682954 429914 711002
rect 429294 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 429914 682954
rect 429294 682634 429914 682718
rect 429294 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 429914 682634
rect 429294 646954 429914 682398
rect 429294 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 429914 646954
rect 429294 646634 429914 646718
rect 429294 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 429914 646634
rect 429294 610954 429914 646398
rect 429294 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 429914 610954
rect 429294 610634 429914 610718
rect 429294 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 429914 610634
rect 429294 574954 429914 610398
rect 429294 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 429914 574954
rect 429294 574634 429914 574718
rect 429294 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 429914 574634
rect 429294 538954 429914 574398
rect 429294 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 429914 538954
rect 429294 538634 429914 538718
rect 429294 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 429914 538634
rect 429294 502954 429914 538398
rect 429294 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 429914 502954
rect 429294 502634 429914 502718
rect 429294 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 429914 502634
rect 429294 466954 429914 502398
rect 429294 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 429914 466954
rect 429294 466634 429914 466718
rect 429294 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 429914 466634
rect 429294 430954 429914 466398
rect 429294 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 429914 430954
rect 429294 430634 429914 430718
rect 429294 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 429914 430634
rect 429294 394954 429914 430398
rect 429294 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 429914 394954
rect 429294 394634 429914 394718
rect 429294 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 429914 394634
rect 429294 358954 429914 394398
rect 429294 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 429914 358954
rect 429294 358634 429914 358718
rect 429294 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 429914 358634
rect 429294 322954 429914 358398
rect 429294 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 429914 322954
rect 429294 322634 429914 322718
rect 429294 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 429914 322634
rect 429294 286954 429914 322398
rect 429294 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 429914 286954
rect 429294 286634 429914 286718
rect 429294 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 429914 286634
rect 429294 250954 429914 286398
rect 429294 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 429914 250954
rect 429294 250634 429914 250718
rect 429294 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 429914 250634
rect 429294 214954 429914 250398
rect 429294 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 429914 214954
rect 429294 214634 429914 214718
rect 429294 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 429914 214634
rect 429294 178954 429914 214398
rect 429294 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 429914 178954
rect 429294 178634 429914 178718
rect 429294 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 429914 178634
rect 429294 142954 429914 178398
rect 429294 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 429914 142954
rect 429294 142634 429914 142718
rect 429294 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 429914 142634
rect 429294 106954 429914 142398
rect 429294 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 429914 106954
rect 429294 106634 429914 106718
rect 429294 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 429914 106634
rect 429294 70954 429914 106398
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7066 429914 34398
rect 429294 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 429914 -7066
rect 429294 -7386 429914 -7302
rect 429294 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 429914 -7386
rect 429294 -7654 429914 -7622
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 438294 705798 438914 711590
rect 438294 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 438914 705798
rect 438294 705478 438914 705562
rect 438294 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 438914 705478
rect 438294 691954 438914 705242
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 655954 438914 691398
rect 438294 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 438914 655954
rect 438294 655634 438914 655718
rect 438294 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 438914 655634
rect 438294 619954 438914 655398
rect 438294 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 438914 619954
rect 438294 619634 438914 619718
rect 438294 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 438914 619634
rect 438294 583954 438914 619398
rect 438294 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 438914 583954
rect 438294 583634 438914 583718
rect 438294 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 438914 583634
rect 438294 547954 438914 583398
rect 438294 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 438914 547954
rect 438294 547634 438914 547718
rect 438294 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 438914 547634
rect 438294 511954 438914 547398
rect 438294 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 438914 511954
rect 438294 511634 438914 511718
rect 438294 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 438914 511634
rect 438294 475954 438914 511398
rect 438294 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 438914 475954
rect 438294 475634 438914 475718
rect 438294 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 438914 475634
rect 438294 439954 438914 475398
rect 438294 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 438914 439954
rect 438294 439634 438914 439718
rect 438294 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 438914 439634
rect 438294 403954 438914 439398
rect 438294 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 438914 403954
rect 438294 403634 438914 403718
rect 438294 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 438914 403634
rect 438294 367954 438914 403398
rect 438294 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 438914 367954
rect 438294 367634 438914 367718
rect 438294 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 438914 367634
rect 438294 331954 438914 367398
rect 438294 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 438914 331954
rect 438294 331634 438914 331718
rect 438294 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 438914 331634
rect 438294 295954 438914 331398
rect 438294 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 438914 295954
rect 438294 295634 438914 295718
rect 438294 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 438914 295634
rect 438294 259954 438914 295398
rect 438294 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 438914 259954
rect 438294 259634 438914 259718
rect 438294 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 438914 259634
rect 438294 223954 438914 259398
rect 438294 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 438914 223954
rect 438294 223634 438914 223718
rect 438294 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 438914 223634
rect 438294 187954 438914 223398
rect 438294 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 438914 187954
rect 438294 187634 438914 187718
rect 438294 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 438914 187634
rect 438294 151954 438914 187398
rect 438294 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 438914 151954
rect 438294 151634 438914 151718
rect 438294 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 438914 151634
rect 438294 115954 438914 151398
rect 438294 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 438914 115954
rect 438294 115634 438914 115718
rect 438294 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 438914 115634
rect 438294 79954 438914 115398
rect 438294 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 438914 79954
rect 438294 79634 438914 79718
rect 438294 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 438914 79634
rect 438294 43954 438914 79398
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1306 438914 7398
rect 438294 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 438914 -1306
rect 438294 -1626 438914 -1542
rect 438294 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 438914 -1626
rect 438294 -7654 438914 -1862
rect 442794 706758 443414 711590
rect 442794 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 443414 706758
rect 442794 706438 443414 706522
rect 442794 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 443414 706438
rect 442794 696454 443414 706202
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 660454 443414 695898
rect 442794 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 443414 660454
rect 442794 660134 443414 660218
rect 442794 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 443414 660134
rect 442794 624454 443414 659898
rect 442794 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 443414 624454
rect 442794 624134 443414 624218
rect 442794 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 443414 624134
rect 442794 588454 443414 623898
rect 442794 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 443414 588454
rect 442794 588134 443414 588218
rect 442794 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 443414 588134
rect 442794 552454 443414 587898
rect 442794 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 443414 552454
rect 442794 552134 443414 552218
rect 442794 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 443414 552134
rect 442794 516454 443414 551898
rect 442794 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 443414 516454
rect 442794 516134 443414 516218
rect 442794 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 443414 516134
rect 442794 480454 443414 515898
rect 442794 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 443414 480454
rect 442794 480134 443414 480218
rect 442794 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 443414 480134
rect 442794 444454 443414 479898
rect 442794 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 443414 444454
rect 442794 444134 443414 444218
rect 442794 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 443414 444134
rect 442794 408454 443414 443898
rect 442794 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 443414 408454
rect 442794 408134 443414 408218
rect 442794 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 443414 408134
rect 442794 372454 443414 407898
rect 442794 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 443414 372454
rect 442794 372134 443414 372218
rect 442794 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 443414 372134
rect 442794 336454 443414 371898
rect 442794 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 443414 336454
rect 442794 336134 443414 336218
rect 442794 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 443414 336134
rect 442794 300454 443414 335898
rect 442794 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 443414 300454
rect 442794 300134 443414 300218
rect 442794 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 443414 300134
rect 442794 264454 443414 299898
rect 442794 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 443414 264454
rect 442794 264134 443414 264218
rect 442794 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 443414 264134
rect 442794 228454 443414 263898
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 192454 443414 227898
rect 442794 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 443414 192454
rect 442794 192134 443414 192218
rect 442794 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 443414 192134
rect 442794 156454 443414 191898
rect 442794 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 443414 156454
rect 442794 156134 443414 156218
rect 442794 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 443414 156134
rect 442794 120454 443414 155898
rect 442794 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 443414 120454
rect 442794 120134 443414 120218
rect 442794 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 443414 120134
rect 442794 84454 443414 119898
rect 442794 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 443414 84454
rect 442794 84134 443414 84218
rect 442794 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 443414 84134
rect 442794 48454 443414 83898
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2266 443414 11898
rect 442794 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 443414 -2266
rect 442794 -2586 443414 -2502
rect 442794 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 443414 -2586
rect 442794 -7654 443414 -2822
rect 447294 707718 447914 711590
rect 447294 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 447914 707718
rect 447294 707398 447914 707482
rect 447294 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 447914 707398
rect 447294 700954 447914 707162
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 664954 447914 700398
rect 447294 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 447914 664954
rect 447294 664634 447914 664718
rect 447294 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 447914 664634
rect 447294 628954 447914 664398
rect 447294 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 447914 628954
rect 447294 628634 447914 628718
rect 447294 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 447914 628634
rect 447294 592954 447914 628398
rect 447294 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 447914 592954
rect 447294 592634 447914 592718
rect 447294 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 447914 592634
rect 447294 556954 447914 592398
rect 447294 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 447914 556954
rect 447294 556634 447914 556718
rect 447294 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 447914 556634
rect 447294 520954 447914 556398
rect 447294 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 447914 520954
rect 447294 520634 447914 520718
rect 447294 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 447914 520634
rect 447294 484954 447914 520398
rect 447294 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 447914 484954
rect 447294 484634 447914 484718
rect 447294 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 447914 484634
rect 447294 448954 447914 484398
rect 447294 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 447914 448954
rect 447294 448634 447914 448718
rect 447294 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 447914 448634
rect 447294 412954 447914 448398
rect 447294 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 447914 412954
rect 447294 412634 447914 412718
rect 447294 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 447914 412634
rect 447294 376954 447914 412398
rect 447294 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 447914 376954
rect 447294 376634 447914 376718
rect 447294 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 447914 376634
rect 447294 340954 447914 376398
rect 447294 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 447914 340954
rect 447294 340634 447914 340718
rect 447294 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 447914 340634
rect 447294 304954 447914 340398
rect 447294 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 447914 304954
rect 447294 304634 447914 304718
rect 447294 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 447914 304634
rect 447294 268954 447914 304398
rect 447294 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 447914 268954
rect 447294 268634 447914 268718
rect 447294 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 447914 268634
rect 447294 232954 447914 268398
rect 447294 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 447914 232954
rect 447294 232634 447914 232718
rect 447294 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 447914 232634
rect 447294 196954 447914 232398
rect 447294 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 447914 196954
rect 447294 196634 447914 196718
rect 447294 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 447914 196634
rect 447294 160954 447914 196398
rect 447294 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 447914 160954
rect 447294 160634 447914 160718
rect 447294 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 447914 160634
rect 447294 124954 447914 160398
rect 447294 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 447914 124954
rect 447294 124634 447914 124718
rect 447294 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 447914 124634
rect 447294 88954 447914 124398
rect 447294 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 447914 88954
rect 447294 88634 447914 88718
rect 447294 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 447914 88634
rect 447294 52954 447914 88398
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3226 447914 16398
rect 447294 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 447914 -3226
rect 447294 -3546 447914 -3462
rect 447294 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 447914 -3546
rect 447294 -7654 447914 -3782
rect 451794 708678 452414 711590
rect 451794 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 452414 708678
rect 451794 708358 452414 708442
rect 451794 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 452414 708358
rect 451794 669454 452414 708122
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4186 452414 20898
rect 451794 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 452414 -4186
rect 451794 -4506 452414 -4422
rect 451794 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 452414 -4506
rect 451794 -7654 452414 -4742
rect 456294 709638 456914 711590
rect 456294 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 456914 709638
rect 456294 709318 456914 709402
rect 456294 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 456914 709318
rect 456294 673954 456914 709082
rect 456294 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 456914 673954
rect 456294 673634 456914 673718
rect 456294 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 456914 673634
rect 456294 637954 456914 673398
rect 456294 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 456914 637954
rect 456294 637634 456914 637718
rect 456294 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 456914 637634
rect 456294 601954 456914 637398
rect 456294 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 456914 601954
rect 456294 601634 456914 601718
rect 456294 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 456914 601634
rect 456294 565954 456914 601398
rect 456294 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 456914 565954
rect 456294 565634 456914 565718
rect 456294 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 456914 565634
rect 456294 529954 456914 565398
rect 456294 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 456914 529954
rect 456294 529634 456914 529718
rect 456294 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 456914 529634
rect 456294 493954 456914 529398
rect 456294 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 456914 493954
rect 456294 493634 456914 493718
rect 456294 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 456914 493634
rect 456294 457954 456914 493398
rect 456294 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 456914 457954
rect 456294 457634 456914 457718
rect 456294 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 456914 457634
rect 456294 421954 456914 457398
rect 456294 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 456914 421954
rect 456294 421634 456914 421718
rect 456294 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 456914 421634
rect 456294 385954 456914 421398
rect 456294 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 456914 385954
rect 456294 385634 456914 385718
rect 456294 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 456914 385634
rect 456294 349954 456914 385398
rect 456294 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 456914 349954
rect 456294 349634 456914 349718
rect 456294 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 456914 349634
rect 456294 313954 456914 349398
rect 456294 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 456914 313954
rect 456294 313634 456914 313718
rect 456294 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 456914 313634
rect 456294 277954 456914 313398
rect 456294 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 456914 277954
rect 456294 277634 456914 277718
rect 456294 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 456914 277634
rect 456294 241954 456914 277398
rect 456294 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 456914 241954
rect 456294 241634 456914 241718
rect 456294 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 456914 241634
rect 456294 205954 456914 241398
rect 456294 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 456914 205954
rect 456294 205634 456914 205718
rect 456294 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 456914 205634
rect 456294 169954 456914 205398
rect 456294 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 456914 169954
rect 456294 169634 456914 169718
rect 456294 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 456914 169634
rect 456294 133954 456914 169398
rect 456294 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 456914 133954
rect 456294 133634 456914 133718
rect 456294 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 456914 133634
rect 456294 97954 456914 133398
rect 456294 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 456914 97954
rect 456294 97634 456914 97718
rect 456294 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 456914 97634
rect 456294 61954 456914 97398
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5146 456914 25398
rect 456294 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 456914 -5146
rect 456294 -5466 456914 -5382
rect 456294 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 456914 -5466
rect 456294 -7654 456914 -5702
rect 460794 710598 461414 711590
rect 460794 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 461414 710598
rect 460794 710278 461414 710362
rect 460794 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 461414 710278
rect 460794 678454 461414 710042
rect 460794 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 461414 678454
rect 460794 678134 461414 678218
rect 460794 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 461414 678134
rect 460794 642454 461414 677898
rect 460794 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 461414 642454
rect 460794 642134 461414 642218
rect 460794 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 461414 642134
rect 460794 606454 461414 641898
rect 460794 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 461414 606454
rect 460794 606134 461414 606218
rect 460794 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 461414 606134
rect 460794 570454 461414 605898
rect 460794 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 461414 570454
rect 460794 570134 461414 570218
rect 460794 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 461414 570134
rect 460794 534454 461414 569898
rect 460794 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 461414 534454
rect 460794 534134 461414 534218
rect 460794 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 461414 534134
rect 460794 498454 461414 533898
rect 460794 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 461414 498454
rect 460794 498134 461414 498218
rect 460794 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 461414 498134
rect 460794 462454 461414 497898
rect 460794 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 461414 462454
rect 460794 462134 461414 462218
rect 460794 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 461414 462134
rect 460794 426454 461414 461898
rect 460794 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 461414 426454
rect 460794 426134 461414 426218
rect 460794 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 461414 426134
rect 460794 390454 461414 425898
rect 460794 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 461414 390454
rect 460794 390134 461414 390218
rect 460794 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 461414 390134
rect 460794 354454 461414 389898
rect 460794 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 461414 354454
rect 460794 354134 461414 354218
rect 460794 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 461414 354134
rect 460794 318454 461414 353898
rect 460794 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 461414 318454
rect 460794 318134 461414 318218
rect 460794 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 461414 318134
rect 460794 282454 461414 317898
rect 460794 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 461414 282454
rect 460794 282134 461414 282218
rect 460794 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 461414 282134
rect 460794 246454 461414 281898
rect 460794 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 461414 246454
rect 460794 246134 461414 246218
rect 460794 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 461414 246134
rect 460794 210454 461414 245898
rect 460794 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 461414 210454
rect 460794 210134 461414 210218
rect 460794 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 461414 210134
rect 460794 174454 461414 209898
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 460794 138454 461414 173898
rect 460794 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 461414 138454
rect 460794 138134 461414 138218
rect 460794 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 461414 138134
rect 460794 102454 461414 137898
rect 460794 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 461414 102454
rect 460794 102134 461414 102218
rect 460794 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 461414 102134
rect 460794 66454 461414 101898
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6106 461414 29898
rect 460794 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 461414 -6106
rect 460794 -6426 461414 -6342
rect 460794 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 461414 -6426
rect 460794 -7654 461414 -6662
rect 465294 711558 465914 711590
rect 465294 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 465914 711558
rect 465294 711238 465914 711322
rect 465294 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 465914 711238
rect 465294 682954 465914 711002
rect 465294 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 465914 682954
rect 465294 682634 465914 682718
rect 465294 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 465914 682634
rect 465294 646954 465914 682398
rect 465294 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 465914 646954
rect 465294 646634 465914 646718
rect 465294 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 465914 646634
rect 465294 610954 465914 646398
rect 465294 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 465914 610954
rect 465294 610634 465914 610718
rect 465294 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 465914 610634
rect 465294 574954 465914 610398
rect 465294 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 465914 574954
rect 465294 574634 465914 574718
rect 465294 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 465914 574634
rect 465294 538954 465914 574398
rect 465294 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 465914 538954
rect 465294 538634 465914 538718
rect 465294 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 465914 538634
rect 465294 502954 465914 538398
rect 465294 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 465914 502954
rect 465294 502634 465914 502718
rect 465294 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 465914 502634
rect 465294 466954 465914 502398
rect 465294 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 465914 466954
rect 465294 466634 465914 466718
rect 465294 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 465914 466634
rect 465294 430954 465914 466398
rect 465294 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 465914 430954
rect 465294 430634 465914 430718
rect 465294 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 465914 430634
rect 465294 394954 465914 430398
rect 465294 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 465914 394954
rect 465294 394634 465914 394718
rect 465294 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 465914 394634
rect 465294 358954 465914 394398
rect 465294 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 465914 358954
rect 465294 358634 465914 358718
rect 465294 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 465914 358634
rect 465294 322954 465914 358398
rect 465294 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 465914 322954
rect 465294 322634 465914 322718
rect 465294 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 465914 322634
rect 465294 286954 465914 322398
rect 465294 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 465914 286954
rect 465294 286634 465914 286718
rect 465294 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 465914 286634
rect 465294 250954 465914 286398
rect 465294 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 465914 250954
rect 465294 250634 465914 250718
rect 465294 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 465914 250634
rect 465294 214954 465914 250398
rect 465294 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 465914 214954
rect 465294 214634 465914 214718
rect 465294 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 465914 214634
rect 465294 178954 465914 214398
rect 465294 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 465914 178954
rect 465294 178634 465914 178718
rect 465294 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 465914 178634
rect 465294 142954 465914 178398
rect 465294 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 465914 142954
rect 465294 142634 465914 142718
rect 465294 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 465914 142634
rect 465294 106954 465914 142398
rect 465294 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 465914 106954
rect 465294 106634 465914 106718
rect 465294 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 465914 106634
rect 465294 70954 465914 106398
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7066 465914 34398
rect 465294 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 465914 -7066
rect 465294 -7386 465914 -7302
rect 465294 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 465914 -7386
rect 465294 -7654 465914 -7622
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 474294 705798 474914 711590
rect 474294 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 474914 705798
rect 474294 705478 474914 705562
rect 474294 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 474914 705478
rect 474294 691954 474914 705242
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 655954 474914 691398
rect 474294 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 474914 655954
rect 474294 655634 474914 655718
rect 474294 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 474914 655634
rect 474294 619954 474914 655398
rect 474294 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 474914 619954
rect 474294 619634 474914 619718
rect 474294 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 474914 619634
rect 474294 583954 474914 619398
rect 474294 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 474914 583954
rect 474294 583634 474914 583718
rect 474294 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 474914 583634
rect 474294 547954 474914 583398
rect 474294 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 474914 547954
rect 474294 547634 474914 547718
rect 474294 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 474914 547634
rect 474294 511954 474914 547398
rect 474294 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 474914 511954
rect 474294 511634 474914 511718
rect 474294 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 474914 511634
rect 474294 475954 474914 511398
rect 474294 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 474914 475954
rect 474294 475634 474914 475718
rect 474294 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 474914 475634
rect 474294 439954 474914 475398
rect 474294 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 474914 439954
rect 474294 439634 474914 439718
rect 474294 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 474914 439634
rect 474294 403954 474914 439398
rect 474294 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 474914 403954
rect 474294 403634 474914 403718
rect 474294 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 474914 403634
rect 474294 367954 474914 403398
rect 474294 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 474914 367954
rect 474294 367634 474914 367718
rect 474294 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 474914 367634
rect 474294 331954 474914 367398
rect 474294 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 474914 331954
rect 474294 331634 474914 331718
rect 474294 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 474914 331634
rect 474294 295954 474914 331398
rect 474294 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 474914 295954
rect 474294 295634 474914 295718
rect 474294 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 474914 295634
rect 474294 259954 474914 295398
rect 474294 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 474914 259954
rect 474294 259634 474914 259718
rect 474294 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 474914 259634
rect 474294 223954 474914 259398
rect 474294 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 474914 223954
rect 474294 223634 474914 223718
rect 474294 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 474914 223634
rect 474294 187954 474914 223398
rect 474294 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 474914 187954
rect 474294 187634 474914 187718
rect 474294 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 474914 187634
rect 474294 151954 474914 187398
rect 474294 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 474914 151954
rect 474294 151634 474914 151718
rect 474294 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 474914 151634
rect 474294 115954 474914 151398
rect 474294 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 474914 115954
rect 474294 115634 474914 115718
rect 474294 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 474914 115634
rect 474294 79954 474914 115398
rect 474294 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 474914 79954
rect 474294 79634 474914 79718
rect 474294 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 474914 79634
rect 474294 43954 474914 79398
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1306 474914 7398
rect 474294 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 474914 -1306
rect 474294 -1626 474914 -1542
rect 474294 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 474914 -1626
rect 474294 -7654 474914 -1862
rect 478794 706758 479414 711590
rect 478794 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 479414 706758
rect 478794 706438 479414 706522
rect 478794 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 479414 706438
rect 478794 696454 479414 706202
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 660454 479414 695898
rect 478794 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 479414 660454
rect 478794 660134 479414 660218
rect 478794 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 479414 660134
rect 478794 624454 479414 659898
rect 478794 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 479414 624454
rect 478794 624134 479414 624218
rect 478794 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 479414 624134
rect 478794 588454 479414 623898
rect 478794 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 479414 588454
rect 478794 588134 479414 588218
rect 478794 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 479414 588134
rect 478794 552454 479414 587898
rect 478794 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 479414 552454
rect 478794 552134 479414 552218
rect 478794 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 479414 552134
rect 478794 516454 479414 551898
rect 478794 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 479414 516454
rect 478794 516134 479414 516218
rect 478794 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 479414 516134
rect 478794 480454 479414 515898
rect 478794 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 479414 480454
rect 478794 480134 479414 480218
rect 478794 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 479414 480134
rect 478794 444454 479414 479898
rect 478794 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 479414 444454
rect 478794 444134 479414 444218
rect 478794 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 479414 444134
rect 478794 408454 479414 443898
rect 478794 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 479414 408454
rect 478794 408134 479414 408218
rect 478794 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 479414 408134
rect 478794 372454 479414 407898
rect 478794 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 479414 372454
rect 478794 372134 479414 372218
rect 478794 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 479414 372134
rect 478794 336454 479414 371898
rect 478794 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 479414 336454
rect 478794 336134 479414 336218
rect 478794 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 479414 336134
rect 478794 300454 479414 335898
rect 478794 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 479414 300454
rect 478794 300134 479414 300218
rect 478794 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 479414 300134
rect 478794 264454 479414 299898
rect 478794 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 479414 264454
rect 478794 264134 479414 264218
rect 478794 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 479414 264134
rect 478794 228454 479414 263898
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 192454 479414 227898
rect 478794 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 479414 192454
rect 478794 192134 479414 192218
rect 478794 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 479414 192134
rect 478794 156454 479414 191898
rect 478794 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 479414 156454
rect 478794 156134 479414 156218
rect 478794 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 479414 156134
rect 478794 120454 479414 155898
rect 478794 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 479414 120454
rect 478794 120134 479414 120218
rect 478794 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 479414 120134
rect 478794 84454 479414 119898
rect 478794 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 479414 84454
rect 478794 84134 479414 84218
rect 478794 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 479414 84134
rect 478794 48454 479414 83898
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2266 479414 11898
rect 478794 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 479414 -2266
rect 478794 -2586 479414 -2502
rect 478794 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 479414 -2586
rect 478794 -7654 479414 -2822
rect 483294 707718 483914 711590
rect 483294 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 483914 707718
rect 483294 707398 483914 707482
rect 483294 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 483914 707398
rect 483294 700954 483914 707162
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 664954 483914 700398
rect 483294 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 483914 664954
rect 483294 664634 483914 664718
rect 483294 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 483914 664634
rect 483294 628954 483914 664398
rect 483294 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 483914 628954
rect 483294 628634 483914 628718
rect 483294 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 483914 628634
rect 483294 592954 483914 628398
rect 483294 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 483914 592954
rect 483294 592634 483914 592718
rect 483294 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 483914 592634
rect 483294 556954 483914 592398
rect 483294 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 483914 556954
rect 483294 556634 483914 556718
rect 483294 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 483914 556634
rect 483294 520954 483914 556398
rect 483294 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 483914 520954
rect 483294 520634 483914 520718
rect 483294 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 483914 520634
rect 483294 484954 483914 520398
rect 483294 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 483914 484954
rect 483294 484634 483914 484718
rect 483294 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 483914 484634
rect 483294 448954 483914 484398
rect 483294 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 483914 448954
rect 483294 448634 483914 448718
rect 483294 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 483914 448634
rect 483294 412954 483914 448398
rect 483294 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 483914 412954
rect 483294 412634 483914 412718
rect 483294 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 483914 412634
rect 483294 376954 483914 412398
rect 483294 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 483914 376954
rect 483294 376634 483914 376718
rect 483294 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 483914 376634
rect 483294 340954 483914 376398
rect 483294 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 483914 340954
rect 483294 340634 483914 340718
rect 483294 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 483914 340634
rect 483294 304954 483914 340398
rect 483294 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 483914 304954
rect 483294 304634 483914 304718
rect 483294 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 483914 304634
rect 483294 268954 483914 304398
rect 483294 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 483914 268954
rect 483294 268634 483914 268718
rect 483294 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 483914 268634
rect 483294 232954 483914 268398
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 124954 483914 160398
rect 483294 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 483914 124954
rect 483294 124634 483914 124718
rect 483294 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 483914 124634
rect 483294 88954 483914 124398
rect 483294 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 483914 88954
rect 483294 88634 483914 88718
rect 483294 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 483914 88634
rect 483294 52954 483914 88398
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3226 483914 16398
rect 483294 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 483914 -3226
rect 483294 -3546 483914 -3462
rect 483294 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 483914 -3546
rect 483294 -7654 483914 -3782
rect 487794 708678 488414 711590
rect 487794 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 488414 708678
rect 487794 708358 488414 708442
rect 487794 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 488414 708358
rect 487794 669454 488414 708122
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4186 488414 20898
rect 487794 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 488414 -4186
rect 487794 -4506 488414 -4422
rect 487794 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 488414 -4506
rect 487794 -7654 488414 -4742
rect 492294 709638 492914 711590
rect 492294 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 492914 709638
rect 492294 709318 492914 709402
rect 492294 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 492914 709318
rect 492294 673954 492914 709082
rect 492294 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 492914 673954
rect 492294 673634 492914 673718
rect 492294 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 492914 673634
rect 492294 637954 492914 673398
rect 492294 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 492914 637954
rect 492294 637634 492914 637718
rect 492294 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 492914 637634
rect 492294 601954 492914 637398
rect 492294 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 492914 601954
rect 492294 601634 492914 601718
rect 492294 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 492914 601634
rect 492294 565954 492914 601398
rect 492294 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 492914 565954
rect 492294 565634 492914 565718
rect 492294 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 492914 565634
rect 492294 529954 492914 565398
rect 492294 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 492914 529954
rect 492294 529634 492914 529718
rect 492294 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 492914 529634
rect 492294 493954 492914 529398
rect 492294 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 492914 493954
rect 492294 493634 492914 493718
rect 492294 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 492914 493634
rect 492294 457954 492914 493398
rect 492294 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 492914 457954
rect 492294 457634 492914 457718
rect 492294 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 492914 457634
rect 492294 421954 492914 457398
rect 492294 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 492914 421954
rect 492294 421634 492914 421718
rect 492294 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 492914 421634
rect 492294 385954 492914 421398
rect 492294 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 492914 385954
rect 492294 385634 492914 385718
rect 492294 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 492914 385634
rect 492294 349954 492914 385398
rect 492294 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 492914 349954
rect 492294 349634 492914 349718
rect 492294 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 492914 349634
rect 492294 313954 492914 349398
rect 492294 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 492914 313954
rect 492294 313634 492914 313718
rect 492294 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 492914 313634
rect 492294 277954 492914 313398
rect 492294 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 492914 277954
rect 492294 277634 492914 277718
rect 492294 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 492914 277634
rect 492294 241954 492914 277398
rect 492294 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 492914 241954
rect 492294 241634 492914 241718
rect 492294 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 492914 241634
rect 492294 205954 492914 241398
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 133954 492914 169398
rect 492294 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 492914 133954
rect 492294 133634 492914 133718
rect 492294 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 492914 133634
rect 492294 97954 492914 133398
rect 492294 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 492914 97954
rect 492294 97634 492914 97718
rect 492294 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 492914 97634
rect 492294 61954 492914 97398
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5146 492914 25398
rect 492294 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 492914 -5146
rect 492294 -5466 492914 -5382
rect 492294 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 492914 -5466
rect 492294 -7654 492914 -5702
rect 496794 710598 497414 711590
rect 496794 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 497414 710598
rect 496794 710278 497414 710362
rect 496794 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 497414 710278
rect 496794 678454 497414 710042
rect 496794 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 497414 678454
rect 496794 678134 497414 678218
rect 496794 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 497414 678134
rect 496794 642454 497414 677898
rect 496794 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 497414 642454
rect 496794 642134 497414 642218
rect 496794 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 497414 642134
rect 496794 606454 497414 641898
rect 496794 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 497414 606454
rect 496794 606134 497414 606218
rect 496794 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 497414 606134
rect 496794 570454 497414 605898
rect 496794 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 497414 570454
rect 496794 570134 497414 570218
rect 496794 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 497414 570134
rect 496794 534454 497414 569898
rect 496794 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 497414 534454
rect 496794 534134 497414 534218
rect 496794 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 497414 534134
rect 496794 498454 497414 533898
rect 496794 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 497414 498454
rect 496794 498134 497414 498218
rect 496794 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 497414 498134
rect 496794 462454 497414 497898
rect 496794 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 497414 462454
rect 496794 462134 497414 462218
rect 496794 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 497414 462134
rect 496794 426454 497414 461898
rect 496794 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 497414 426454
rect 496794 426134 497414 426218
rect 496794 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 497414 426134
rect 496794 390454 497414 425898
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 354454 497414 389898
rect 496794 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 497414 354454
rect 496794 354134 497414 354218
rect 496794 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 497414 354134
rect 496794 318454 497414 353898
rect 496794 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 497414 318454
rect 496794 318134 497414 318218
rect 496794 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 497414 318134
rect 496794 282454 497414 317898
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 246454 497414 281898
rect 496794 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 497414 246454
rect 496794 246134 497414 246218
rect 496794 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 497414 246134
rect 496794 210454 497414 245898
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 138454 497414 173898
rect 496794 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 497414 138454
rect 496794 138134 497414 138218
rect 496794 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 497414 138134
rect 496794 102454 497414 137898
rect 496794 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 497414 102454
rect 496794 102134 497414 102218
rect 496794 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 497414 102134
rect 496794 66454 497414 101898
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6106 497414 29898
rect 496794 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 497414 -6106
rect 496794 -6426 497414 -6342
rect 496794 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 497414 -6426
rect 496794 -7654 497414 -6662
rect 501294 711558 501914 711590
rect 501294 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 501914 711558
rect 501294 711238 501914 711322
rect 501294 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 501914 711238
rect 501294 682954 501914 711002
rect 501294 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 501914 682954
rect 501294 682634 501914 682718
rect 501294 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 501914 682634
rect 501294 646954 501914 682398
rect 501294 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 501914 646954
rect 501294 646634 501914 646718
rect 501294 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 501914 646634
rect 501294 610954 501914 646398
rect 501294 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 501914 610954
rect 501294 610634 501914 610718
rect 501294 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 501914 610634
rect 501294 574954 501914 610398
rect 501294 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 501914 574954
rect 501294 574634 501914 574718
rect 501294 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 501914 574634
rect 501294 538954 501914 574398
rect 501294 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 501914 538954
rect 501294 538634 501914 538718
rect 501294 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 501914 538634
rect 501294 502954 501914 538398
rect 501294 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 501914 502954
rect 501294 502634 501914 502718
rect 501294 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 501914 502634
rect 501294 466954 501914 502398
rect 501294 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 501914 466954
rect 501294 466634 501914 466718
rect 501294 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 501914 466634
rect 501294 430954 501914 466398
rect 501294 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 501914 430954
rect 501294 430634 501914 430718
rect 501294 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 501914 430634
rect 501294 394954 501914 430398
rect 501294 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 501914 394954
rect 501294 394634 501914 394718
rect 501294 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 501914 394634
rect 501294 358954 501914 394398
rect 501294 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 501914 358954
rect 501294 358634 501914 358718
rect 501294 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 501914 358634
rect 501294 322954 501914 358398
rect 501294 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 501914 322954
rect 501294 322634 501914 322718
rect 501294 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 501914 322634
rect 501294 286954 501914 322398
rect 501294 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 501914 286954
rect 501294 286634 501914 286718
rect 501294 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 501914 286634
rect 501294 250954 501914 286398
rect 501294 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 501914 250954
rect 501294 250634 501914 250718
rect 501294 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 501914 250634
rect 501294 214954 501914 250398
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 142954 501914 178398
rect 501294 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 501914 142954
rect 501294 142634 501914 142718
rect 501294 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 501914 142634
rect 501294 106954 501914 142398
rect 501294 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 501914 106954
rect 501294 106634 501914 106718
rect 501294 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 501914 106634
rect 501294 70954 501914 106398
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7066 501914 34398
rect 501294 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 501914 -7066
rect 501294 -7386 501914 -7302
rect 501294 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 501914 -7386
rect 501294 -7654 501914 -7622
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 510294 705798 510914 711590
rect 510294 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 510914 705798
rect 510294 705478 510914 705562
rect 510294 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 510914 705478
rect 510294 691954 510914 705242
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 655954 510914 691398
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 619954 510914 655398
rect 510294 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 510914 619954
rect 510294 619634 510914 619718
rect 510294 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 510914 619634
rect 510294 583954 510914 619398
rect 510294 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 510914 583954
rect 510294 583634 510914 583718
rect 510294 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 510914 583634
rect 510294 547954 510914 583398
rect 510294 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 510914 547954
rect 510294 547634 510914 547718
rect 510294 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 510914 547634
rect 510294 511954 510914 547398
rect 510294 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 510914 511954
rect 510294 511634 510914 511718
rect 510294 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 510914 511634
rect 510294 475954 510914 511398
rect 510294 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 510914 475954
rect 510294 475634 510914 475718
rect 510294 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 510914 475634
rect 510294 439954 510914 475398
rect 510294 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 510914 439954
rect 510294 439634 510914 439718
rect 510294 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 510914 439634
rect 510294 403954 510914 439398
rect 510294 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 510914 403954
rect 510294 403634 510914 403718
rect 510294 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 510914 403634
rect 510294 367954 510914 403398
rect 510294 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 510914 367954
rect 510294 367634 510914 367718
rect 510294 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 510914 367634
rect 510294 331954 510914 367398
rect 510294 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 510914 331954
rect 510294 331634 510914 331718
rect 510294 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 510914 331634
rect 510294 295954 510914 331398
rect 510294 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 510914 295954
rect 510294 295634 510914 295718
rect 510294 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 510914 295634
rect 510294 259954 510914 295398
rect 510294 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 510914 259954
rect 510294 259634 510914 259718
rect 510294 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 510914 259634
rect 510294 223954 510914 259398
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 151954 510914 187398
rect 510294 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 510914 151954
rect 510294 151634 510914 151718
rect 510294 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 510914 151634
rect 510294 115954 510914 151398
rect 510294 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 510914 115954
rect 510294 115634 510914 115718
rect 510294 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 510914 115634
rect 510294 79954 510914 115398
rect 510294 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 510914 79954
rect 510294 79634 510914 79718
rect 510294 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 510914 79634
rect 510294 43954 510914 79398
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1306 510914 7398
rect 510294 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 510914 -1306
rect 510294 -1626 510914 -1542
rect 510294 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 510914 -1626
rect 510294 -7654 510914 -1862
rect 514794 706758 515414 711590
rect 514794 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 515414 706758
rect 514794 706438 515414 706522
rect 514794 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 515414 706438
rect 514794 696454 515414 706202
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 624454 515414 659898
rect 514794 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 515414 624454
rect 514794 624134 515414 624218
rect 514794 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 515414 624134
rect 514794 588454 515414 623898
rect 514794 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 515414 588454
rect 514794 588134 515414 588218
rect 514794 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 515414 588134
rect 514794 552454 515414 587898
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 514794 516454 515414 551898
rect 514794 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 515414 516454
rect 514794 516134 515414 516218
rect 514794 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 515414 516134
rect 514794 480454 515414 515898
rect 514794 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 515414 480454
rect 514794 480134 515414 480218
rect 514794 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 515414 480134
rect 514794 444454 515414 479898
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 514794 408454 515414 443898
rect 514794 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 515414 408454
rect 514794 408134 515414 408218
rect 514794 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 515414 408134
rect 514794 372454 515414 407898
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 514794 264454 515414 299898
rect 514794 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 515414 264454
rect 514794 264134 515414 264218
rect 514794 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 515414 264134
rect 514794 228454 515414 263898
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 120454 515414 155898
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 514794 84454 515414 119898
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2266 515414 11898
rect 514794 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 515414 -2266
rect 514794 -2586 515414 -2502
rect 514794 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 515414 -2586
rect 514794 -7654 515414 -2822
rect 519294 707718 519914 711590
rect 519294 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 519914 707718
rect 519294 707398 519914 707482
rect 519294 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 519914 707398
rect 519294 700954 519914 707162
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 628954 519914 664398
rect 519294 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 519914 628954
rect 519294 628634 519914 628718
rect 519294 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 519914 628634
rect 519294 592954 519914 628398
rect 519294 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 519914 592954
rect 519294 592634 519914 592718
rect 519294 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 519914 592634
rect 519294 556954 519914 592398
rect 519294 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 519914 556954
rect 519294 556634 519914 556718
rect 519294 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 519914 556634
rect 519294 520954 519914 556398
rect 519294 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 519914 520954
rect 519294 520634 519914 520718
rect 519294 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 519914 520634
rect 519294 484954 519914 520398
rect 519294 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 519914 484954
rect 519294 484634 519914 484718
rect 519294 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 519914 484634
rect 519294 448954 519914 484398
rect 519294 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 519914 448954
rect 519294 448634 519914 448718
rect 519294 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 519914 448634
rect 519294 412954 519914 448398
rect 519294 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 519914 412954
rect 519294 412634 519914 412718
rect 519294 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 519914 412634
rect 519294 376954 519914 412398
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 268954 519914 304398
rect 519294 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 519914 268954
rect 519294 268634 519914 268718
rect 519294 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 519914 268634
rect 519294 232954 519914 268398
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 124954 519914 160398
rect 519294 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 519914 124954
rect 519294 124634 519914 124718
rect 519294 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 519914 124634
rect 519294 88954 519914 124398
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3226 519914 16398
rect 519294 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 519914 -3226
rect 519294 -3546 519914 -3462
rect 519294 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 519914 -3546
rect 519294 -7654 519914 -3782
rect 523794 708678 524414 711590
rect 523794 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 524414 708678
rect 523794 708358 524414 708442
rect 523794 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 524414 708358
rect 523794 669454 524414 708122
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4186 524414 20898
rect 523794 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 524414 -4186
rect 523794 -4506 524414 -4422
rect 523794 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 524414 -4506
rect 523794 -7654 524414 -4742
rect 528294 709638 528914 711590
rect 528294 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 528914 709638
rect 528294 709318 528914 709402
rect 528294 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 528914 709318
rect 528294 673954 528914 709082
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 528294 565954 528914 601398
rect 528294 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 528914 565954
rect 528294 565634 528914 565718
rect 528294 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 528914 565634
rect 528294 529954 528914 565398
rect 528294 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 528914 529954
rect 528294 529634 528914 529718
rect 528294 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 528914 529634
rect 528294 493954 528914 529398
rect 528294 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 528914 493954
rect 528294 493634 528914 493718
rect 528294 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 528914 493634
rect 528294 457954 528914 493398
rect 528294 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 528914 457954
rect 528294 457634 528914 457718
rect 528294 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 528914 457634
rect 528294 421954 528914 457398
rect 528294 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 528914 421954
rect 528294 421634 528914 421718
rect 528294 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 528914 421634
rect 528294 385954 528914 421398
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 277954 528914 313398
rect 528294 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 528914 277954
rect 528294 277634 528914 277718
rect 528294 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 528914 277634
rect 528294 241954 528914 277398
rect 528294 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 528914 241954
rect 528294 241634 528914 241718
rect 528294 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 528914 241634
rect 528294 205954 528914 241398
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 133954 528914 169398
rect 528294 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 528914 133954
rect 528294 133634 528914 133718
rect 528294 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 528914 133634
rect 528294 97954 528914 133398
rect 528294 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 528914 97954
rect 528294 97634 528914 97718
rect 528294 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 528914 97634
rect 528294 61954 528914 97398
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5146 528914 25398
rect 528294 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 528914 -5146
rect 528294 -5466 528914 -5382
rect 528294 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 528914 -5466
rect 528294 -7654 528914 -5702
rect 532794 710598 533414 711590
rect 532794 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 533414 710598
rect 532794 710278 533414 710362
rect 532794 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 533414 710278
rect 532794 678454 533414 710042
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 570454 533414 605898
rect 532794 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 533414 570454
rect 532794 570134 533414 570218
rect 532794 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 533414 570134
rect 532794 534454 533414 569898
rect 532794 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 533414 534454
rect 532794 534134 533414 534218
rect 532794 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 533414 534134
rect 532794 498454 533414 533898
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 462454 533414 497898
rect 532794 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 533414 462454
rect 532794 462134 533414 462218
rect 532794 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 533414 462134
rect 532794 426454 533414 461898
rect 532794 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 533414 426454
rect 532794 426134 533414 426218
rect 532794 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 533414 426134
rect 532794 390454 533414 425898
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 246454 533414 281898
rect 532794 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 533414 246454
rect 532794 246134 533414 246218
rect 532794 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 533414 246134
rect 532794 210454 533414 245898
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 138454 533414 173898
rect 532794 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 533414 138454
rect 532794 138134 533414 138218
rect 532794 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 533414 138134
rect 532794 102454 533414 137898
rect 532794 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 533414 102454
rect 532794 102134 533414 102218
rect 532794 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 533414 102134
rect 532794 66454 533414 101898
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6106 533414 29898
rect 532794 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 533414 -6106
rect 532794 -6426 533414 -6342
rect 532794 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 533414 -6426
rect 532794 -7654 533414 -6662
rect 537294 711558 537914 711590
rect 537294 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 537914 711558
rect 537294 711238 537914 711322
rect 537294 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 537914 711238
rect 537294 682954 537914 711002
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 537294 574954 537914 610398
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 250954 537914 286398
rect 537294 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 537914 250954
rect 537294 250634 537914 250718
rect 537294 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 537914 250634
rect 537294 214954 537914 250398
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 142954 537914 178398
rect 537294 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 537914 142954
rect 537294 142634 537914 142718
rect 537294 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 537914 142634
rect 537294 106954 537914 142398
rect 537294 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 537914 106954
rect 537294 106634 537914 106718
rect 537294 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 537914 106634
rect 537294 70954 537914 106398
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7066 537914 34398
rect 537294 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 537914 -7066
rect 537294 -7386 537914 -7302
rect 537294 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 537914 -7386
rect 537294 -7654 537914 -7622
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 546294 705798 546914 711590
rect 546294 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 546914 705798
rect 546294 705478 546914 705562
rect 546294 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 546914 705478
rect 546294 691954 546914 705242
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 295954 546914 331398
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 259954 546914 295398
rect 546294 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 546914 259954
rect 546294 259634 546914 259718
rect 546294 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 546914 259634
rect 546294 223954 546914 259398
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1306 546914 7398
rect 546294 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 546914 -1306
rect 546294 -1626 546914 -1542
rect 546294 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 546914 -1626
rect 546294 -7654 546914 -1862
rect 550794 706758 551414 711590
rect 550794 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 551414 706758
rect 550794 706438 551414 706522
rect 550794 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 551414 706438
rect 550794 696454 551414 706202
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 300454 551414 335898
rect 550794 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 551414 300454
rect 550794 300134 551414 300218
rect 550794 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 551414 300134
rect 550794 264454 551414 299898
rect 550794 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 551414 264454
rect 550794 264134 551414 264218
rect 550794 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 551414 264134
rect 550794 228454 551414 263898
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2266 551414 11898
rect 550794 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 551414 -2266
rect 550794 -2586 551414 -2502
rect 550794 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 551414 -2586
rect 550794 -7654 551414 -2822
rect 555294 707718 555914 711590
rect 555294 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 555914 707718
rect 555294 707398 555914 707482
rect 555294 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 555914 707398
rect 555294 700954 555914 707162
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3226 555914 16398
rect 555294 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 555914 -3226
rect 555294 -3546 555914 -3462
rect 555294 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 555914 -3546
rect 555294 -7654 555914 -3782
rect 559794 708678 560414 711590
rect 559794 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 560414 708678
rect 559794 708358 560414 708442
rect 559794 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 560414 708358
rect 559794 669454 560414 708122
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4186 560414 20898
rect 559794 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 560414 -4186
rect 559794 -4506 560414 -4422
rect 559794 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 560414 -4506
rect 559794 -7654 560414 -4742
rect 564294 709638 564914 711590
rect 564294 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 564914 709638
rect 564294 709318 564914 709402
rect 564294 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 564914 709318
rect 564294 673954 564914 709082
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5146 564914 25398
rect 564294 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 564914 -5146
rect 564294 -5466 564914 -5382
rect 564294 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 564914 -5466
rect 564294 -7654 564914 -5702
rect 568794 710598 569414 711590
rect 568794 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 569414 710598
rect 568794 710278 569414 710362
rect 568794 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 569414 710278
rect 568794 678454 569414 710042
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6106 569414 29898
rect 568794 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 569414 -6106
rect 568794 -6426 569414 -6342
rect 568794 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 569414 -6426
rect 568794 -7654 569414 -6662
rect 573294 711558 573914 711590
rect 573294 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 573914 711558
rect 573294 711238 573914 711322
rect 573294 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 573914 711238
rect 573294 682954 573914 711002
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7066 573914 34398
rect 573294 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 573914 -7066
rect 573294 -7386 573914 -7302
rect 573294 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 573914 -7386
rect 573294 -7654 573914 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect 582294 691954 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1306 582914 7398
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691954 586890 705242
rect 586270 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 586890 691954
rect 586270 691634 586890 691718
rect 586270 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 586890 691634
rect 586270 655954 586890 691398
rect 586270 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 586890 655954
rect 586270 655634 586890 655718
rect 586270 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 586890 655634
rect 586270 619954 586890 655398
rect 586270 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 586890 619954
rect 586270 619634 586890 619718
rect 586270 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 586890 619634
rect 586270 583954 586890 619398
rect 586270 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 586890 583954
rect 586270 583634 586890 583718
rect 586270 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 586890 583634
rect 586270 547954 586890 583398
rect 586270 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 586890 547954
rect 586270 547634 586890 547718
rect 586270 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 586890 547634
rect 586270 511954 586890 547398
rect 586270 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 586890 511954
rect 586270 511634 586890 511718
rect 586270 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 586890 511634
rect 586270 475954 586890 511398
rect 586270 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 586890 475954
rect 586270 475634 586890 475718
rect 586270 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 586890 475634
rect 586270 439954 586890 475398
rect 586270 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 586890 439954
rect 586270 439634 586890 439718
rect 586270 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 586890 439634
rect 586270 403954 586890 439398
rect 586270 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 586890 403954
rect 586270 403634 586890 403718
rect 586270 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 586890 403634
rect 586270 367954 586890 403398
rect 586270 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 586890 367954
rect 586270 367634 586890 367718
rect 586270 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 586890 367634
rect 586270 331954 586890 367398
rect 586270 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 586890 331954
rect 586270 331634 586890 331718
rect 586270 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 586890 331634
rect 586270 295954 586890 331398
rect 586270 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 586890 295954
rect 586270 295634 586890 295718
rect 586270 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 586890 295634
rect 586270 259954 586890 295398
rect 586270 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 586890 259954
rect 586270 259634 586890 259718
rect 586270 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 586890 259634
rect 586270 223954 586890 259398
rect 586270 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 586890 223954
rect 586270 223634 586890 223718
rect 586270 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 586890 223634
rect 586270 187954 586890 223398
rect 586270 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 586890 187954
rect 586270 187634 586890 187718
rect 586270 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 586890 187634
rect 586270 151954 586890 187398
rect 586270 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 586890 151954
rect 586270 151634 586890 151718
rect 586270 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 586890 151634
rect 586270 115954 586890 151398
rect 586270 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 586890 115954
rect 586270 115634 586890 115718
rect 586270 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 586890 115634
rect 586270 79954 586890 115398
rect 586270 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 586890 79954
rect 586270 79634 586890 79718
rect 586270 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 586890 79634
rect 586270 43954 586890 79398
rect 586270 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 586890 43954
rect 586270 43634 586890 43718
rect 586270 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 586890 43634
rect 586270 7954 586890 43398
rect 586270 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 586890 7954
rect 586270 7634 586890 7718
rect 586270 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 586890 7634
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 7398
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 696454 587850 706202
rect 587230 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 587850 696454
rect 587230 696134 587850 696218
rect 587230 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 587850 696134
rect 587230 660454 587850 695898
rect 587230 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 587850 660454
rect 587230 660134 587850 660218
rect 587230 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 587850 660134
rect 587230 624454 587850 659898
rect 587230 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 587850 624454
rect 587230 624134 587850 624218
rect 587230 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 587850 624134
rect 587230 588454 587850 623898
rect 587230 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 587850 588454
rect 587230 588134 587850 588218
rect 587230 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 587850 588134
rect 587230 552454 587850 587898
rect 587230 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 587850 552454
rect 587230 552134 587850 552218
rect 587230 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 587850 552134
rect 587230 516454 587850 551898
rect 587230 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 587850 516454
rect 587230 516134 587850 516218
rect 587230 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 587850 516134
rect 587230 480454 587850 515898
rect 587230 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 587850 480454
rect 587230 480134 587850 480218
rect 587230 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 587850 480134
rect 587230 444454 587850 479898
rect 587230 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 587850 444454
rect 587230 444134 587850 444218
rect 587230 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 587850 444134
rect 587230 408454 587850 443898
rect 587230 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 587850 408454
rect 587230 408134 587850 408218
rect 587230 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 587850 408134
rect 587230 372454 587850 407898
rect 587230 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 587850 372454
rect 587230 372134 587850 372218
rect 587230 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 587850 372134
rect 587230 336454 587850 371898
rect 587230 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 587850 336454
rect 587230 336134 587850 336218
rect 587230 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 587850 336134
rect 587230 300454 587850 335898
rect 587230 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 587850 300454
rect 587230 300134 587850 300218
rect 587230 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 587850 300134
rect 587230 264454 587850 299898
rect 587230 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 587850 264454
rect 587230 264134 587850 264218
rect 587230 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 587850 264134
rect 587230 228454 587850 263898
rect 587230 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 587850 228454
rect 587230 228134 587850 228218
rect 587230 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 587850 228134
rect 587230 192454 587850 227898
rect 587230 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 587850 192454
rect 587230 192134 587850 192218
rect 587230 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 587850 192134
rect 587230 156454 587850 191898
rect 587230 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 587850 156454
rect 587230 156134 587850 156218
rect 587230 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 587850 156134
rect 587230 120454 587850 155898
rect 587230 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 587850 120454
rect 587230 120134 587850 120218
rect 587230 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 587850 120134
rect 587230 84454 587850 119898
rect 587230 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 587850 84454
rect 587230 84134 587850 84218
rect 587230 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 587850 84134
rect 587230 48454 587850 83898
rect 587230 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 587850 48454
rect 587230 48134 587850 48218
rect 587230 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 587850 48134
rect 587230 12454 587850 47898
rect 587230 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 587850 12454
rect 587230 12134 587850 12218
rect 587230 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 587850 12134
rect 587230 -2266 587850 11898
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 700954 588810 707162
rect 588190 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 588810 700954
rect 588190 700634 588810 700718
rect 588190 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 588810 700634
rect 588190 664954 588810 700398
rect 588190 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 588810 664954
rect 588190 664634 588810 664718
rect 588190 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 588810 664634
rect 588190 628954 588810 664398
rect 588190 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 588810 628954
rect 588190 628634 588810 628718
rect 588190 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 588810 628634
rect 588190 592954 588810 628398
rect 588190 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 588810 592954
rect 588190 592634 588810 592718
rect 588190 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 588810 592634
rect 588190 556954 588810 592398
rect 588190 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect 588190 556634 588810 556718
rect 588190 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 588810 556634
rect 588190 520954 588810 556398
rect 588190 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 588810 520954
rect 588190 520634 588810 520718
rect 588190 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 588810 520634
rect 588190 484954 588810 520398
rect 588190 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 588810 484954
rect 588190 484634 588810 484718
rect 588190 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 588810 484634
rect 588190 448954 588810 484398
rect 588190 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 588810 448954
rect 588190 448634 588810 448718
rect 588190 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 588810 448634
rect 588190 412954 588810 448398
rect 588190 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 588810 412954
rect 588190 412634 588810 412718
rect 588190 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 588810 412634
rect 588190 376954 588810 412398
rect 588190 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect 588190 376634 588810 376718
rect 588190 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 588810 376634
rect 588190 340954 588810 376398
rect 588190 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 588810 340954
rect 588190 340634 588810 340718
rect 588190 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 588810 340634
rect 588190 304954 588810 340398
rect 588190 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 588810 304954
rect 588190 304634 588810 304718
rect 588190 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 588810 304634
rect 588190 268954 588810 304398
rect 588190 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 588810 268954
rect 588190 268634 588810 268718
rect 588190 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 588810 268634
rect 588190 232954 588810 268398
rect 588190 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 588810 232954
rect 588190 232634 588810 232718
rect 588190 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 588810 232634
rect 588190 196954 588810 232398
rect 588190 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect 588190 196634 588810 196718
rect 588190 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 588810 196634
rect 588190 160954 588810 196398
rect 588190 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 588810 160954
rect 588190 160634 588810 160718
rect 588190 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 588810 160634
rect 588190 124954 588810 160398
rect 588190 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 588810 124954
rect 588190 124634 588810 124718
rect 588190 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 588810 124634
rect 588190 88954 588810 124398
rect 588190 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 588810 88954
rect 588190 88634 588810 88718
rect 588190 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 588810 88634
rect 588190 52954 588810 88398
rect 588190 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 588810 52954
rect 588190 52634 588810 52718
rect 588190 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 588810 52634
rect 588190 16954 588810 52398
rect 588190 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect 588190 16634 588810 16718
rect 588190 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 588810 16634
rect 588190 -3226 588810 16398
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 669454 589770 708122
rect 589150 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 589770 669454
rect 589150 669134 589770 669218
rect 589150 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 589770 669134
rect 589150 633454 589770 668898
rect 589150 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 589770 633454
rect 589150 633134 589770 633218
rect 589150 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 589770 633134
rect 589150 597454 589770 632898
rect 589150 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 589770 597454
rect 589150 597134 589770 597218
rect 589150 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 589770 597134
rect 589150 561454 589770 596898
rect 589150 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 589770 561454
rect 589150 561134 589770 561218
rect 589150 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 589770 561134
rect 589150 525454 589770 560898
rect 589150 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 589770 525454
rect 589150 525134 589770 525218
rect 589150 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 589770 525134
rect 589150 489454 589770 524898
rect 589150 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 589770 489454
rect 589150 489134 589770 489218
rect 589150 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 589770 489134
rect 589150 453454 589770 488898
rect 589150 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 589770 453454
rect 589150 453134 589770 453218
rect 589150 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 589770 453134
rect 589150 417454 589770 452898
rect 589150 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 589770 417454
rect 589150 417134 589770 417218
rect 589150 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 589770 417134
rect 589150 381454 589770 416898
rect 589150 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 589770 381454
rect 589150 381134 589770 381218
rect 589150 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 589770 381134
rect 589150 345454 589770 380898
rect 589150 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 589770 345454
rect 589150 345134 589770 345218
rect 589150 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 589770 345134
rect 589150 309454 589770 344898
rect 589150 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 589770 309454
rect 589150 309134 589770 309218
rect 589150 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 589770 309134
rect 589150 273454 589770 308898
rect 589150 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 589770 273454
rect 589150 273134 589770 273218
rect 589150 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 589770 273134
rect 589150 237454 589770 272898
rect 589150 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 589770 237454
rect 589150 237134 589770 237218
rect 589150 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 589770 237134
rect 589150 201454 589770 236898
rect 589150 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 589770 201454
rect 589150 201134 589770 201218
rect 589150 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 589770 201134
rect 589150 165454 589770 200898
rect 589150 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 589770 165454
rect 589150 165134 589770 165218
rect 589150 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 589770 165134
rect 589150 129454 589770 164898
rect 589150 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 589770 129454
rect 589150 129134 589770 129218
rect 589150 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 589770 129134
rect 589150 93454 589770 128898
rect 589150 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 589770 93454
rect 589150 93134 589770 93218
rect 589150 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 589770 93134
rect 589150 57454 589770 92898
rect 589150 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 589770 57454
rect 589150 57134 589770 57218
rect 589150 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 589770 57134
rect 589150 21454 589770 56898
rect 589150 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 589770 21454
rect 589150 21134 589770 21218
rect 589150 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 589770 21134
rect 589150 -4186 589770 20898
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 673954 590730 709082
rect 590110 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 590730 673954
rect 590110 673634 590730 673718
rect 590110 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 590730 673634
rect 590110 637954 590730 673398
rect 590110 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 590730 637954
rect 590110 637634 590730 637718
rect 590110 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 590730 637634
rect 590110 601954 590730 637398
rect 590110 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 590730 601954
rect 590110 601634 590730 601718
rect 590110 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 590730 601634
rect 590110 565954 590730 601398
rect 590110 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 590730 565954
rect 590110 565634 590730 565718
rect 590110 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 590730 565634
rect 590110 529954 590730 565398
rect 590110 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 590730 529954
rect 590110 529634 590730 529718
rect 590110 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 590730 529634
rect 590110 493954 590730 529398
rect 590110 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 590730 493954
rect 590110 493634 590730 493718
rect 590110 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 590730 493634
rect 590110 457954 590730 493398
rect 590110 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 590730 457954
rect 590110 457634 590730 457718
rect 590110 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 590730 457634
rect 590110 421954 590730 457398
rect 590110 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 590730 421954
rect 590110 421634 590730 421718
rect 590110 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 590730 421634
rect 590110 385954 590730 421398
rect 590110 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 590730 385954
rect 590110 385634 590730 385718
rect 590110 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 590730 385634
rect 590110 349954 590730 385398
rect 590110 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 590730 349954
rect 590110 349634 590730 349718
rect 590110 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 590730 349634
rect 590110 313954 590730 349398
rect 590110 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 590730 313954
rect 590110 313634 590730 313718
rect 590110 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 590730 313634
rect 590110 277954 590730 313398
rect 590110 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 590730 277954
rect 590110 277634 590730 277718
rect 590110 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 590730 277634
rect 590110 241954 590730 277398
rect 590110 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 590730 241954
rect 590110 241634 590730 241718
rect 590110 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 590730 241634
rect 590110 205954 590730 241398
rect 590110 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 590730 205954
rect 590110 205634 590730 205718
rect 590110 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 590730 205634
rect 590110 169954 590730 205398
rect 590110 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 590730 169954
rect 590110 169634 590730 169718
rect 590110 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 590730 169634
rect 590110 133954 590730 169398
rect 590110 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 590730 133954
rect 590110 133634 590730 133718
rect 590110 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 590730 133634
rect 590110 97954 590730 133398
rect 590110 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 590730 97954
rect 590110 97634 590730 97718
rect 590110 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 590730 97634
rect 590110 61954 590730 97398
rect 590110 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 590730 61954
rect 590110 61634 590730 61718
rect 590110 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 590730 61634
rect 590110 25954 590730 61398
rect 590110 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 590730 25954
rect 590110 25634 590730 25718
rect 590110 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 590730 25634
rect 590110 -5146 590730 25398
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 678454 591690 710042
rect 591070 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 591690 678454
rect 591070 678134 591690 678218
rect 591070 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 591690 678134
rect 591070 642454 591690 677898
rect 591070 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 591690 642454
rect 591070 642134 591690 642218
rect 591070 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 591690 642134
rect 591070 606454 591690 641898
rect 591070 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 591690 606454
rect 591070 606134 591690 606218
rect 591070 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 591690 606134
rect 591070 570454 591690 605898
rect 591070 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 591690 570454
rect 591070 570134 591690 570218
rect 591070 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 591690 570134
rect 591070 534454 591690 569898
rect 591070 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 591690 534454
rect 591070 534134 591690 534218
rect 591070 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 591690 534134
rect 591070 498454 591690 533898
rect 591070 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 591690 498454
rect 591070 498134 591690 498218
rect 591070 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 591690 498134
rect 591070 462454 591690 497898
rect 591070 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 591690 462454
rect 591070 462134 591690 462218
rect 591070 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 591690 462134
rect 591070 426454 591690 461898
rect 591070 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 591690 426454
rect 591070 426134 591690 426218
rect 591070 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 591690 426134
rect 591070 390454 591690 425898
rect 591070 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 591690 390454
rect 591070 390134 591690 390218
rect 591070 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 591690 390134
rect 591070 354454 591690 389898
rect 591070 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 591690 354454
rect 591070 354134 591690 354218
rect 591070 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 591690 354134
rect 591070 318454 591690 353898
rect 591070 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 591690 318454
rect 591070 318134 591690 318218
rect 591070 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 591690 318134
rect 591070 282454 591690 317898
rect 591070 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 591690 282454
rect 591070 282134 591690 282218
rect 591070 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 591690 282134
rect 591070 246454 591690 281898
rect 591070 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 591690 246454
rect 591070 246134 591690 246218
rect 591070 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 591690 246134
rect 591070 210454 591690 245898
rect 591070 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 591690 210454
rect 591070 210134 591690 210218
rect 591070 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 591690 210134
rect 591070 174454 591690 209898
rect 591070 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 591690 174454
rect 591070 174134 591690 174218
rect 591070 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 591690 174134
rect 591070 138454 591690 173898
rect 591070 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 591690 138454
rect 591070 138134 591690 138218
rect 591070 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 591690 138134
rect 591070 102454 591690 137898
rect 591070 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 591690 102454
rect 591070 102134 591690 102218
rect 591070 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 591690 102134
rect 591070 66454 591690 101898
rect 591070 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 591690 66454
rect 591070 66134 591690 66218
rect 591070 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 591690 66134
rect 591070 30454 591690 65898
rect 591070 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 591690 30454
rect 591070 30134 591690 30218
rect 591070 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 591690 30134
rect 591070 -6106 591690 29898
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 682954 592650 711002
rect 592030 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect 592030 682634 592650 682718
rect 592030 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect 592030 646954 592650 682398
rect 592030 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect 592030 646634 592650 646718
rect 592030 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect 592030 610954 592650 646398
rect 592030 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect 592030 610634 592650 610718
rect 592030 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect 592030 574954 592650 610398
rect 592030 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect 592030 574634 592650 574718
rect 592030 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect 592030 538954 592650 574398
rect 592030 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect 592030 538634 592650 538718
rect 592030 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect 592030 502954 592650 538398
rect 592030 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect 592030 502634 592650 502718
rect 592030 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect 592030 466954 592650 502398
rect 592030 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect 592030 466634 592650 466718
rect 592030 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect 592030 430954 592650 466398
rect 592030 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect 592030 430634 592650 430718
rect 592030 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect 592030 394954 592650 430398
rect 592030 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect 592030 394634 592650 394718
rect 592030 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect 592030 358954 592650 394398
rect 592030 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect 592030 358634 592650 358718
rect 592030 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect 592030 322954 592650 358398
rect 592030 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect 592030 322634 592650 322718
rect 592030 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect 592030 286954 592650 322398
rect 592030 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect 592030 286634 592650 286718
rect 592030 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect 592030 250954 592650 286398
rect 592030 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect 592030 250634 592650 250718
rect 592030 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect 592030 214954 592650 250398
rect 592030 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect 592030 214634 592650 214718
rect 592030 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect 592030 178954 592650 214398
rect 592030 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect 592030 178634 592650 178718
rect 592030 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect 592030 142954 592650 178398
rect 592030 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect 592030 142634 592650 142718
rect 592030 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect 592030 106954 592650 142398
rect 592030 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect 592030 106634 592650 106718
rect 592030 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect 592030 70954 592650 106398
rect 592030 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect 592030 70634 592650 70718
rect 592030 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect 592030 34954 592650 70398
rect 592030 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect 592030 34634 592650 34718
rect 592030 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect 592030 -7066 592650 34398
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 682718 -8458 682954
rect -8374 682718 -8138 682954
rect -8694 682398 -8458 682634
rect -8374 682398 -8138 682634
rect -8694 646718 -8458 646954
rect -8374 646718 -8138 646954
rect -8694 646398 -8458 646634
rect -8374 646398 -8138 646634
rect -8694 610718 -8458 610954
rect -8374 610718 -8138 610954
rect -8694 610398 -8458 610634
rect -8374 610398 -8138 610634
rect -8694 574718 -8458 574954
rect -8374 574718 -8138 574954
rect -8694 574398 -8458 574634
rect -8374 574398 -8138 574634
rect -8694 538718 -8458 538954
rect -8374 538718 -8138 538954
rect -8694 538398 -8458 538634
rect -8374 538398 -8138 538634
rect -8694 502718 -8458 502954
rect -8374 502718 -8138 502954
rect -8694 502398 -8458 502634
rect -8374 502398 -8138 502634
rect -8694 466718 -8458 466954
rect -8374 466718 -8138 466954
rect -8694 466398 -8458 466634
rect -8374 466398 -8138 466634
rect -8694 430718 -8458 430954
rect -8374 430718 -8138 430954
rect -8694 430398 -8458 430634
rect -8374 430398 -8138 430634
rect -8694 394718 -8458 394954
rect -8374 394718 -8138 394954
rect -8694 394398 -8458 394634
rect -8374 394398 -8138 394634
rect -8694 358718 -8458 358954
rect -8374 358718 -8138 358954
rect -8694 358398 -8458 358634
rect -8374 358398 -8138 358634
rect -8694 322718 -8458 322954
rect -8374 322718 -8138 322954
rect -8694 322398 -8458 322634
rect -8374 322398 -8138 322634
rect -8694 286718 -8458 286954
rect -8374 286718 -8138 286954
rect -8694 286398 -8458 286634
rect -8374 286398 -8138 286634
rect -8694 250718 -8458 250954
rect -8374 250718 -8138 250954
rect -8694 250398 -8458 250634
rect -8374 250398 -8138 250634
rect -8694 214718 -8458 214954
rect -8374 214718 -8138 214954
rect -8694 214398 -8458 214634
rect -8374 214398 -8138 214634
rect -8694 178718 -8458 178954
rect -8374 178718 -8138 178954
rect -8694 178398 -8458 178634
rect -8374 178398 -8138 178634
rect -8694 142718 -8458 142954
rect -8374 142718 -8138 142954
rect -8694 142398 -8458 142634
rect -8374 142398 -8138 142634
rect -8694 106718 -8458 106954
rect -8374 106718 -8138 106954
rect -8694 106398 -8458 106634
rect -8374 106398 -8138 106634
rect -8694 70718 -8458 70954
rect -8374 70718 -8138 70954
rect -8694 70398 -8458 70634
rect -8374 70398 -8138 70634
rect -8694 34718 -8458 34954
rect -8374 34718 -8138 34954
rect -8694 34398 -8458 34634
rect -8374 34398 -8138 34634
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 678218 -7498 678454
rect -7414 678218 -7178 678454
rect -7734 677898 -7498 678134
rect -7414 677898 -7178 678134
rect -7734 642218 -7498 642454
rect -7414 642218 -7178 642454
rect -7734 641898 -7498 642134
rect -7414 641898 -7178 642134
rect -7734 606218 -7498 606454
rect -7414 606218 -7178 606454
rect -7734 605898 -7498 606134
rect -7414 605898 -7178 606134
rect -7734 570218 -7498 570454
rect -7414 570218 -7178 570454
rect -7734 569898 -7498 570134
rect -7414 569898 -7178 570134
rect -7734 534218 -7498 534454
rect -7414 534218 -7178 534454
rect -7734 533898 -7498 534134
rect -7414 533898 -7178 534134
rect -7734 498218 -7498 498454
rect -7414 498218 -7178 498454
rect -7734 497898 -7498 498134
rect -7414 497898 -7178 498134
rect -7734 462218 -7498 462454
rect -7414 462218 -7178 462454
rect -7734 461898 -7498 462134
rect -7414 461898 -7178 462134
rect -7734 426218 -7498 426454
rect -7414 426218 -7178 426454
rect -7734 425898 -7498 426134
rect -7414 425898 -7178 426134
rect -7734 390218 -7498 390454
rect -7414 390218 -7178 390454
rect -7734 389898 -7498 390134
rect -7414 389898 -7178 390134
rect -7734 354218 -7498 354454
rect -7414 354218 -7178 354454
rect -7734 353898 -7498 354134
rect -7414 353898 -7178 354134
rect -7734 318218 -7498 318454
rect -7414 318218 -7178 318454
rect -7734 317898 -7498 318134
rect -7414 317898 -7178 318134
rect -7734 282218 -7498 282454
rect -7414 282218 -7178 282454
rect -7734 281898 -7498 282134
rect -7414 281898 -7178 282134
rect -7734 246218 -7498 246454
rect -7414 246218 -7178 246454
rect -7734 245898 -7498 246134
rect -7414 245898 -7178 246134
rect -7734 210218 -7498 210454
rect -7414 210218 -7178 210454
rect -7734 209898 -7498 210134
rect -7414 209898 -7178 210134
rect -7734 174218 -7498 174454
rect -7414 174218 -7178 174454
rect -7734 173898 -7498 174134
rect -7414 173898 -7178 174134
rect -7734 138218 -7498 138454
rect -7414 138218 -7178 138454
rect -7734 137898 -7498 138134
rect -7414 137898 -7178 138134
rect -7734 102218 -7498 102454
rect -7414 102218 -7178 102454
rect -7734 101898 -7498 102134
rect -7414 101898 -7178 102134
rect -7734 66218 -7498 66454
rect -7414 66218 -7178 66454
rect -7734 65898 -7498 66134
rect -7414 65898 -7178 66134
rect -7734 30218 -7498 30454
rect -7414 30218 -7178 30454
rect -7734 29898 -7498 30134
rect -7414 29898 -7178 30134
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 673718 -6538 673954
rect -6454 673718 -6218 673954
rect -6774 673398 -6538 673634
rect -6454 673398 -6218 673634
rect -6774 637718 -6538 637954
rect -6454 637718 -6218 637954
rect -6774 637398 -6538 637634
rect -6454 637398 -6218 637634
rect -6774 601718 -6538 601954
rect -6454 601718 -6218 601954
rect -6774 601398 -6538 601634
rect -6454 601398 -6218 601634
rect -6774 565718 -6538 565954
rect -6454 565718 -6218 565954
rect -6774 565398 -6538 565634
rect -6454 565398 -6218 565634
rect -6774 529718 -6538 529954
rect -6454 529718 -6218 529954
rect -6774 529398 -6538 529634
rect -6454 529398 -6218 529634
rect -6774 493718 -6538 493954
rect -6454 493718 -6218 493954
rect -6774 493398 -6538 493634
rect -6454 493398 -6218 493634
rect -6774 457718 -6538 457954
rect -6454 457718 -6218 457954
rect -6774 457398 -6538 457634
rect -6454 457398 -6218 457634
rect -6774 421718 -6538 421954
rect -6454 421718 -6218 421954
rect -6774 421398 -6538 421634
rect -6454 421398 -6218 421634
rect -6774 385718 -6538 385954
rect -6454 385718 -6218 385954
rect -6774 385398 -6538 385634
rect -6454 385398 -6218 385634
rect -6774 349718 -6538 349954
rect -6454 349718 -6218 349954
rect -6774 349398 -6538 349634
rect -6454 349398 -6218 349634
rect -6774 313718 -6538 313954
rect -6454 313718 -6218 313954
rect -6774 313398 -6538 313634
rect -6454 313398 -6218 313634
rect -6774 277718 -6538 277954
rect -6454 277718 -6218 277954
rect -6774 277398 -6538 277634
rect -6454 277398 -6218 277634
rect -6774 241718 -6538 241954
rect -6454 241718 -6218 241954
rect -6774 241398 -6538 241634
rect -6454 241398 -6218 241634
rect -6774 205718 -6538 205954
rect -6454 205718 -6218 205954
rect -6774 205398 -6538 205634
rect -6454 205398 -6218 205634
rect -6774 169718 -6538 169954
rect -6454 169718 -6218 169954
rect -6774 169398 -6538 169634
rect -6454 169398 -6218 169634
rect -6774 133718 -6538 133954
rect -6454 133718 -6218 133954
rect -6774 133398 -6538 133634
rect -6454 133398 -6218 133634
rect -6774 97718 -6538 97954
rect -6454 97718 -6218 97954
rect -6774 97398 -6538 97634
rect -6454 97398 -6218 97634
rect -6774 61718 -6538 61954
rect -6454 61718 -6218 61954
rect -6774 61398 -6538 61634
rect -6454 61398 -6218 61634
rect -6774 25718 -6538 25954
rect -6454 25718 -6218 25954
rect -6774 25398 -6538 25634
rect -6454 25398 -6218 25634
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 669218 -5578 669454
rect -5494 669218 -5258 669454
rect -5814 668898 -5578 669134
rect -5494 668898 -5258 669134
rect -5814 633218 -5578 633454
rect -5494 633218 -5258 633454
rect -5814 632898 -5578 633134
rect -5494 632898 -5258 633134
rect -5814 597218 -5578 597454
rect -5494 597218 -5258 597454
rect -5814 596898 -5578 597134
rect -5494 596898 -5258 597134
rect -5814 561218 -5578 561454
rect -5494 561218 -5258 561454
rect -5814 560898 -5578 561134
rect -5494 560898 -5258 561134
rect -5814 525218 -5578 525454
rect -5494 525218 -5258 525454
rect -5814 524898 -5578 525134
rect -5494 524898 -5258 525134
rect -5814 489218 -5578 489454
rect -5494 489218 -5258 489454
rect -5814 488898 -5578 489134
rect -5494 488898 -5258 489134
rect -5814 453218 -5578 453454
rect -5494 453218 -5258 453454
rect -5814 452898 -5578 453134
rect -5494 452898 -5258 453134
rect -5814 417218 -5578 417454
rect -5494 417218 -5258 417454
rect -5814 416898 -5578 417134
rect -5494 416898 -5258 417134
rect -5814 381218 -5578 381454
rect -5494 381218 -5258 381454
rect -5814 380898 -5578 381134
rect -5494 380898 -5258 381134
rect -5814 345218 -5578 345454
rect -5494 345218 -5258 345454
rect -5814 344898 -5578 345134
rect -5494 344898 -5258 345134
rect -5814 309218 -5578 309454
rect -5494 309218 -5258 309454
rect -5814 308898 -5578 309134
rect -5494 308898 -5258 309134
rect -5814 273218 -5578 273454
rect -5494 273218 -5258 273454
rect -5814 272898 -5578 273134
rect -5494 272898 -5258 273134
rect -5814 237218 -5578 237454
rect -5494 237218 -5258 237454
rect -5814 236898 -5578 237134
rect -5494 236898 -5258 237134
rect -5814 201218 -5578 201454
rect -5494 201218 -5258 201454
rect -5814 200898 -5578 201134
rect -5494 200898 -5258 201134
rect -5814 165218 -5578 165454
rect -5494 165218 -5258 165454
rect -5814 164898 -5578 165134
rect -5494 164898 -5258 165134
rect -5814 129218 -5578 129454
rect -5494 129218 -5258 129454
rect -5814 128898 -5578 129134
rect -5494 128898 -5258 129134
rect -5814 93218 -5578 93454
rect -5494 93218 -5258 93454
rect -5814 92898 -5578 93134
rect -5494 92898 -5258 93134
rect -5814 57218 -5578 57454
rect -5494 57218 -5258 57454
rect -5814 56898 -5578 57134
rect -5494 56898 -5258 57134
rect -5814 21218 -5578 21454
rect -5494 21218 -5258 21454
rect -5814 20898 -5578 21134
rect -5494 20898 -5258 21134
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 700718 -4618 700954
rect -4534 700718 -4298 700954
rect -4854 700398 -4618 700634
rect -4534 700398 -4298 700634
rect -4854 664718 -4618 664954
rect -4534 664718 -4298 664954
rect -4854 664398 -4618 664634
rect -4534 664398 -4298 664634
rect -4854 628718 -4618 628954
rect -4534 628718 -4298 628954
rect -4854 628398 -4618 628634
rect -4534 628398 -4298 628634
rect -4854 592718 -4618 592954
rect -4534 592718 -4298 592954
rect -4854 592398 -4618 592634
rect -4534 592398 -4298 592634
rect -4854 556718 -4618 556954
rect -4534 556718 -4298 556954
rect -4854 556398 -4618 556634
rect -4534 556398 -4298 556634
rect -4854 520718 -4618 520954
rect -4534 520718 -4298 520954
rect -4854 520398 -4618 520634
rect -4534 520398 -4298 520634
rect -4854 484718 -4618 484954
rect -4534 484718 -4298 484954
rect -4854 484398 -4618 484634
rect -4534 484398 -4298 484634
rect -4854 448718 -4618 448954
rect -4534 448718 -4298 448954
rect -4854 448398 -4618 448634
rect -4534 448398 -4298 448634
rect -4854 412718 -4618 412954
rect -4534 412718 -4298 412954
rect -4854 412398 -4618 412634
rect -4534 412398 -4298 412634
rect -4854 376718 -4618 376954
rect -4534 376718 -4298 376954
rect -4854 376398 -4618 376634
rect -4534 376398 -4298 376634
rect -4854 340718 -4618 340954
rect -4534 340718 -4298 340954
rect -4854 340398 -4618 340634
rect -4534 340398 -4298 340634
rect -4854 304718 -4618 304954
rect -4534 304718 -4298 304954
rect -4854 304398 -4618 304634
rect -4534 304398 -4298 304634
rect -4854 268718 -4618 268954
rect -4534 268718 -4298 268954
rect -4854 268398 -4618 268634
rect -4534 268398 -4298 268634
rect -4854 232718 -4618 232954
rect -4534 232718 -4298 232954
rect -4854 232398 -4618 232634
rect -4534 232398 -4298 232634
rect -4854 196718 -4618 196954
rect -4534 196718 -4298 196954
rect -4854 196398 -4618 196634
rect -4534 196398 -4298 196634
rect -4854 160718 -4618 160954
rect -4534 160718 -4298 160954
rect -4854 160398 -4618 160634
rect -4534 160398 -4298 160634
rect -4854 124718 -4618 124954
rect -4534 124718 -4298 124954
rect -4854 124398 -4618 124634
rect -4534 124398 -4298 124634
rect -4854 88718 -4618 88954
rect -4534 88718 -4298 88954
rect -4854 88398 -4618 88634
rect -4534 88398 -4298 88634
rect -4854 52718 -4618 52954
rect -4534 52718 -4298 52954
rect -4854 52398 -4618 52634
rect -4534 52398 -4298 52634
rect -4854 16718 -4618 16954
rect -4534 16718 -4298 16954
rect -4854 16398 -4618 16634
rect -4534 16398 -4298 16634
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 696218 -3658 696454
rect -3574 696218 -3338 696454
rect -3894 695898 -3658 696134
rect -3574 695898 -3338 696134
rect -3894 660218 -3658 660454
rect -3574 660218 -3338 660454
rect -3894 659898 -3658 660134
rect -3574 659898 -3338 660134
rect -3894 624218 -3658 624454
rect -3574 624218 -3338 624454
rect -3894 623898 -3658 624134
rect -3574 623898 -3338 624134
rect -3894 588218 -3658 588454
rect -3574 588218 -3338 588454
rect -3894 587898 -3658 588134
rect -3574 587898 -3338 588134
rect -3894 552218 -3658 552454
rect -3574 552218 -3338 552454
rect -3894 551898 -3658 552134
rect -3574 551898 -3338 552134
rect -3894 516218 -3658 516454
rect -3574 516218 -3338 516454
rect -3894 515898 -3658 516134
rect -3574 515898 -3338 516134
rect -3894 480218 -3658 480454
rect -3574 480218 -3338 480454
rect -3894 479898 -3658 480134
rect -3574 479898 -3338 480134
rect -3894 444218 -3658 444454
rect -3574 444218 -3338 444454
rect -3894 443898 -3658 444134
rect -3574 443898 -3338 444134
rect -3894 408218 -3658 408454
rect -3574 408218 -3338 408454
rect -3894 407898 -3658 408134
rect -3574 407898 -3338 408134
rect -3894 372218 -3658 372454
rect -3574 372218 -3338 372454
rect -3894 371898 -3658 372134
rect -3574 371898 -3338 372134
rect -3894 336218 -3658 336454
rect -3574 336218 -3338 336454
rect -3894 335898 -3658 336134
rect -3574 335898 -3338 336134
rect -3894 300218 -3658 300454
rect -3574 300218 -3338 300454
rect -3894 299898 -3658 300134
rect -3574 299898 -3338 300134
rect -3894 264218 -3658 264454
rect -3574 264218 -3338 264454
rect -3894 263898 -3658 264134
rect -3574 263898 -3338 264134
rect -3894 228218 -3658 228454
rect -3574 228218 -3338 228454
rect -3894 227898 -3658 228134
rect -3574 227898 -3338 228134
rect -3894 192218 -3658 192454
rect -3574 192218 -3338 192454
rect -3894 191898 -3658 192134
rect -3574 191898 -3338 192134
rect -3894 156218 -3658 156454
rect -3574 156218 -3338 156454
rect -3894 155898 -3658 156134
rect -3574 155898 -3338 156134
rect -3894 120218 -3658 120454
rect -3574 120218 -3338 120454
rect -3894 119898 -3658 120134
rect -3574 119898 -3338 120134
rect -3894 84218 -3658 84454
rect -3574 84218 -3338 84454
rect -3894 83898 -3658 84134
rect -3574 83898 -3338 84134
rect -3894 48218 -3658 48454
rect -3574 48218 -3338 48454
rect -3894 47898 -3658 48134
rect -3574 47898 -3338 48134
rect -3894 12218 -3658 12454
rect -3574 12218 -3338 12454
rect -3894 11898 -3658 12134
rect -3574 11898 -3338 12134
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 691718 -2698 691954
rect -2614 691718 -2378 691954
rect -2934 691398 -2698 691634
rect -2614 691398 -2378 691634
rect -2934 655718 -2698 655954
rect -2614 655718 -2378 655954
rect -2934 655398 -2698 655634
rect -2614 655398 -2378 655634
rect -2934 619718 -2698 619954
rect -2614 619718 -2378 619954
rect -2934 619398 -2698 619634
rect -2614 619398 -2378 619634
rect -2934 583718 -2698 583954
rect -2614 583718 -2378 583954
rect -2934 583398 -2698 583634
rect -2614 583398 -2378 583634
rect -2934 547718 -2698 547954
rect -2614 547718 -2378 547954
rect -2934 547398 -2698 547634
rect -2614 547398 -2378 547634
rect -2934 511718 -2698 511954
rect -2614 511718 -2378 511954
rect -2934 511398 -2698 511634
rect -2614 511398 -2378 511634
rect -2934 475718 -2698 475954
rect -2614 475718 -2378 475954
rect -2934 475398 -2698 475634
rect -2614 475398 -2378 475634
rect -2934 439718 -2698 439954
rect -2614 439718 -2378 439954
rect -2934 439398 -2698 439634
rect -2614 439398 -2378 439634
rect -2934 403718 -2698 403954
rect -2614 403718 -2378 403954
rect -2934 403398 -2698 403634
rect -2614 403398 -2378 403634
rect -2934 367718 -2698 367954
rect -2614 367718 -2378 367954
rect -2934 367398 -2698 367634
rect -2614 367398 -2378 367634
rect -2934 331718 -2698 331954
rect -2614 331718 -2378 331954
rect -2934 331398 -2698 331634
rect -2614 331398 -2378 331634
rect -2934 295718 -2698 295954
rect -2614 295718 -2378 295954
rect -2934 295398 -2698 295634
rect -2614 295398 -2378 295634
rect -2934 259718 -2698 259954
rect -2614 259718 -2378 259954
rect -2934 259398 -2698 259634
rect -2614 259398 -2378 259634
rect -2934 223718 -2698 223954
rect -2614 223718 -2378 223954
rect -2934 223398 -2698 223634
rect -2614 223398 -2378 223634
rect -2934 187718 -2698 187954
rect -2614 187718 -2378 187954
rect -2934 187398 -2698 187634
rect -2614 187398 -2378 187634
rect -2934 151718 -2698 151954
rect -2614 151718 -2378 151954
rect -2934 151398 -2698 151634
rect -2614 151398 -2378 151634
rect -2934 115718 -2698 115954
rect -2614 115718 -2378 115954
rect -2934 115398 -2698 115634
rect -2614 115398 -2378 115634
rect -2934 79718 -2698 79954
rect -2614 79718 -2378 79954
rect -2934 79398 -2698 79634
rect -2614 79398 -2378 79634
rect -2934 43718 -2698 43954
rect -2614 43718 -2378 43954
rect -2934 43398 -2698 43634
rect -2614 43398 -2378 43634
rect -2934 7718 -2698 7954
rect -2614 7718 -2378 7954
rect -2934 7398 -2698 7634
rect -2614 7398 -2378 7634
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 6326 705562 6562 705798
rect 6646 705562 6882 705798
rect 6326 705242 6562 705478
rect 6646 705242 6882 705478
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1542 6562 -1306
rect 6646 -1542 6882 -1306
rect 6326 -1862 6562 -1626
rect 6646 -1862 6882 -1626
rect 10826 706522 11062 706758
rect 11146 706522 11382 706758
rect 10826 706202 11062 706438
rect 11146 706202 11382 706438
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2502 11062 -2266
rect 11146 -2502 11382 -2266
rect 10826 -2822 11062 -2586
rect 11146 -2822 11382 -2586
rect 15326 707482 15562 707718
rect 15646 707482 15882 707718
rect 15326 707162 15562 707398
rect 15646 707162 15882 707398
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3462 15562 -3226
rect 15646 -3462 15882 -3226
rect 15326 -3782 15562 -3546
rect 15646 -3782 15882 -3546
rect 19826 708442 20062 708678
rect 20146 708442 20382 708678
rect 19826 708122 20062 708358
rect 20146 708122 20382 708358
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4422 20062 -4186
rect 20146 -4422 20382 -4186
rect 19826 -4742 20062 -4506
rect 20146 -4742 20382 -4506
rect 24326 709402 24562 709638
rect 24646 709402 24882 709638
rect 24326 709082 24562 709318
rect 24646 709082 24882 709318
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 24326 133718 24562 133954
rect 24646 133718 24882 133954
rect 24326 133398 24562 133634
rect 24646 133398 24882 133634
rect 24326 97718 24562 97954
rect 24646 97718 24882 97954
rect 24326 97398 24562 97634
rect 24646 97398 24882 97634
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5382 24562 -5146
rect 24646 -5382 24882 -5146
rect 24326 -5702 24562 -5466
rect 24646 -5702 24882 -5466
rect 28826 710362 29062 710598
rect 29146 710362 29382 710598
rect 28826 710042 29062 710278
rect 29146 710042 29382 710278
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 28826 138218 29062 138454
rect 29146 138218 29382 138454
rect 28826 137898 29062 138134
rect 29146 137898 29382 138134
rect 28826 102218 29062 102454
rect 29146 102218 29382 102454
rect 28826 101898 29062 102134
rect 29146 101898 29382 102134
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6342 29062 -6106
rect 29146 -6342 29382 -6106
rect 28826 -6662 29062 -6426
rect 29146 -6662 29382 -6426
rect 33326 711322 33562 711558
rect 33646 711322 33882 711558
rect 33326 711002 33562 711238
rect 33646 711002 33882 711238
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 33326 646718 33562 646954
rect 33646 646718 33882 646954
rect 33326 646398 33562 646634
rect 33646 646398 33882 646634
rect 33326 610718 33562 610954
rect 33646 610718 33882 610954
rect 33326 610398 33562 610634
rect 33646 610398 33882 610634
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 33326 142718 33562 142954
rect 33646 142718 33882 142954
rect 33326 142398 33562 142634
rect 33646 142398 33882 142634
rect 33326 106718 33562 106954
rect 33646 106718 33882 106954
rect 33326 106398 33562 106634
rect 33646 106398 33882 106634
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7302 33562 -7066
rect 33646 -7302 33882 -7066
rect 33326 -7622 33562 -7386
rect 33646 -7622 33882 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 42326 705562 42562 705798
rect 42646 705562 42882 705798
rect 42326 705242 42562 705478
rect 42646 705242 42882 705478
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 42326 655718 42562 655954
rect 42646 655718 42882 655954
rect 42326 655398 42562 655634
rect 42646 655398 42882 655634
rect 42326 619718 42562 619954
rect 42646 619718 42882 619954
rect 42326 619398 42562 619634
rect 42646 619398 42882 619634
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 42326 151718 42562 151954
rect 42646 151718 42882 151954
rect 42326 151398 42562 151634
rect 42646 151398 42882 151634
rect 42326 115718 42562 115954
rect 42646 115718 42882 115954
rect 42326 115398 42562 115634
rect 42646 115398 42882 115634
rect 42326 79718 42562 79954
rect 42646 79718 42882 79954
rect 42326 79398 42562 79634
rect 42646 79398 42882 79634
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1542 42562 -1306
rect 42646 -1542 42882 -1306
rect 42326 -1862 42562 -1626
rect 42646 -1862 42882 -1626
rect 46826 706522 47062 706758
rect 47146 706522 47382 706758
rect 46826 706202 47062 706438
rect 47146 706202 47382 706438
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 46826 660218 47062 660454
rect 47146 660218 47382 660454
rect 46826 659898 47062 660134
rect 47146 659898 47382 660134
rect 46826 624218 47062 624454
rect 47146 624218 47382 624454
rect 46826 623898 47062 624134
rect 47146 623898 47382 624134
rect 46826 588218 47062 588454
rect 47146 588218 47382 588454
rect 46826 587898 47062 588134
rect 47146 587898 47382 588134
rect 46826 552218 47062 552454
rect 47146 552218 47382 552454
rect 46826 551898 47062 552134
rect 47146 551898 47382 552134
rect 46826 516218 47062 516454
rect 47146 516218 47382 516454
rect 46826 515898 47062 516134
rect 47146 515898 47382 516134
rect 46826 480218 47062 480454
rect 47146 480218 47382 480454
rect 46826 479898 47062 480134
rect 47146 479898 47382 480134
rect 46826 444218 47062 444454
rect 47146 444218 47382 444454
rect 46826 443898 47062 444134
rect 47146 443898 47382 444134
rect 46826 408218 47062 408454
rect 47146 408218 47382 408454
rect 46826 407898 47062 408134
rect 47146 407898 47382 408134
rect 46826 372218 47062 372454
rect 47146 372218 47382 372454
rect 46826 371898 47062 372134
rect 47146 371898 47382 372134
rect 46826 336218 47062 336454
rect 47146 336218 47382 336454
rect 46826 335898 47062 336134
rect 47146 335898 47382 336134
rect 46826 300218 47062 300454
rect 47146 300218 47382 300454
rect 46826 299898 47062 300134
rect 47146 299898 47382 300134
rect 46826 264218 47062 264454
rect 47146 264218 47382 264454
rect 46826 263898 47062 264134
rect 47146 263898 47382 264134
rect 46826 228218 47062 228454
rect 47146 228218 47382 228454
rect 46826 227898 47062 228134
rect 47146 227898 47382 228134
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 46826 84218 47062 84454
rect 47146 84218 47382 84454
rect 46826 83898 47062 84134
rect 47146 83898 47382 84134
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2502 47062 -2266
rect 47146 -2502 47382 -2266
rect 46826 -2822 47062 -2586
rect 47146 -2822 47382 -2586
rect 51326 707482 51562 707718
rect 51646 707482 51882 707718
rect 51326 707162 51562 707398
rect 51646 707162 51882 707398
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 51326 664718 51562 664954
rect 51646 664718 51882 664954
rect 51326 664398 51562 664634
rect 51646 664398 51882 664634
rect 51326 628718 51562 628954
rect 51646 628718 51882 628954
rect 51326 628398 51562 628634
rect 51646 628398 51882 628634
rect 51326 592718 51562 592954
rect 51646 592718 51882 592954
rect 51326 592398 51562 592634
rect 51646 592398 51882 592634
rect 51326 556718 51562 556954
rect 51646 556718 51882 556954
rect 51326 556398 51562 556634
rect 51646 556398 51882 556634
rect 51326 520718 51562 520954
rect 51646 520718 51882 520954
rect 51326 520398 51562 520634
rect 51646 520398 51882 520634
rect 51326 484718 51562 484954
rect 51646 484718 51882 484954
rect 51326 484398 51562 484634
rect 51646 484398 51882 484634
rect 51326 448718 51562 448954
rect 51646 448718 51882 448954
rect 51326 448398 51562 448634
rect 51646 448398 51882 448634
rect 51326 412718 51562 412954
rect 51646 412718 51882 412954
rect 51326 412398 51562 412634
rect 51646 412398 51882 412634
rect 51326 376718 51562 376954
rect 51646 376718 51882 376954
rect 51326 376398 51562 376634
rect 51646 376398 51882 376634
rect 51326 340718 51562 340954
rect 51646 340718 51882 340954
rect 51326 340398 51562 340634
rect 51646 340398 51882 340634
rect 51326 304718 51562 304954
rect 51646 304718 51882 304954
rect 51326 304398 51562 304634
rect 51646 304398 51882 304634
rect 51326 268718 51562 268954
rect 51646 268718 51882 268954
rect 51326 268398 51562 268634
rect 51646 268398 51882 268634
rect 51326 232718 51562 232954
rect 51646 232718 51882 232954
rect 51326 232398 51562 232634
rect 51646 232398 51882 232634
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 51326 124718 51562 124954
rect 51646 124718 51882 124954
rect 51326 124398 51562 124634
rect 51646 124398 51882 124634
rect 51326 88718 51562 88954
rect 51646 88718 51882 88954
rect 51326 88398 51562 88634
rect 51646 88398 51882 88634
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3462 51562 -3226
rect 51646 -3462 51882 -3226
rect 51326 -3782 51562 -3546
rect 51646 -3782 51882 -3546
rect 55826 708442 56062 708678
rect 56146 708442 56382 708678
rect 55826 708122 56062 708358
rect 56146 708122 56382 708358
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4422 56062 -4186
rect 56146 -4422 56382 -4186
rect 55826 -4742 56062 -4506
rect 56146 -4742 56382 -4506
rect 60326 709402 60562 709638
rect 60646 709402 60882 709638
rect 60326 709082 60562 709318
rect 60646 709082 60882 709318
rect 60326 673718 60562 673954
rect 60646 673718 60882 673954
rect 60326 673398 60562 673634
rect 60646 673398 60882 673634
rect 60326 637718 60562 637954
rect 60646 637718 60882 637954
rect 60326 637398 60562 637634
rect 60646 637398 60882 637634
rect 60326 601718 60562 601954
rect 60646 601718 60882 601954
rect 60326 601398 60562 601634
rect 60646 601398 60882 601634
rect 60326 565718 60562 565954
rect 60646 565718 60882 565954
rect 60326 565398 60562 565634
rect 60646 565398 60882 565634
rect 60326 529718 60562 529954
rect 60646 529718 60882 529954
rect 60326 529398 60562 529634
rect 60646 529398 60882 529634
rect 60326 493718 60562 493954
rect 60646 493718 60882 493954
rect 60326 493398 60562 493634
rect 60646 493398 60882 493634
rect 60326 457718 60562 457954
rect 60646 457718 60882 457954
rect 60326 457398 60562 457634
rect 60646 457398 60882 457634
rect 60326 421718 60562 421954
rect 60646 421718 60882 421954
rect 60326 421398 60562 421634
rect 60646 421398 60882 421634
rect 60326 385718 60562 385954
rect 60646 385718 60882 385954
rect 60326 385398 60562 385634
rect 60646 385398 60882 385634
rect 60326 349718 60562 349954
rect 60646 349718 60882 349954
rect 60326 349398 60562 349634
rect 60646 349398 60882 349634
rect 60326 313718 60562 313954
rect 60646 313718 60882 313954
rect 60326 313398 60562 313634
rect 60646 313398 60882 313634
rect 60326 277718 60562 277954
rect 60646 277718 60882 277954
rect 60326 277398 60562 277634
rect 60646 277398 60882 277634
rect 60326 241718 60562 241954
rect 60646 241718 60882 241954
rect 60326 241398 60562 241634
rect 60646 241398 60882 241634
rect 60326 205718 60562 205954
rect 60646 205718 60882 205954
rect 60326 205398 60562 205634
rect 60646 205398 60882 205634
rect 60326 169718 60562 169954
rect 60646 169718 60882 169954
rect 60326 169398 60562 169634
rect 60646 169398 60882 169634
rect 60326 133718 60562 133954
rect 60646 133718 60882 133954
rect 60326 133398 60562 133634
rect 60646 133398 60882 133634
rect 60326 97718 60562 97954
rect 60646 97718 60882 97954
rect 60326 97398 60562 97634
rect 60646 97398 60882 97634
rect 60326 61718 60562 61954
rect 60646 61718 60882 61954
rect 60326 61398 60562 61634
rect 60646 61398 60882 61634
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 60326 -5382 60562 -5146
rect 60646 -5382 60882 -5146
rect 60326 -5702 60562 -5466
rect 60646 -5702 60882 -5466
rect 64826 710362 65062 710598
rect 65146 710362 65382 710598
rect 64826 710042 65062 710278
rect 65146 710042 65382 710278
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 64826 642218 65062 642454
rect 65146 642218 65382 642454
rect 64826 641898 65062 642134
rect 65146 641898 65382 642134
rect 64826 606218 65062 606454
rect 65146 606218 65382 606454
rect 64826 605898 65062 606134
rect 65146 605898 65382 606134
rect 64826 570218 65062 570454
rect 65146 570218 65382 570454
rect 64826 569898 65062 570134
rect 65146 569898 65382 570134
rect 64826 534218 65062 534454
rect 65146 534218 65382 534454
rect 64826 533898 65062 534134
rect 65146 533898 65382 534134
rect 64826 498218 65062 498454
rect 65146 498218 65382 498454
rect 64826 497898 65062 498134
rect 65146 497898 65382 498134
rect 64826 462218 65062 462454
rect 65146 462218 65382 462454
rect 64826 461898 65062 462134
rect 65146 461898 65382 462134
rect 64826 426218 65062 426454
rect 65146 426218 65382 426454
rect 64826 425898 65062 426134
rect 65146 425898 65382 426134
rect 64826 390218 65062 390454
rect 65146 390218 65382 390454
rect 64826 389898 65062 390134
rect 65146 389898 65382 390134
rect 64826 354218 65062 354454
rect 65146 354218 65382 354454
rect 64826 353898 65062 354134
rect 65146 353898 65382 354134
rect 64826 318218 65062 318454
rect 65146 318218 65382 318454
rect 64826 317898 65062 318134
rect 65146 317898 65382 318134
rect 64826 282218 65062 282454
rect 65146 282218 65382 282454
rect 64826 281898 65062 282134
rect 65146 281898 65382 282134
rect 64826 246218 65062 246454
rect 65146 246218 65382 246454
rect 64826 245898 65062 246134
rect 65146 245898 65382 246134
rect 64826 210218 65062 210454
rect 65146 210218 65382 210454
rect 64826 209898 65062 210134
rect 65146 209898 65382 210134
rect 64826 174218 65062 174454
rect 65146 174218 65382 174454
rect 64826 173898 65062 174134
rect 65146 173898 65382 174134
rect 64826 138218 65062 138454
rect 65146 138218 65382 138454
rect 64826 137898 65062 138134
rect 65146 137898 65382 138134
rect 64826 102218 65062 102454
rect 65146 102218 65382 102454
rect 64826 101898 65062 102134
rect 65146 101898 65382 102134
rect 64826 66218 65062 66454
rect 65146 66218 65382 66454
rect 64826 65898 65062 66134
rect 65146 65898 65382 66134
rect 64826 30218 65062 30454
rect 65146 30218 65382 30454
rect 64826 29898 65062 30134
rect 65146 29898 65382 30134
rect 64826 -6342 65062 -6106
rect 65146 -6342 65382 -6106
rect 64826 -6662 65062 -6426
rect 65146 -6662 65382 -6426
rect 69326 711322 69562 711558
rect 69646 711322 69882 711558
rect 69326 711002 69562 711238
rect 69646 711002 69882 711238
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 69326 646718 69562 646954
rect 69646 646718 69882 646954
rect 69326 646398 69562 646634
rect 69646 646398 69882 646634
rect 69326 610718 69562 610954
rect 69646 610718 69882 610954
rect 69326 610398 69562 610634
rect 69646 610398 69882 610634
rect 69326 574718 69562 574954
rect 69646 574718 69882 574954
rect 69326 574398 69562 574634
rect 69646 574398 69882 574634
rect 69326 538718 69562 538954
rect 69646 538718 69882 538954
rect 69326 538398 69562 538634
rect 69646 538398 69882 538634
rect 69326 502718 69562 502954
rect 69646 502718 69882 502954
rect 69326 502398 69562 502634
rect 69646 502398 69882 502634
rect 69326 466718 69562 466954
rect 69646 466718 69882 466954
rect 69326 466398 69562 466634
rect 69646 466398 69882 466634
rect 69326 430718 69562 430954
rect 69646 430718 69882 430954
rect 69326 430398 69562 430634
rect 69646 430398 69882 430634
rect 69326 394718 69562 394954
rect 69646 394718 69882 394954
rect 69326 394398 69562 394634
rect 69646 394398 69882 394634
rect 69326 358718 69562 358954
rect 69646 358718 69882 358954
rect 69326 358398 69562 358634
rect 69646 358398 69882 358634
rect 69326 322718 69562 322954
rect 69646 322718 69882 322954
rect 69326 322398 69562 322634
rect 69646 322398 69882 322634
rect 69326 286718 69562 286954
rect 69646 286718 69882 286954
rect 69326 286398 69562 286634
rect 69646 286398 69882 286634
rect 69326 250718 69562 250954
rect 69646 250718 69882 250954
rect 69326 250398 69562 250634
rect 69646 250398 69882 250634
rect 69326 214718 69562 214954
rect 69646 214718 69882 214954
rect 69326 214398 69562 214634
rect 69646 214398 69882 214634
rect 69326 178718 69562 178954
rect 69646 178718 69882 178954
rect 69326 178398 69562 178634
rect 69646 178398 69882 178634
rect 69326 142718 69562 142954
rect 69646 142718 69882 142954
rect 69326 142398 69562 142634
rect 69646 142398 69882 142634
rect 69326 106718 69562 106954
rect 69646 106718 69882 106954
rect 69326 106398 69562 106634
rect 69646 106398 69882 106634
rect 69326 70718 69562 70954
rect 69646 70718 69882 70954
rect 69326 70398 69562 70634
rect 69646 70398 69882 70634
rect 69326 34718 69562 34954
rect 69646 34718 69882 34954
rect 69326 34398 69562 34634
rect 69646 34398 69882 34634
rect 69326 -7302 69562 -7066
rect 69646 -7302 69882 -7066
rect 69326 -7622 69562 -7386
rect 69646 -7622 69882 -7386
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 78326 705562 78562 705798
rect 78646 705562 78882 705798
rect 78326 705242 78562 705478
rect 78646 705242 78882 705478
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 78326 655718 78562 655954
rect 78646 655718 78882 655954
rect 78326 655398 78562 655634
rect 78646 655398 78882 655634
rect 78326 619718 78562 619954
rect 78646 619718 78882 619954
rect 78326 619398 78562 619634
rect 78646 619398 78882 619634
rect 78326 583718 78562 583954
rect 78646 583718 78882 583954
rect 78326 583398 78562 583634
rect 78646 583398 78882 583634
rect 78326 547718 78562 547954
rect 78646 547718 78882 547954
rect 78326 547398 78562 547634
rect 78646 547398 78882 547634
rect 78326 511718 78562 511954
rect 78646 511718 78882 511954
rect 78326 511398 78562 511634
rect 78646 511398 78882 511634
rect 78326 475718 78562 475954
rect 78646 475718 78882 475954
rect 78326 475398 78562 475634
rect 78646 475398 78882 475634
rect 78326 439718 78562 439954
rect 78646 439718 78882 439954
rect 78326 439398 78562 439634
rect 78646 439398 78882 439634
rect 78326 403718 78562 403954
rect 78646 403718 78882 403954
rect 78326 403398 78562 403634
rect 78646 403398 78882 403634
rect 78326 367718 78562 367954
rect 78646 367718 78882 367954
rect 78326 367398 78562 367634
rect 78646 367398 78882 367634
rect 78326 331718 78562 331954
rect 78646 331718 78882 331954
rect 78326 331398 78562 331634
rect 78646 331398 78882 331634
rect 78326 295718 78562 295954
rect 78646 295718 78882 295954
rect 78326 295398 78562 295634
rect 78646 295398 78882 295634
rect 78326 259718 78562 259954
rect 78646 259718 78882 259954
rect 78326 259398 78562 259634
rect 78646 259398 78882 259634
rect 78326 223718 78562 223954
rect 78646 223718 78882 223954
rect 78326 223398 78562 223634
rect 78646 223398 78882 223634
rect 78326 187718 78562 187954
rect 78646 187718 78882 187954
rect 78326 187398 78562 187634
rect 78646 187398 78882 187634
rect 78326 151718 78562 151954
rect 78646 151718 78882 151954
rect 78326 151398 78562 151634
rect 78646 151398 78882 151634
rect 78326 115718 78562 115954
rect 78646 115718 78882 115954
rect 78326 115398 78562 115634
rect 78646 115398 78882 115634
rect 78326 79718 78562 79954
rect 78646 79718 78882 79954
rect 78326 79398 78562 79634
rect 78646 79398 78882 79634
rect 78326 43718 78562 43954
rect 78646 43718 78882 43954
rect 78326 43398 78562 43634
rect 78646 43398 78882 43634
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1542 78562 -1306
rect 78646 -1542 78882 -1306
rect 78326 -1862 78562 -1626
rect 78646 -1862 78882 -1626
rect 82826 706522 83062 706758
rect 83146 706522 83382 706758
rect 82826 706202 83062 706438
rect 83146 706202 83382 706438
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 82826 660218 83062 660454
rect 83146 660218 83382 660454
rect 82826 659898 83062 660134
rect 83146 659898 83382 660134
rect 82826 624218 83062 624454
rect 83146 624218 83382 624454
rect 82826 623898 83062 624134
rect 83146 623898 83382 624134
rect 82826 588218 83062 588454
rect 83146 588218 83382 588454
rect 82826 587898 83062 588134
rect 83146 587898 83382 588134
rect 82826 552218 83062 552454
rect 83146 552218 83382 552454
rect 82826 551898 83062 552134
rect 83146 551898 83382 552134
rect 82826 516218 83062 516454
rect 83146 516218 83382 516454
rect 82826 515898 83062 516134
rect 83146 515898 83382 516134
rect 82826 480218 83062 480454
rect 83146 480218 83382 480454
rect 82826 479898 83062 480134
rect 83146 479898 83382 480134
rect 82826 444218 83062 444454
rect 83146 444218 83382 444454
rect 82826 443898 83062 444134
rect 83146 443898 83382 444134
rect 82826 408218 83062 408454
rect 83146 408218 83382 408454
rect 82826 407898 83062 408134
rect 83146 407898 83382 408134
rect 82826 372218 83062 372454
rect 83146 372218 83382 372454
rect 82826 371898 83062 372134
rect 83146 371898 83382 372134
rect 82826 336218 83062 336454
rect 83146 336218 83382 336454
rect 82826 335898 83062 336134
rect 83146 335898 83382 336134
rect 82826 300218 83062 300454
rect 83146 300218 83382 300454
rect 82826 299898 83062 300134
rect 83146 299898 83382 300134
rect 82826 264218 83062 264454
rect 83146 264218 83382 264454
rect 82826 263898 83062 264134
rect 83146 263898 83382 264134
rect 82826 228218 83062 228454
rect 83146 228218 83382 228454
rect 82826 227898 83062 228134
rect 83146 227898 83382 228134
rect 82826 192218 83062 192454
rect 83146 192218 83382 192454
rect 82826 191898 83062 192134
rect 83146 191898 83382 192134
rect 82826 156218 83062 156454
rect 83146 156218 83382 156454
rect 82826 155898 83062 156134
rect 83146 155898 83382 156134
rect 82826 120218 83062 120454
rect 83146 120218 83382 120454
rect 82826 119898 83062 120134
rect 83146 119898 83382 120134
rect 82826 84218 83062 84454
rect 83146 84218 83382 84454
rect 82826 83898 83062 84134
rect 83146 83898 83382 84134
rect 82826 48218 83062 48454
rect 83146 48218 83382 48454
rect 82826 47898 83062 48134
rect 83146 47898 83382 48134
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2502 83062 -2266
rect 83146 -2502 83382 -2266
rect 82826 -2822 83062 -2586
rect 83146 -2822 83382 -2586
rect 87326 707482 87562 707718
rect 87646 707482 87882 707718
rect 87326 707162 87562 707398
rect 87646 707162 87882 707398
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 87326 664718 87562 664954
rect 87646 664718 87882 664954
rect 87326 664398 87562 664634
rect 87646 664398 87882 664634
rect 87326 628718 87562 628954
rect 87646 628718 87882 628954
rect 87326 628398 87562 628634
rect 87646 628398 87882 628634
rect 87326 592718 87562 592954
rect 87646 592718 87882 592954
rect 87326 592398 87562 592634
rect 87646 592398 87882 592634
rect 87326 556718 87562 556954
rect 87646 556718 87882 556954
rect 87326 556398 87562 556634
rect 87646 556398 87882 556634
rect 87326 520718 87562 520954
rect 87646 520718 87882 520954
rect 87326 520398 87562 520634
rect 87646 520398 87882 520634
rect 87326 484718 87562 484954
rect 87646 484718 87882 484954
rect 87326 484398 87562 484634
rect 87646 484398 87882 484634
rect 87326 448718 87562 448954
rect 87646 448718 87882 448954
rect 87326 448398 87562 448634
rect 87646 448398 87882 448634
rect 87326 412718 87562 412954
rect 87646 412718 87882 412954
rect 87326 412398 87562 412634
rect 87646 412398 87882 412634
rect 87326 376718 87562 376954
rect 87646 376718 87882 376954
rect 87326 376398 87562 376634
rect 87646 376398 87882 376634
rect 87326 340718 87562 340954
rect 87646 340718 87882 340954
rect 87326 340398 87562 340634
rect 87646 340398 87882 340634
rect 87326 304718 87562 304954
rect 87646 304718 87882 304954
rect 87326 304398 87562 304634
rect 87646 304398 87882 304634
rect 87326 268718 87562 268954
rect 87646 268718 87882 268954
rect 87326 268398 87562 268634
rect 87646 268398 87882 268634
rect 87326 232718 87562 232954
rect 87646 232718 87882 232954
rect 87326 232398 87562 232634
rect 87646 232398 87882 232634
rect 87326 196718 87562 196954
rect 87646 196718 87882 196954
rect 87326 196398 87562 196634
rect 87646 196398 87882 196634
rect 87326 160718 87562 160954
rect 87646 160718 87882 160954
rect 87326 160398 87562 160634
rect 87646 160398 87882 160634
rect 87326 124718 87562 124954
rect 87646 124718 87882 124954
rect 87326 124398 87562 124634
rect 87646 124398 87882 124634
rect 87326 88718 87562 88954
rect 87646 88718 87882 88954
rect 87326 88398 87562 88634
rect 87646 88398 87882 88634
rect 87326 52718 87562 52954
rect 87646 52718 87882 52954
rect 87326 52398 87562 52634
rect 87646 52398 87882 52634
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3462 87562 -3226
rect 87646 -3462 87882 -3226
rect 87326 -3782 87562 -3546
rect 87646 -3782 87882 -3546
rect 91826 708442 92062 708678
rect 92146 708442 92382 708678
rect 91826 708122 92062 708358
rect 92146 708122 92382 708358
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4422 92062 -4186
rect 92146 -4422 92382 -4186
rect 91826 -4742 92062 -4506
rect 92146 -4742 92382 -4506
rect 96326 709402 96562 709638
rect 96646 709402 96882 709638
rect 96326 709082 96562 709318
rect 96646 709082 96882 709318
rect 96326 673718 96562 673954
rect 96646 673718 96882 673954
rect 96326 673398 96562 673634
rect 96646 673398 96882 673634
rect 96326 637718 96562 637954
rect 96646 637718 96882 637954
rect 96326 637398 96562 637634
rect 96646 637398 96882 637634
rect 96326 601718 96562 601954
rect 96646 601718 96882 601954
rect 96326 601398 96562 601634
rect 96646 601398 96882 601634
rect 96326 565718 96562 565954
rect 96646 565718 96882 565954
rect 96326 565398 96562 565634
rect 96646 565398 96882 565634
rect 96326 529718 96562 529954
rect 96646 529718 96882 529954
rect 96326 529398 96562 529634
rect 96646 529398 96882 529634
rect 96326 493718 96562 493954
rect 96646 493718 96882 493954
rect 96326 493398 96562 493634
rect 96646 493398 96882 493634
rect 96326 457718 96562 457954
rect 96646 457718 96882 457954
rect 96326 457398 96562 457634
rect 96646 457398 96882 457634
rect 96326 421718 96562 421954
rect 96646 421718 96882 421954
rect 96326 421398 96562 421634
rect 96646 421398 96882 421634
rect 96326 385718 96562 385954
rect 96646 385718 96882 385954
rect 96326 385398 96562 385634
rect 96646 385398 96882 385634
rect 96326 349718 96562 349954
rect 96646 349718 96882 349954
rect 96326 349398 96562 349634
rect 96646 349398 96882 349634
rect 96326 313718 96562 313954
rect 96646 313718 96882 313954
rect 96326 313398 96562 313634
rect 96646 313398 96882 313634
rect 96326 277718 96562 277954
rect 96646 277718 96882 277954
rect 96326 277398 96562 277634
rect 96646 277398 96882 277634
rect 96326 241718 96562 241954
rect 96646 241718 96882 241954
rect 96326 241398 96562 241634
rect 96646 241398 96882 241634
rect 96326 205718 96562 205954
rect 96646 205718 96882 205954
rect 96326 205398 96562 205634
rect 96646 205398 96882 205634
rect 100826 710362 101062 710598
rect 101146 710362 101382 710598
rect 100826 710042 101062 710278
rect 101146 710042 101382 710278
rect 100826 678218 101062 678454
rect 101146 678218 101382 678454
rect 100826 677898 101062 678134
rect 101146 677898 101382 678134
rect 100826 642218 101062 642454
rect 101146 642218 101382 642454
rect 100826 641898 101062 642134
rect 101146 641898 101382 642134
rect 100826 606218 101062 606454
rect 101146 606218 101382 606454
rect 100826 605898 101062 606134
rect 101146 605898 101382 606134
rect 100826 570218 101062 570454
rect 101146 570218 101382 570454
rect 100826 569898 101062 570134
rect 101146 569898 101382 570134
rect 100826 534218 101062 534454
rect 101146 534218 101382 534454
rect 100826 533898 101062 534134
rect 101146 533898 101382 534134
rect 100826 498218 101062 498454
rect 101146 498218 101382 498454
rect 100826 497898 101062 498134
rect 101146 497898 101382 498134
rect 100826 462218 101062 462454
rect 101146 462218 101382 462454
rect 100826 461898 101062 462134
rect 101146 461898 101382 462134
rect 100826 426218 101062 426454
rect 101146 426218 101382 426454
rect 100826 425898 101062 426134
rect 101146 425898 101382 426134
rect 100826 390218 101062 390454
rect 101146 390218 101382 390454
rect 100826 389898 101062 390134
rect 101146 389898 101382 390134
rect 100826 354218 101062 354454
rect 101146 354218 101382 354454
rect 100826 353898 101062 354134
rect 101146 353898 101382 354134
rect 100826 318218 101062 318454
rect 101146 318218 101382 318454
rect 100826 317898 101062 318134
rect 101146 317898 101382 318134
rect 100826 282218 101062 282454
rect 101146 282218 101382 282454
rect 100826 281898 101062 282134
rect 101146 281898 101382 282134
rect 100826 246218 101062 246454
rect 101146 246218 101382 246454
rect 100826 245898 101062 246134
rect 101146 245898 101382 246134
rect 100826 210218 101062 210454
rect 101146 210218 101382 210454
rect 100826 209898 101062 210134
rect 101146 209898 101382 210134
rect 96326 169718 96562 169954
rect 96646 169718 96882 169954
rect 96326 169398 96562 169634
rect 96646 169398 96882 169634
rect 96326 133718 96562 133954
rect 96646 133718 96882 133954
rect 96326 133398 96562 133634
rect 96646 133398 96882 133634
rect 96326 97718 96562 97954
rect 96646 97718 96882 97954
rect 96326 97398 96562 97634
rect 96646 97398 96882 97634
rect 96326 61718 96562 61954
rect 96646 61718 96882 61954
rect 96326 61398 96562 61634
rect 96646 61398 96882 61634
rect 105326 711322 105562 711558
rect 105646 711322 105882 711558
rect 105326 711002 105562 711238
rect 105646 711002 105882 711238
rect 105326 682718 105562 682954
rect 105646 682718 105882 682954
rect 105326 682398 105562 682634
rect 105646 682398 105882 682634
rect 105326 646718 105562 646954
rect 105646 646718 105882 646954
rect 105326 646398 105562 646634
rect 105646 646398 105882 646634
rect 105326 610718 105562 610954
rect 105646 610718 105882 610954
rect 105326 610398 105562 610634
rect 105646 610398 105882 610634
rect 105326 574718 105562 574954
rect 105646 574718 105882 574954
rect 105326 574398 105562 574634
rect 105646 574398 105882 574634
rect 105326 538718 105562 538954
rect 105646 538718 105882 538954
rect 105326 538398 105562 538634
rect 105646 538398 105882 538634
rect 105326 502718 105562 502954
rect 105646 502718 105882 502954
rect 105326 502398 105562 502634
rect 105646 502398 105882 502634
rect 105326 466718 105562 466954
rect 105646 466718 105882 466954
rect 105326 466398 105562 466634
rect 105646 466398 105882 466634
rect 105326 430718 105562 430954
rect 105646 430718 105882 430954
rect 105326 430398 105562 430634
rect 105646 430398 105882 430634
rect 105326 394718 105562 394954
rect 105646 394718 105882 394954
rect 105326 394398 105562 394634
rect 105646 394398 105882 394634
rect 105326 358718 105562 358954
rect 105646 358718 105882 358954
rect 105326 358398 105562 358634
rect 105646 358398 105882 358634
rect 105326 322718 105562 322954
rect 105646 322718 105882 322954
rect 105326 322398 105562 322634
rect 105646 322398 105882 322634
rect 105326 286718 105562 286954
rect 105646 286718 105882 286954
rect 105326 286398 105562 286634
rect 105646 286398 105882 286634
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 105326 250718 105562 250954
rect 105646 250718 105882 250954
rect 105326 250398 105562 250634
rect 105646 250398 105882 250634
rect 105326 214718 105562 214954
rect 105646 214718 105882 214954
rect 105326 214398 105562 214634
rect 105646 214398 105882 214634
rect 100826 174218 101062 174454
rect 101146 174218 101382 174454
rect 100826 173898 101062 174134
rect 101146 173898 101382 174134
rect 100826 138218 101062 138454
rect 101146 138218 101382 138454
rect 100826 137898 101062 138134
rect 101146 137898 101382 138134
rect 100826 102218 101062 102454
rect 101146 102218 101382 102454
rect 100826 101898 101062 102134
rect 101146 101898 101382 102134
rect 100826 66218 101062 66454
rect 101146 66218 101382 66454
rect 100826 65898 101062 66134
rect 101146 65898 101382 66134
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 96326 -5382 96562 -5146
rect 96646 -5382 96882 -5146
rect 96326 -5702 96562 -5466
rect 96646 -5702 96882 -5466
rect 105326 178718 105562 178954
rect 105646 178718 105882 178954
rect 105326 178398 105562 178634
rect 105646 178398 105882 178634
rect 105326 142718 105562 142954
rect 105646 142718 105882 142954
rect 105326 142398 105562 142634
rect 105646 142398 105882 142634
rect 105326 106718 105562 106954
rect 105646 106718 105882 106954
rect 105326 106398 105562 106634
rect 105646 106398 105882 106634
rect 105326 70718 105562 70954
rect 105646 70718 105882 70954
rect 105326 70398 105562 70634
rect 105646 70398 105882 70634
rect 100826 30218 101062 30454
rect 101146 30218 101382 30454
rect 100826 29898 101062 30134
rect 101146 29898 101382 30134
rect 100826 -6342 101062 -6106
rect 101146 -6342 101382 -6106
rect 100826 -6662 101062 -6426
rect 101146 -6662 101382 -6426
rect 114326 705562 114562 705798
rect 114646 705562 114882 705798
rect 114326 705242 114562 705478
rect 114646 705242 114882 705478
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 114326 655718 114562 655954
rect 114646 655718 114882 655954
rect 114326 655398 114562 655634
rect 114646 655398 114882 655634
rect 114326 619718 114562 619954
rect 114646 619718 114882 619954
rect 114326 619398 114562 619634
rect 114646 619398 114882 619634
rect 114326 583718 114562 583954
rect 114646 583718 114882 583954
rect 114326 583398 114562 583634
rect 114646 583398 114882 583634
rect 114326 547718 114562 547954
rect 114646 547718 114882 547954
rect 114326 547398 114562 547634
rect 114646 547398 114882 547634
rect 114326 511718 114562 511954
rect 114646 511718 114882 511954
rect 114326 511398 114562 511634
rect 114646 511398 114882 511634
rect 114326 475718 114562 475954
rect 114646 475718 114882 475954
rect 114326 475398 114562 475634
rect 114646 475398 114882 475634
rect 114326 439718 114562 439954
rect 114646 439718 114882 439954
rect 114326 439398 114562 439634
rect 114646 439398 114882 439634
rect 114326 403718 114562 403954
rect 114646 403718 114882 403954
rect 114326 403398 114562 403634
rect 114646 403398 114882 403634
rect 114326 367718 114562 367954
rect 114646 367718 114882 367954
rect 114326 367398 114562 367634
rect 114646 367398 114882 367634
rect 114326 331718 114562 331954
rect 114646 331718 114882 331954
rect 114326 331398 114562 331634
rect 114646 331398 114882 331634
rect 114326 295718 114562 295954
rect 114646 295718 114882 295954
rect 114326 295398 114562 295634
rect 114646 295398 114882 295634
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 105326 -7302 105562 -7066
rect 105646 -7302 105882 -7066
rect 105326 -7622 105562 -7386
rect 105646 -7622 105882 -7386
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 118826 706522 119062 706758
rect 119146 706522 119382 706758
rect 118826 706202 119062 706438
rect 119146 706202 119382 706438
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 118826 660218 119062 660454
rect 119146 660218 119382 660454
rect 118826 659898 119062 660134
rect 119146 659898 119382 660134
rect 118826 624218 119062 624454
rect 119146 624218 119382 624454
rect 118826 623898 119062 624134
rect 119146 623898 119382 624134
rect 118826 588218 119062 588454
rect 119146 588218 119382 588454
rect 118826 587898 119062 588134
rect 119146 587898 119382 588134
rect 118826 552218 119062 552454
rect 119146 552218 119382 552454
rect 118826 551898 119062 552134
rect 119146 551898 119382 552134
rect 118826 516218 119062 516454
rect 119146 516218 119382 516454
rect 118826 515898 119062 516134
rect 119146 515898 119382 516134
rect 118826 480218 119062 480454
rect 119146 480218 119382 480454
rect 118826 479898 119062 480134
rect 119146 479898 119382 480134
rect 118826 444218 119062 444454
rect 119146 444218 119382 444454
rect 118826 443898 119062 444134
rect 119146 443898 119382 444134
rect 118826 408218 119062 408454
rect 119146 408218 119382 408454
rect 118826 407898 119062 408134
rect 119146 407898 119382 408134
rect 118826 372218 119062 372454
rect 119146 372218 119382 372454
rect 118826 371898 119062 372134
rect 119146 371898 119382 372134
rect 118826 336218 119062 336454
rect 119146 336218 119382 336454
rect 118826 335898 119062 336134
rect 119146 335898 119382 336134
rect 118826 300218 119062 300454
rect 119146 300218 119382 300454
rect 118826 299898 119062 300134
rect 119146 299898 119382 300134
rect 114326 259718 114562 259954
rect 114646 259718 114882 259954
rect 114326 259398 114562 259634
rect 114646 259398 114882 259634
rect 114326 223718 114562 223954
rect 114646 223718 114882 223954
rect 114326 223398 114562 223634
rect 114646 223398 114882 223634
rect 114326 187718 114562 187954
rect 114646 187718 114882 187954
rect 114326 187398 114562 187634
rect 114646 187398 114882 187634
rect 114326 151718 114562 151954
rect 114646 151718 114882 151954
rect 114326 151398 114562 151634
rect 114646 151398 114882 151634
rect 114326 115718 114562 115954
rect 114646 115718 114882 115954
rect 114326 115398 114562 115634
rect 114646 115398 114882 115634
rect 114326 79718 114562 79954
rect 114646 79718 114882 79954
rect 114326 79398 114562 79634
rect 114646 79398 114882 79634
rect 118826 264218 119062 264454
rect 119146 264218 119382 264454
rect 118826 263898 119062 264134
rect 119146 263898 119382 264134
rect 123326 707482 123562 707718
rect 123646 707482 123882 707718
rect 123326 707162 123562 707398
rect 123646 707162 123882 707398
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 123326 664718 123562 664954
rect 123646 664718 123882 664954
rect 123326 664398 123562 664634
rect 123646 664398 123882 664634
rect 123326 628718 123562 628954
rect 123646 628718 123882 628954
rect 123326 628398 123562 628634
rect 123646 628398 123882 628634
rect 123326 592718 123562 592954
rect 123646 592718 123882 592954
rect 123326 592398 123562 592634
rect 123646 592398 123882 592634
rect 123326 556718 123562 556954
rect 123646 556718 123882 556954
rect 123326 556398 123562 556634
rect 123646 556398 123882 556634
rect 123326 520718 123562 520954
rect 123646 520718 123882 520954
rect 123326 520398 123562 520634
rect 123646 520398 123882 520634
rect 123326 484718 123562 484954
rect 123646 484718 123882 484954
rect 123326 484398 123562 484634
rect 123646 484398 123882 484634
rect 123326 448718 123562 448954
rect 123646 448718 123882 448954
rect 123326 448398 123562 448634
rect 123646 448398 123882 448634
rect 123326 412718 123562 412954
rect 123646 412718 123882 412954
rect 123326 412398 123562 412634
rect 123646 412398 123882 412634
rect 123326 376718 123562 376954
rect 123646 376718 123882 376954
rect 123326 376398 123562 376634
rect 123646 376398 123882 376634
rect 123326 340718 123562 340954
rect 123646 340718 123882 340954
rect 123326 340398 123562 340634
rect 123646 340398 123882 340634
rect 123326 304718 123562 304954
rect 123646 304718 123882 304954
rect 123326 304398 123562 304634
rect 123646 304398 123882 304634
rect 123326 268718 123562 268954
rect 123646 268718 123882 268954
rect 123326 268398 123562 268634
rect 123646 268398 123882 268634
rect 118826 192218 119062 192454
rect 119146 192218 119382 192454
rect 118826 191898 119062 192134
rect 119146 191898 119382 192134
rect 118826 156218 119062 156454
rect 119146 156218 119382 156454
rect 118826 155898 119062 156134
rect 119146 155898 119382 156134
rect 127826 708442 128062 708678
rect 128146 708442 128382 708678
rect 127826 708122 128062 708358
rect 128146 708122 128382 708358
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 132326 709402 132562 709638
rect 132646 709402 132882 709638
rect 132326 709082 132562 709318
rect 132646 709082 132882 709318
rect 132326 673718 132562 673954
rect 132646 673718 132882 673954
rect 132326 673398 132562 673634
rect 132646 673398 132882 673634
rect 132326 637718 132562 637954
rect 132646 637718 132882 637954
rect 132326 637398 132562 637634
rect 132646 637398 132882 637634
rect 132326 601718 132562 601954
rect 132646 601718 132882 601954
rect 132326 601398 132562 601634
rect 132646 601398 132882 601634
rect 132326 565718 132562 565954
rect 132646 565718 132882 565954
rect 132326 565398 132562 565634
rect 132646 565398 132882 565634
rect 132326 529718 132562 529954
rect 132646 529718 132882 529954
rect 132326 529398 132562 529634
rect 132646 529398 132882 529634
rect 132326 493718 132562 493954
rect 132646 493718 132882 493954
rect 132326 493398 132562 493634
rect 132646 493398 132882 493634
rect 132326 457718 132562 457954
rect 132646 457718 132882 457954
rect 132326 457398 132562 457634
rect 132646 457398 132882 457634
rect 132326 421718 132562 421954
rect 132646 421718 132882 421954
rect 132326 421398 132562 421634
rect 132646 421398 132882 421634
rect 132326 385718 132562 385954
rect 132646 385718 132882 385954
rect 132326 385398 132562 385634
rect 132646 385398 132882 385634
rect 132326 349718 132562 349954
rect 132646 349718 132882 349954
rect 132326 349398 132562 349634
rect 132646 349398 132882 349634
rect 132326 313718 132562 313954
rect 132646 313718 132882 313954
rect 132326 313398 132562 313634
rect 132646 313398 132882 313634
rect 132326 277718 132562 277954
rect 132646 277718 132882 277954
rect 132326 277398 132562 277634
rect 132646 277398 132882 277634
rect 136826 710362 137062 710598
rect 137146 710362 137382 710598
rect 136826 710042 137062 710278
rect 137146 710042 137382 710278
rect 136826 678218 137062 678454
rect 137146 678218 137382 678454
rect 136826 677898 137062 678134
rect 137146 677898 137382 678134
rect 136826 642218 137062 642454
rect 137146 642218 137382 642454
rect 136826 641898 137062 642134
rect 137146 641898 137382 642134
rect 136826 606218 137062 606454
rect 137146 606218 137382 606454
rect 136826 605898 137062 606134
rect 137146 605898 137382 606134
rect 136826 570218 137062 570454
rect 137146 570218 137382 570454
rect 136826 569898 137062 570134
rect 137146 569898 137382 570134
rect 136826 534218 137062 534454
rect 137146 534218 137382 534454
rect 136826 533898 137062 534134
rect 137146 533898 137382 534134
rect 136826 498218 137062 498454
rect 137146 498218 137382 498454
rect 136826 497898 137062 498134
rect 137146 497898 137382 498134
rect 136826 462218 137062 462454
rect 137146 462218 137382 462454
rect 136826 461898 137062 462134
rect 137146 461898 137382 462134
rect 136826 426218 137062 426454
rect 137146 426218 137382 426454
rect 136826 425898 137062 426134
rect 137146 425898 137382 426134
rect 136826 390218 137062 390454
rect 137146 390218 137382 390454
rect 136826 389898 137062 390134
rect 137146 389898 137382 390134
rect 136826 354218 137062 354454
rect 137146 354218 137382 354454
rect 136826 353898 137062 354134
rect 137146 353898 137382 354134
rect 136826 318218 137062 318454
rect 137146 318218 137382 318454
rect 136826 317898 137062 318134
rect 137146 317898 137382 318134
rect 136826 282218 137062 282454
rect 137146 282218 137382 282454
rect 136826 281898 137062 282134
rect 137146 281898 137382 282134
rect 141326 711322 141562 711558
rect 141646 711322 141882 711558
rect 141326 711002 141562 711238
rect 141646 711002 141882 711238
rect 141326 682718 141562 682954
rect 141646 682718 141882 682954
rect 141326 682398 141562 682634
rect 141646 682398 141882 682634
rect 141326 646718 141562 646954
rect 141646 646718 141882 646954
rect 141326 646398 141562 646634
rect 141646 646398 141882 646634
rect 141326 610718 141562 610954
rect 141646 610718 141882 610954
rect 141326 610398 141562 610634
rect 141646 610398 141882 610634
rect 141326 574718 141562 574954
rect 141646 574718 141882 574954
rect 141326 574398 141562 574634
rect 141646 574398 141882 574634
rect 141326 538718 141562 538954
rect 141646 538718 141882 538954
rect 141326 538398 141562 538634
rect 141646 538398 141882 538634
rect 141326 502718 141562 502954
rect 141646 502718 141882 502954
rect 141326 502398 141562 502634
rect 141646 502398 141882 502634
rect 141326 466718 141562 466954
rect 141646 466718 141882 466954
rect 141326 466398 141562 466634
rect 141646 466398 141882 466634
rect 141326 430718 141562 430954
rect 141646 430718 141882 430954
rect 141326 430398 141562 430634
rect 141646 430398 141882 430634
rect 141326 394718 141562 394954
rect 141646 394718 141882 394954
rect 141326 394398 141562 394634
rect 141646 394398 141882 394634
rect 141326 358718 141562 358954
rect 141646 358718 141882 358954
rect 141326 358398 141562 358634
rect 141646 358398 141882 358634
rect 141326 322718 141562 322954
rect 141646 322718 141882 322954
rect 141326 322398 141562 322634
rect 141646 322398 141882 322634
rect 141326 286718 141562 286954
rect 141646 286718 141882 286954
rect 141326 286398 141562 286634
rect 141646 286398 141882 286634
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 150326 705562 150562 705798
rect 150646 705562 150882 705798
rect 150326 705242 150562 705478
rect 150646 705242 150882 705478
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 150326 655718 150562 655954
rect 150646 655718 150882 655954
rect 150326 655398 150562 655634
rect 150646 655398 150882 655634
rect 150326 619718 150562 619954
rect 150646 619718 150882 619954
rect 150326 619398 150562 619634
rect 150646 619398 150882 619634
rect 150326 583718 150562 583954
rect 150646 583718 150882 583954
rect 150326 583398 150562 583634
rect 150646 583398 150882 583634
rect 150326 547718 150562 547954
rect 150646 547718 150882 547954
rect 150326 547398 150562 547634
rect 150646 547398 150882 547634
rect 150326 511718 150562 511954
rect 150646 511718 150882 511954
rect 150326 511398 150562 511634
rect 150646 511398 150882 511634
rect 150326 475718 150562 475954
rect 150646 475718 150882 475954
rect 150326 475398 150562 475634
rect 150646 475398 150882 475634
rect 150326 439718 150562 439954
rect 150646 439718 150882 439954
rect 150326 439398 150562 439634
rect 150646 439398 150882 439634
rect 150326 403718 150562 403954
rect 150646 403718 150882 403954
rect 150326 403398 150562 403634
rect 150646 403398 150882 403634
rect 150326 367718 150562 367954
rect 150646 367718 150882 367954
rect 150326 367398 150562 367634
rect 150646 367398 150882 367634
rect 150326 331718 150562 331954
rect 150646 331718 150882 331954
rect 150326 331398 150562 331634
rect 150646 331398 150882 331634
rect 150326 295718 150562 295954
rect 150646 295718 150882 295954
rect 150326 295398 150562 295634
rect 150646 295398 150882 295634
rect 154826 706522 155062 706758
rect 155146 706522 155382 706758
rect 154826 706202 155062 706438
rect 155146 706202 155382 706438
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 154826 660218 155062 660454
rect 155146 660218 155382 660454
rect 154826 659898 155062 660134
rect 155146 659898 155382 660134
rect 154826 624218 155062 624454
rect 155146 624218 155382 624454
rect 154826 623898 155062 624134
rect 155146 623898 155382 624134
rect 154826 588218 155062 588454
rect 155146 588218 155382 588454
rect 154826 587898 155062 588134
rect 155146 587898 155382 588134
rect 154826 552218 155062 552454
rect 155146 552218 155382 552454
rect 154826 551898 155062 552134
rect 155146 551898 155382 552134
rect 154826 516218 155062 516454
rect 155146 516218 155382 516454
rect 154826 515898 155062 516134
rect 155146 515898 155382 516134
rect 154826 480218 155062 480454
rect 155146 480218 155382 480454
rect 154826 479898 155062 480134
rect 155146 479898 155382 480134
rect 154826 444218 155062 444454
rect 155146 444218 155382 444454
rect 154826 443898 155062 444134
rect 155146 443898 155382 444134
rect 154826 408218 155062 408454
rect 155146 408218 155382 408454
rect 154826 407898 155062 408134
rect 155146 407898 155382 408134
rect 154826 372218 155062 372454
rect 155146 372218 155382 372454
rect 154826 371898 155062 372134
rect 155146 371898 155382 372134
rect 154826 336218 155062 336454
rect 155146 336218 155382 336454
rect 154826 335898 155062 336134
rect 155146 335898 155382 336134
rect 154826 300218 155062 300454
rect 155146 300218 155382 300454
rect 154826 299898 155062 300134
rect 155146 299898 155382 300134
rect 154826 264218 155062 264454
rect 155146 264218 155382 264454
rect 154826 263898 155062 264134
rect 155146 263898 155382 264134
rect 159326 707482 159562 707718
rect 159646 707482 159882 707718
rect 159326 707162 159562 707398
rect 159646 707162 159882 707398
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 159326 664718 159562 664954
rect 159646 664718 159882 664954
rect 159326 664398 159562 664634
rect 159646 664398 159882 664634
rect 159326 628718 159562 628954
rect 159646 628718 159882 628954
rect 159326 628398 159562 628634
rect 159646 628398 159882 628634
rect 159326 592718 159562 592954
rect 159646 592718 159882 592954
rect 159326 592398 159562 592634
rect 159646 592398 159882 592634
rect 159326 556718 159562 556954
rect 159646 556718 159882 556954
rect 159326 556398 159562 556634
rect 159646 556398 159882 556634
rect 159326 520718 159562 520954
rect 159646 520718 159882 520954
rect 159326 520398 159562 520634
rect 159646 520398 159882 520634
rect 159326 484718 159562 484954
rect 159646 484718 159882 484954
rect 159326 484398 159562 484634
rect 159646 484398 159882 484634
rect 159326 448718 159562 448954
rect 159646 448718 159882 448954
rect 159326 448398 159562 448634
rect 159646 448398 159882 448634
rect 159326 412718 159562 412954
rect 159646 412718 159882 412954
rect 159326 412398 159562 412634
rect 159646 412398 159882 412634
rect 159326 376718 159562 376954
rect 159646 376718 159882 376954
rect 159326 376398 159562 376634
rect 159646 376398 159882 376634
rect 159326 340718 159562 340954
rect 159646 340718 159882 340954
rect 159326 340398 159562 340634
rect 159646 340398 159882 340634
rect 159326 304718 159562 304954
rect 159646 304718 159882 304954
rect 159326 304398 159562 304634
rect 159646 304398 159882 304634
rect 159326 268718 159562 268954
rect 159646 268718 159882 268954
rect 159326 268398 159562 268634
rect 159646 268398 159882 268634
rect 163826 708442 164062 708678
rect 164146 708442 164382 708678
rect 163826 708122 164062 708358
rect 164146 708122 164382 708358
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 168326 709402 168562 709638
rect 168646 709402 168882 709638
rect 168326 709082 168562 709318
rect 168646 709082 168882 709318
rect 168326 673718 168562 673954
rect 168646 673718 168882 673954
rect 168326 673398 168562 673634
rect 168646 673398 168882 673634
rect 168326 637718 168562 637954
rect 168646 637718 168882 637954
rect 168326 637398 168562 637634
rect 168646 637398 168882 637634
rect 168326 601718 168562 601954
rect 168646 601718 168882 601954
rect 168326 601398 168562 601634
rect 168646 601398 168882 601634
rect 168326 565718 168562 565954
rect 168646 565718 168882 565954
rect 168326 565398 168562 565634
rect 168646 565398 168882 565634
rect 168326 529718 168562 529954
rect 168646 529718 168882 529954
rect 168326 529398 168562 529634
rect 168646 529398 168882 529634
rect 168326 493718 168562 493954
rect 168646 493718 168882 493954
rect 168326 493398 168562 493634
rect 168646 493398 168882 493634
rect 168326 457718 168562 457954
rect 168646 457718 168882 457954
rect 168326 457398 168562 457634
rect 168646 457398 168882 457634
rect 168326 421718 168562 421954
rect 168646 421718 168882 421954
rect 168326 421398 168562 421634
rect 168646 421398 168882 421634
rect 168326 385718 168562 385954
rect 168646 385718 168882 385954
rect 168326 385398 168562 385634
rect 168646 385398 168882 385634
rect 168326 349718 168562 349954
rect 168646 349718 168882 349954
rect 168326 349398 168562 349634
rect 168646 349398 168882 349634
rect 168326 313718 168562 313954
rect 168646 313718 168882 313954
rect 168326 313398 168562 313634
rect 168646 313398 168882 313634
rect 168326 277718 168562 277954
rect 168646 277718 168882 277954
rect 168326 277398 168562 277634
rect 168646 277398 168882 277634
rect 172826 710362 173062 710598
rect 173146 710362 173382 710598
rect 172826 710042 173062 710278
rect 173146 710042 173382 710278
rect 172826 678218 173062 678454
rect 173146 678218 173382 678454
rect 172826 677898 173062 678134
rect 173146 677898 173382 678134
rect 172826 642218 173062 642454
rect 173146 642218 173382 642454
rect 172826 641898 173062 642134
rect 173146 641898 173382 642134
rect 172826 606218 173062 606454
rect 173146 606218 173382 606454
rect 172826 605898 173062 606134
rect 173146 605898 173382 606134
rect 172826 570218 173062 570454
rect 173146 570218 173382 570454
rect 172826 569898 173062 570134
rect 173146 569898 173382 570134
rect 172826 534218 173062 534454
rect 173146 534218 173382 534454
rect 172826 533898 173062 534134
rect 173146 533898 173382 534134
rect 172826 498218 173062 498454
rect 173146 498218 173382 498454
rect 172826 497898 173062 498134
rect 173146 497898 173382 498134
rect 172826 462218 173062 462454
rect 173146 462218 173382 462454
rect 172826 461898 173062 462134
rect 173146 461898 173382 462134
rect 172826 426218 173062 426454
rect 173146 426218 173382 426454
rect 172826 425898 173062 426134
rect 173146 425898 173382 426134
rect 172826 390218 173062 390454
rect 173146 390218 173382 390454
rect 172826 389898 173062 390134
rect 173146 389898 173382 390134
rect 172826 354218 173062 354454
rect 173146 354218 173382 354454
rect 172826 353898 173062 354134
rect 173146 353898 173382 354134
rect 172826 318218 173062 318454
rect 173146 318218 173382 318454
rect 172826 317898 173062 318134
rect 173146 317898 173382 318134
rect 172826 282218 173062 282454
rect 173146 282218 173382 282454
rect 172826 281898 173062 282134
rect 173146 281898 173382 282134
rect 177326 711322 177562 711558
rect 177646 711322 177882 711558
rect 177326 711002 177562 711238
rect 177646 711002 177882 711238
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 177326 646718 177562 646954
rect 177646 646718 177882 646954
rect 177326 646398 177562 646634
rect 177646 646398 177882 646634
rect 177326 610718 177562 610954
rect 177646 610718 177882 610954
rect 177326 610398 177562 610634
rect 177646 610398 177882 610634
rect 177326 574718 177562 574954
rect 177646 574718 177882 574954
rect 177326 574398 177562 574634
rect 177646 574398 177882 574634
rect 177326 538718 177562 538954
rect 177646 538718 177882 538954
rect 177326 538398 177562 538634
rect 177646 538398 177882 538634
rect 177326 502718 177562 502954
rect 177646 502718 177882 502954
rect 177326 502398 177562 502634
rect 177646 502398 177882 502634
rect 177326 466718 177562 466954
rect 177646 466718 177882 466954
rect 177326 466398 177562 466634
rect 177646 466398 177882 466634
rect 177326 430718 177562 430954
rect 177646 430718 177882 430954
rect 177326 430398 177562 430634
rect 177646 430398 177882 430634
rect 177326 394718 177562 394954
rect 177646 394718 177882 394954
rect 177326 394398 177562 394634
rect 177646 394398 177882 394634
rect 177326 358718 177562 358954
rect 177646 358718 177882 358954
rect 177326 358398 177562 358634
rect 177646 358398 177882 358634
rect 177326 322718 177562 322954
rect 177646 322718 177882 322954
rect 177326 322398 177562 322634
rect 177646 322398 177882 322634
rect 177326 286718 177562 286954
rect 177646 286718 177882 286954
rect 177326 286398 177562 286634
rect 177646 286398 177882 286634
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 186326 705562 186562 705798
rect 186646 705562 186882 705798
rect 186326 705242 186562 705478
rect 186646 705242 186882 705478
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 186326 655718 186562 655954
rect 186646 655718 186882 655954
rect 186326 655398 186562 655634
rect 186646 655398 186882 655634
rect 186326 619718 186562 619954
rect 186646 619718 186882 619954
rect 186326 619398 186562 619634
rect 186646 619398 186882 619634
rect 186326 583718 186562 583954
rect 186646 583718 186882 583954
rect 186326 583398 186562 583634
rect 186646 583398 186882 583634
rect 186326 547718 186562 547954
rect 186646 547718 186882 547954
rect 186326 547398 186562 547634
rect 186646 547398 186882 547634
rect 186326 511718 186562 511954
rect 186646 511718 186882 511954
rect 186326 511398 186562 511634
rect 186646 511398 186882 511634
rect 186326 475718 186562 475954
rect 186646 475718 186882 475954
rect 186326 475398 186562 475634
rect 186646 475398 186882 475634
rect 186326 439718 186562 439954
rect 186646 439718 186882 439954
rect 186326 439398 186562 439634
rect 186646 439398 186882 439634
rect 186326 403718 186562 403954
rect 186646 403718 186882 403954
rect 186326 403398 186562 403634
rect 186646 403398 186882 403634
rect 186326 367718 186562 367954
rect 186646 367718 186882 367954
rect 186326 367398 186562 367634
rect 186646 367398 186882 367634
rect 186326 331718 186562 331954
rect 186646 331718 186882 331954
rect 186326 331398 186562 331634
rect 186646 331398 186882 331634
rect 186326 295718 186562 295954
rect 186646 295718 186882 295954
rect 186326 295398 186562 295634
rect 186646 295398 186882 295634
rect 190826 706522 191062 706758
rect 191146 706522 191382 706758
rect 190826 706202 191062 706438
rect 191146 706202 191382 706438
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 190826 660218 191062 660454
rect 191146 660218 191382 660454
rect 190826 659898 191062 660134
rect 191146 659898 191382 660134
rect 190826 624218 191062 624454
rect 191146 624218 191382 624454
rect 190826 623898 191062 624134
rect 191146 623898 191382 624134
rect 190826 588218 191062 588454
rect 191146 588218 191382 588454
rect 190826 587898 191062 588134
rect 191146 587898 191382 588134
rect 190826 552218 191062 552454
rect 191146 552218 191382 552454
rect 190826 551898 191062 552134
rect 191146 551898 191382 552134
rect 190826 516218 191062 516454
rect 191146 516218 191382 516454
rect 190826 515898 191062 516134
rect 191146 515898 191382 516134
rect 190826 480218 191062 480454
rect 191146 480218 191382 480454
rect 190826 479898 191062 480134
rect 191146 479898 191382 480134
rect 190826 444218 191062 444454
rect 191146 444218 191382 444454
rect 190826 443898 191062 444134
rect 191146 443898 191382 444134
rect 190826 408218 191062 408454
rect 191146 408218 191382 408454
rect 190826 407898 191062 408134
rect 191146 407898 191382 408134
rect 190826 372218 191062 372454
rect 191146 372218 191382 372454
rect 190826 371898 191062 372134
rect 191146 371898 191382 372134
rect 190826 336218 191062 336454
rect 191146 336218 191382 336454
rect 190826 335898 191062 336134
rect 191146 335898 191382 336134
rect 190826 300218 191062 300454
rect 191146 300218 191382 300454
rect 190826 299898 191062 300134
rect 191146 299898 191382 300134
rect 124250 255218 124486 255454
rect 124250 254898 124486 255134
rect 154970 255218 155206 255454
rect 154970 254898 155206 255134
rect 185690 255218 185926 255454
rect 185690 254898 185926 255134
rect 139610 223718 139846 223954
rect 139610 223398 139846 223634
rect 170330 223718 170566 223954
rect 170330 223398 170566 223634
rect 124250 219218 124486 219454
rect 124250 218898 124486 219134
rect 154970 219218 155206 219454
rect 154970 218898 155206 219134
rect 185690 219218 185926 219454
rect 185690 218898 185926 219134
rect 123326 196718 123562 196954
rect 123646 196718 123882 196954
rect 123326 196398 123562 196634
rect 123646 196398 123882 196634
rect 123326 160718 123562 160954
rect 123646 160718 123882 160954
rect 123326 160398 123562 160634
rect 123646 160398 123882 160634
rect 141326 178718 141562 178954
rect 141646 178718 141882 178954
rect 141326 178398 141562 178634
rect 141646 178398 141882 178634
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 141326 142718 141562 142954
rect 141646 142718 141882 142954
rect 141326 142398 141562 142634
rect 141646 142398 141882 142634
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1542 114562 -1306
rect 114646 -1542 114882 -1306
rect 114326 -1862 114562 -1626
rect 114646 -1862 114882 -1626
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2502 119062 -2266
rect 119146 -2502 119382 -2266
rect 118826 -2822 119062 -2586
rect 119146 -2822 119382 -2586
rect 150326 187718 150562 187954
rect 150646 187718 150882 187954
rect 150326 187398 150562 187634
rect 150646 187398 150882 187634
rect 150326 151718 150562 151954
rect 150646 151718 150882 151954
rect 150326 151398 150562 151634
rect 150646 151398 150882 151634
rect 154826 192218 155062 192454
rect 155146 192218 155382 192454
rect 154826 191898 155062 192134
rect 155146 191898 155382 192134
rect 154826 156218 155062 156454
rect 155146 156218 155382 156454
rect 154826 155898 155062 156134
rect 155146 155898 155382 156134
rect 159326 196718 159562 196954
rect 159646 196718 159882 196954
rect 159326 196398 159562 196634
rect 159646 196398 159882 196634
rect 159326 160718 159562 160954
rect 159646 160718 159882 160954
rect 159326 160398 159562 160634
rect 159646 160398 159882 160634
rect 177326 178718 177562 178954
rect 177646 178718 177882 178954
rect 177326 178398 177562 178634
rect 177646 178398 177882 178634
rect 177326 142718 177562 142954
rect 177646 142718 177882 142954
rect 177326 142398 177562 142634
rect 177646 142398 177882 142634
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 139610 115718 139846 115954
rect 139610 115398 139846 115634
rect 170330 115718 170566 115954
rect 170330 115398 170566 115634
rect 124250 111218 124486 111454
rect 124250 110898 124486 111134
rect 154970 111218 155206 111454
rect 154970 110898 155206 111134
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 123326 -3462 123562 -3226
rect 123646 -3462 123882 -3226
rect 123326 -3782 123562 -3546
rect 123646 -3782 123882 -3546
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -4422 128062 -4186
rect 128146 -4422 128382 -4186
rect 127826 -4742 128062 -4506
rect 128146 -4742 128382 -4506
rect 132326 61718 132562 61954
rect 132646 61718 132882 61954
rect 132326 61398 132562 61634
rect 132646 61398 132882 61634
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 132326 -5382 132562 -5146
rect 132646 -5382 132882 -5146
rect 132326 -5702 132562 -5466
rect 132646 -5702 132882 -5466
rect 141326 70718 141562 70954
rect 141646 70718 141882 70954
rect 141326 70398 141562 70634
rect 141646 70398 141882 70634
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 136826 -6342 137062 -6106
rect 137146 -6342 137382 -6106
rect 136826 -6662 137062 -6426
rect 137146 -6662 137382 -6426
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 141326 -7302 141562 -7066
rect 141646 -7302 141882 -7066
rect 141326 -7622 141562 -7386
rect 141646 -7622 141882 -7386
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 150326 -1542 150562 -1306
rect 150646 -1542 150882 -1306
rect 150326 -1862 150562 -1626
rect 150646 -1862 150882 -1626
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 154826 -2502 155062 -2266
rect 155146 -2502 155382 -2266
rect 154826 -2822 155062 -2586
rect 155146 -2822 155382 -2586
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 159326 -3462 159562 -3226
rect 159646 -3462 159882 -3226
rect 159326 -3782 159562 -3546
rect 159646 -3782 159882 -3546
rect 168326 61718 168562 61954
rect 168646 61718 168882 61954
rect 168326 61398 168562 61634
rect 168646 61398 168882 61634
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -4422 164062 -4186
rect 164146 -4422 164382 -4186
rect 163826 -4742 164062 -4506
rect 164146 -4742 164382 -4506
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 168326 -5382 168562 -5146
rect 168646 -5382 168882 -5146
rect 168326 -5702 168562 -5466
rect 168646 -5702 168882 -5466
rect 177326 70718 177562 70954
rect 177646 70718 177882 70954
rect 177326 70398 177562 70634
rect 177646 70398 177882 70634
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 172826 -6342 173062 -6106
rect 173146 -6342 173382 -6106
rect 172826 -6662 173062 -6426
rect 173146 -6662 173382 -6426
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 177326 -7302 177562 -7066
rect 177646 -7302 177882 -7066
rect 177326 -7622 177562 -7386
rect 177646 -7622 177882 -7386
rect 185690 111218 185926 111454
rect 185690 110898 185926 111134
rect 186326 187718 186562 187954
rect 186646 187718 186882 187954
rect 186326 187398 186562 187634
rect 186646 187398 186882 187634
rect 186326 151718 186562 151954
rect 186646 151718 186882 151954
rect 186326 151398 186562 151634
rect 186646 151398 186882 151634
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 190826 264218 191062 264454
rect 191146 264218 191382 264454
rect 190826 263898 191062 264134
rect 191146 263898 191382 264134
rect 195326 707482 195562 707718
rect 195646 707482 195882 707718
rect 195326 707162 195562 707398
rect 195646 707162 195882 707398
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 195326 664718 195562 664954
rect 195646 664718 195882 664954
rect 195326 664398 195562 664634
rect 195646 664398 195882 664634
rect 195326 628718 195562 628954
rect 195646 628718 195882 628954
rect 195326 628398 195562 628634
rect 195646 628398 195882 628634
rect 195326 592718 195562 592954
rect 195646 592718 195882 592954
rect 195326 592398 195562 592634
rect 195646 592398 195882 592634
rect 195326 556718 195562 556954
rect 195646 556718 195882 556954
rect 195326 556398 195562 556634
rect 195646 556398 195882 556634
rect 195326 520718 195562 520954
rect 195646 520718 195882 520954
rect 195326 520398 195562 520634
rect 195646 520398 195882 520634
rect 195326 484718 195562 484954
rect 195646 484718 195882 484954
rect 195326 484398 195562 484634
rect 195646 484398 195882 484634
rect 195326 448718 195562 448954
rect 195646 448718 195882 448954
rect 195326 448398 195562 448634
rect 195646 448398 195882 448634
rect 195326 412718 195562 412954
rect 195646 412718 195882 412954
rect 195326 412398 195562 412634
rect 195646 412398 195882 412634
rect 195326 376718 195562 376954
rect 195646 376718 195882 376954
rect 195326 376398 195562 376634
rect 195646 376398 195882 376634
rect 195326 340718 195562 340954
rect 195646 340718 195882 340954
rect 195326 340398 195562 340634
rect 195646 340398 195882 340634
rect 195326 304718 195562 304954
rect 195646 304718 195882 304954
rect 195326 304398 195562 304634
rect 195646 304398 195882 304634
rect 195326 268718 195562 268954
rect 195646 268718 195882 268954
rect 195326 268398 195562 268634
rect 195646 268398 195882 268634
rect 190826 192218 191062 192454
rect 191146 192218 191382 192454
rect 190826 191898 191062 192134
rect 191146 191898 191382 192134
rect 190826 156218 191062 156454
rect 191146 156218 191382 156454
rect 190826 155898 191062 156134
rect 191146 155898 191382 156134
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1542 186562 -1306
rect 186646 -1542 186882 -1306
rect 186326 -1862 186562 -1626
rect 186646 -1862 186882 -1626
rect 199826 708442 200062 708678
rect 200146 708442 200382 708678
rect 199826 708122 200062 708358
rect 200146 708122 200382 708358
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 195326 232718 195562 232954
rect 195646 232718 195882 232954
rect 195326 232398 195562 232634
rect 195646 232398 195882 232634
rect 195326 196718 195562 196954
rect 195646 196718 195882 196954
rect 195326 196398 195562 196634
rect 195646 196398 195882 196634
rect 195326 160718 195562 160954
rect 195646 160718 195882 160954
rect 195326 160398 195562 160634
rect 195646 160398 195882 160634
rect 195326 124718 195562 124954
rect 195646 124718 195882 124954
rect 195326 124398 195562 124634
rect 195646 124398 195882 124634
rect 195326 88718 195562 88954
rect 195646 88718 195882 88954
rect 195326 88398 195562 88634
rect 195646 88398 195882 88634
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2502 191062 -2266
rect 191146 -2502 191382 -2266
rect 190826 -2822 191062 -2586
rect 191146 -2822 191382 -2586
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 204326 709402 204562 709638
rect 204646 709402 204882 709638
rect 204326 709082 204562 709318
rect 204646 709082 204882 709318
rect 204326 673718 204562 673954
rect 204646 673718 204882 673954
rect 204326 673398 204562 673634
rect 204646 673398 204882 673634
rect 204326 637718 204562 637954
rect 204646 637718 204882 637954
rect 204326 637398 204562 637634
rect 204646 637398 204882 637634
rect 204326 601718 204562 601954
rect 204646 601718 204882 601954
rect 204326 601398 204562 601634
rect 204646 601398 204882 601634
rect 204326 565718 204562 565954
rect 204646 565718 204882 565954
rect 204326 565398 204562 565634
rect 204646 565398 204882 565634
rect 204326 529718 204562 529954
rect 204646 529718 204882 529954
rect 204326 529398 204562 529634
rect 204646 529398 204882 529634
rect 204326 493718 204562 493954
rect 204646 493718 204882 493954
rect 204326 493398 204562 493634
rect 204646 493398 204882 493634
rect 204326 457718 204562 457954
rect 204646 457718 204882 457954
rect 204326 457398 204562 457634
rect 204646 457398 204882 457634
rect 204326 421718 204562 421954
rect 204646 421718 204882 421954
rect 204326 421398 204562 421634
rect 204646 421398 204882 421634
rect 204326 385718 204562 385954
rect 204646 385718 204882 385954
rect 204326 385398 204562 385634
rect 204646 385398 204882 385634
rect 204326 349718 204562 349954
rect 204646 349718 204882 349954
rect 204326 349398 204562 349634
rect 204646 349398 204882 349634
rect 204326 313718 204562 313954
rect 204646 313718 204882 313954
rect 204326 313398 204562 313634
rect 204646 313398 204882 313634
rect 204326 277718 204562 277954
rect 204646 277718 204882 277954
rect 204326 277398 204562 277634
rect 204646 277398 204882 277634
rect 204326 241718 204562 241954
rect 204646 241718 204882 241954
rect 204326 241398 204562 241634
rect 204646 241398 204882 241634
rect 204326 205718 204562 205954
rect 204646 205718 204882 205954
rect 204326 205398 204562 205634
rect 204646 205398 204882 205634
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3462 195562 -3226
rect 195646 -3462 195882 -3226
rect 195326 -3782 195562 -3546
rect 195646 -3782 195882 -3546
rect 208826 710362 209062 710598
rect 209146 710362 209382 710598
rect 208826 710042 209062 710278
rect 209146 710042 209382 710278
rect 208826 678218 209062 678454
rect 209146 678218 209382 678454
rect 208826 677898 209062 678134
rect 209146 677898 209382 678134
rect 208826 642218 209062 642454
rect 209146 642218 209382 642454
rect 208826 641898 209062 642134
rect 209146 641898 209382 642134
rect 208826 606218 209062 606454
rect 209146 606218 209382 606454
rect 208826 605898 209062 606134
rect 209146 605898 209382 606134
rect 208826 570218 209062 570454
rect 209146 570218 209382 570454
rect 208826 569898 209062 570134
rect 209146 569898 209382 570134
rect 208826 534218 209062 534454
rect 209146 534218 209382 534454
rect 208826 533898 209062 534134
rect 209146 533898 209382 534134
rect 208826 498218 209062 498454
rect 209146 498218 209382 498454
rect 208826 497898 209062 498134
rect 209146 497898 209382 498134
rect 208826 462218 209062 462454
rect 209146 462218 209382 462454
rect 208826 461898 209062 462134
rect 209146 461898 209382 462134
rect 208826 426218 209062 426454
rect 209146 426218 209382 426454
rect 208826 425898 209062 426134
rect 209146 425898 209382 426134
rect 208826 390218 209062 390454
rect 209146 390218 209382 390454
rect 208826 389898 209062 390134
rect 209146 389898 209382 390134
rect 208826 354218 209062 354454
rect 209146 354218 209382 354454
rect 208826 353898 209062 354134
rect 209146 353898 209382 354134
rect 208826 318218 209062 318454
rect 209146 318218 209382 318454
rect 208826 317898 209062 318134
rect 209146 317898 209382 318134
rect 208826 282218 209062 282454
rect 209146 282218 209382 282454
rect 208826 281898 209062 282134
rect 209146 281898 209382 282134
rect 208826 246218 209062 246454
rect 209146 246218 209382 246454
rect 208826 245898 209062 246134
rect 209146 245898 209382 246134
rect 208826 210218 209062 210454
rect 209146 210218 209382 210454
rect 208826 209898 209062 210134
rect 209146 209898 209382 210134
rect 204326 169718 204562 169954
rect 204646 169718 204882 169954
rect 204326 169398 204562 169634
rect 204646 169398 204882 169634
rect 204326 133718 204562 133954
rect 204646 133718 204882 133954
rect 204326 133398 204562 133634
rect 204646 133398 204882 133634
rect 204326 97718 204562 97954
rect 204646 97718 204882 97954
rect 204326 97398 204562 97634
rect 204646 97398 204882 97634
rect 204326 61718 204562 61954
rect 204646 61718 204882 61954
rect 204326 61398 204562 61634
rect 204646 61398 204882 61634
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4422 200062 -4186
rect 200146 -4422 200382 -4186
rect 199826 -4742 200062 -4506
rect 200146 -4742 200382 -4506
rect 213326 711322 213562 711558
rect 213646 711322 213882 711558
rect 213326 711002 213562 711238
rect 213646 711002 213882 711238
rect 213326 682718 213562 682954
rect 213646 682718 213882 682954
rect 213326 682398 213562 682634
rect 213646 682398 213882 682634
rect 213326 646718 213562 646954
rect 213646 646718 213882 646954
rect 213326 646398 213562 646634
rect 213646 646398 213882 646634
rect 213326 610718 213562 610954
rect 213646 610718 213882 610954
rect 213326 610398 213562 610634
rect 213646 610398 213882 610634
rect 213326 574718 213562 574954
rect 213646 574718 213882 574954
rect 213326 574398 213562 574634
rect 213646 574398 213882 574634
rect 213326 538718 213562 538954
rect 213646 538718 213882 538954
rect 213326 538398 213562 538634
rect 213646 538398 213882 538634
rect 213326 502718 213562 502954
rect 213646 502718 213882 502954
rect 213326 502398 213562 502634
rect 213646 502398 213882 502634
rect 213326 466718 213562 466954
rect 213646 466718 213882 466954
rect 213326 466398 213562 466634
rect 213646 466398 213882 466634
rect 213326 430718 213562 430954
rect 213646 430718 213882 430954
rect 213326 430398 213562 430634
rect 213646 430398 213882 430634
rect 213326 394718 213562 394954
rect 213646 394718 213882 394954
rect 213326 394398 213562 394634
rect 213646 394398 213882 394634
rect 213326 358718 213562 358954
rect 213646 358718 213882 358954
rect 213326 358398 213562 358634
rect 213646 358398 213882 358634
rect 213326 322718 213562 322954
rect 213646 322718 213882 322954
rect 213326 322398 213562 322634
rect 213646 322398 213882 322634
rect 213326 286718 213562 286954
rect 213646 286718 213882 286954
rect 213326 286398 213562 286634
rect 213646 286398 213882 286634
rect 213326 250718 213562 250954
rect 213646 250718 213882 250954
rect 213326 250398 213562 250634
rect 213646 250398 213882 250634
rect 213326 214718 213562 214954
rect 213646 214718 213882 214954
rect 213326 214398 213562 214634
rect 213646 214398 213882 214634
rect 208826 174218 209062 174454
rect 209146 174218 209382 174454
rect 208826 173898 209062 174134
rect 209146 173898 209382 174134
rect 208826 138218 209062 138454
rect 209146 138218 209382 138454
rect 208826 137898 209062 138134
rect 209146 137898 209382 138134
rect 208826 102218 209062 102454
rect 209146 102218 209382 102454
rect 208826 101898 209062 102134
rect 209146 101898 209382 102134
rect 208826 66218 209062 66454
rect 209146 66218 209382 66454
rect 208826 65898 209062 66134
rect 209146 65898 209382 66134
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 204326 -5382 204562 -5146
rect 204646 -5382 204882 -5146
rect 204326 -5702 204562 -5466
rect 204646 -5702 204882 -5466
rect 213326 178718 213562 178954
rect 213646 178718 213882 178954
rect 213326 178398 213562 178634
rect 213646 178398 213882 178634
rect 213326 142718 213562 142954
rect 213646 142718 213882 142954
rect 213326 142398 213562 142634
rect 213646 142398 213882 142634
rect 213326 106718 213562 106954
rect 213646 106718 213882 106954
rect 213326 106398 213562 106634
rect 213646 106398 213882 106634
rect 213326 70718 213562 70954
rect 213646 70718 213882 70954
rect 213326 70398 213562 70634
rect 213646 70398 213882 70634
rect 208826 30218 209062 30454
rect 209146 30218 209382 30454
rect 208826 29898 209062 30134
rect 209146 29898 209382 30134
rect 208826 -6342 209062 -6106
rect 209146 -6342 209382 -6106
rect 208826 -6662 209062 -6426
rect 209146 -6662 209382 -6426
rect 213326 34718 213562 34954
rect 213646 34718 213882 34954
rect 213326 34398 213562 34634
rect 213646 34398 213882 34634
rect 213326 -7302 213562 -7066
rect 213646 -7302 213882 -7066
rect 213326 -7622 213562 -7386
rect 213646 -7622 213882 -7386
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 222326 705562 222562 705798
rect 222646 705562 222882 705798
rect 222326 705242 222562 705478
rect 222646 705242 222882 705478
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 222326 655718 222562 655954
rect 222646 655718 222882 655954
rect 222326 655398 222562 655634
rect 222646 655398 222882 655634
rect 222326 619718 222562 619954
rect 222646 619718 222882 619954
rect 222326 619398 222562 619634
rect 222646 619398 222882 619634
rect 222326 583718 222562 583954
rect 222646 583718 222882 583954
rect 222326 583398 222562 583634
rect 222646 583398 222882 583634
rect 222326 547718 222562 547954
rect 222646 547718 222882 547954
rect 222326 547398 222562 547634
rect 222646 547398 222882 547634
rect 222326 511718 222562 511954
rect 222646 511718 222882 511954
rect 222326 511398 222562 511634
rect 222646 511398 222882 511634
rect 222326 475718 222562 475954
rect 222646 475718 222882 475954
rect 222326 475398 222562 475634
rect 222646 475398 222882 475634
rect 222326 439718 222562 439954
rect 222646 439718 222882 439954
rect 222326 439398 222562 439634
rect 222646 439398 222882 439634
rect 222326 403718 222562 403954
rect 222646 403718 222882 403954
rect 222326 403398 222562 403634
rect 222646 403398 222882 403634
rect 222326 367718 222562 367954
rect 222646 367718 222882 367954
rect 222326 367398 222562 367634
rect 222646 367398 222882 367634
rect 222326 331718 222562 331954
rect 222646 331718 222882 331954
rect 222326 331398 222562 331634
rect 222646 331398 222882 331634
rect 222326 295718 222562 295954
rect 222646 295718 222882 295954
rect 222326 295398 222562 295634
rect 222646 295398 222882 295634
rect 222326 259718 222562 259954
rect 222646 259718 222882 259954
rect 222326 259398 222562 259634
rect 222646 259398 222882 259634
rect 222326 223718 222562 223954
rect 222646 223718 222882 223954
rect 222326 223398 222562 223634
rect 222646 223398 222882 223634
rect 222326 187718 222562 187954
rect 222646 187718 222882 187954
rect 222326 187398 222562 187634
rect 222646 187398 222882 187634
rect 222326 151718 222562 151954
rect 222646 151718 222882 151954
rect 222326 151398 222562 151634
rect 222646 151398 222882 151634
rect 222326 115718 222562 115954
rect 222646 115718 222882 115954
rect 222326 115398 222562 115634
rect 222646 115398 222882 115634
rect 222326 79718 222562 79954
rect 222646 79718 222882 79954
rect 222326 79398 222562 79634
rect 222646 79398 222882 79634
rect 222326 43718 222562 43954
rect 222646 43718 222882 43954
rect 222326 43398 222562 43634
rect 222646 43398 222882 43634
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 222326 -1542 222562 -1306
rect 222646 -1542 222882 -1306
rect 222326 -1862 222562 -1626
rect 222646 -1862 222882 -1626
rect 226826 706522 227062 706758
rect 227146 706522 227382 706758
rect 226826 706202 227062 706438
rect 227146 706202 227382 706438
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 226826 660218 227062 660454
rect 227146 660218 227382 660454
rect 226826 659898 227062 660134
rect 227146 659898 227382 660134
rect 226826 624218 227062 624454
rect 227146 624218 227382 624454
rect 226826 623898 227062 624134
rect 227146 623898 227382 624134
rect 226826 588218 227062 588454
rect 227146 588218 227382 588454
rect 226826 587898 227062 588134
rect 227146 587898 227382 588134
rect 226826 552218 227062 552454
rect 227146 552218 227382 552454
rect 226826 551898 227062 552134
rect 227146 551898 227382 552134
rect 226826 516218 227062 516454
rect 227146 516218 227382 516454
rect 226826 515898 227062 516134
rect 227146 515898 227382 516134
rect 226826 480218 227062 480454
rect 227146 480218 227382 480454
rect 226826 479898 227062 480134
rect 227146 479898 227382 480134
rect 226826 444218 227062 444454
rect 227146 444218 227382 444454
rect 226826 443898 227062 444134
rect 227146 443898 227382 444134
rect 226826 408218 227062 408454
rect 227146 408218 227382 408454
rect 226826 407898 227062 408134
rect 227146 407898 227382 408134
rect 226826 372218 227062 372454
rect 227146 372218 227382 372454
rect 226826 371898 227062 372134
rect 227146 371898 227382 372134
rect 226826 336218 227062 336454
rect 227146 336218 227382 336454
rect 226826 335898 227062 336134
rect 227146 335898 227382 336134
rect 226826 300218 227062 300454
rect 227146 300218 227382 300454
rect 226826 299898 227062 300134
rect 227146 299898 227382 300134
rect 226826 264218 227062 264454
rect 227146 264218 227382 264454
rect 226826 263898 227062 264134
rect 227146 263898 227382 264134
rect 226826 228218 227062 228454
rect 227146 228218 227382 228454
rect 226826 227898 227062 228134
rect 227146 227898 227382 228134
rect 226826 192218 227062 192454
rect 227146 192218 227382 192454
rect 226826 191898 227062 192134
rect 227146 191898 227382 192134
rect 226826 156218 227062 156454
rect 227146 156218 227382 156454
rect 226826 155898 227062 156134
rect 227146 155898 227382 156134
rect 226826 120218 227062 120454
rect 227146 120218 227382 120454
rect 226826 119898 227062 120134
rect 227146 119898 227382 120134
rect 226826 84218 227062 84454
rect 227146 84218 227382 84454
rect 226826 83898 227062 84134
rect 227146 83898 227382 84134
rect 226826 48218 227062 48454
rect 227146 48218 227382 48454
rect 226826 47898 227062 48134
rect 227146 47898 227382 48134
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2502 227062 -2266
rect 227146 -2502 227382 -2266
rect 226826 -2822 227062 -2586
rect 227146 -2822 227382 -2586
rect 231326 707482 231562 707718
rect 231646 707482 231882 707718
rect 231326 707162 231562 707398
rect 231646 707162 231882 707398
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 231326 664718 231562 664954
rect 231646 664718 231882 664954
rect 231326 664398 231562 664634
rect 231646 664398 231882 664634
rect 231326 628718 231562 628954
rect 231646 628718 231882 628954
rect 231326 628398 231562 628634
rect 231646 628398 231882 628634
rect 231326 592718 231562 592954
rect 231646 592718 231882 592954
rect 231326 592398 231562 592634
rect 231646 592398 231882 592634
rect 231326 556718 231562 556954
rect 231646 556718 231882 556954
rect 231326 556398 231562 556634
rect 231646 556398 231882 556634
rect 231326 520718 231562 520954
rect 231646 520718 231882 520954
rect 231326 520398 231562 520634
rect 231646 520398 231882 520634
rect 231326 484718 231562 484954
rect 231646 484718 231882 484954
rect 231326 484398 231562 484634
rect 231646 484398 231882 484634
rect 231326 448718 231562 448954
rect 231646 448718 231882 448954
rect 231326 448398 231562 448634
rect 231646 448398 231882 448634
rect 231326 412718 231562 412954
rect 231646 412718 231882 412954
rect 231326 412398 231562 412634
rect 231646 412398 231882 412634
rect 231326 376718 231562 376954
rect 231646 376718 231882 376954
rect 231326 376398 231562 376634
rect 231646 376398 231882 376634
rect 231326 340718 231562 340954
rect 231646 340718 231882 340954
rect 231326 340398 231562 340634
rect 231646 340398 231882 340634
rect 231326 304718 231562 304954
rect 231646 304718 231882 304954
rect 231326 304398 231562 304634
rect 231646 304398 231882 304634
rect 231326 268718 231562 268954
rect 231646 268718 231882 268954
rect 231326 268398 231562 268634
rect 231646 268398 231882 268634
rect 231326 232718 231562 232954
rect 231646 232718 231882 232954
rect 231326 232398 231562 232634
rect 231646 232398 231882 232634
rect 231326 196718 231562 196954
rect 231646 196718 231882 196954
rect 231326 196398 231562 196634
rect 231646 196398 231882 196634
rect 231326 160718 231562 160954
rect 231646 160718 231882 160954
rect 231326 160398 231562 160634
rect 231646 160398 231882 160634
rect 231326 124718 231562 124954
rect 231646 124718 231882 124954
rect 231326 124398 231562 124634
rect 231646 124398 231882 124634
rect 231326 88718 231562 88954
rect 231646 88718 231882 88954
rect 231326 88398 231562 88634
rect 231646 88398 231882 88634
rect 231326 52718 231562 52954
rect 231646 52718 231882 52954
rect 231326 52398 231562 52634
rect 231646 52398 231882 52634
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3462 231562 -3226
rect 231646 -3462 231882 -3226
rect 231326 -3782 231562 -3546
rect 231646 -3782 231882 -3546
rect 235826 708442 236062 708678
rect 236146 708442 236382 708678
rect 235826 708122 236062 708358
rect 236146 708122 236382 708358
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4422 236062 -4186
rect 236146 -4422 236382 -4186
rect 235826 -4742 236062 -4506
rect 236146 -4742 236382 -4506
rect 240326 709402 240562 709638
rect 240646 709402 240882 709638
rect 240326 709082 240562 709318
rect 240646 709082 240882 709318
rect 240326 673718 240562 673954
rect 240646 673718 240882 673954
rect 240326 673398 240562 673634
rect 240646 673398 240882 673634
rect 240326 637718 240562 637954
rect 240646 637718 240882 637954
rect 240326 637398 240562 637634
rect 240646 637398 240882 637634
rect 240326 601718 240562 601954
rect 240646 601718 240882 601954
rect 240326 601398 240562 601634
rect 240646 601398 240882 601634
rect 240326 565718 240562 565954
rect 240646 565718 240882 565954
rect 240326 565398 240562 565634
rect 240646 565398 240882 565634
rect 240326 529718 240562 529954
rect 240646 529718 240882 529954
rect 240326 529398 240562 529634
rect 240646 529398 240882 529634
rect 240326 493718 240562 493954
rect 240646 493718 240882 493954
rect 240326 493398 240562 493634
rect 240646 493398 240882 493634
rect 240326 457718 240562 457954
rect 240646 457718 240882 457954
rect 240326 457398 240562 457634
rect 240646 457398 240882 457634
rect 240326 421718 240562 421954
rect 240646 421718 240882 421954
rect 240326 421398 240562 421634
rect 240646 421398 240882 421634
rect 240326 385718 240562 385954
rect 240646 385718 240882 385954
rect 240326 385398 240562 385634
rect 240646 385398 240882 385634
rect 240326 349718 240562 349954
rect 240646 349718 240882 349954
rect 240326 349398 240562 349634
rect 240646 349398 240882 349634
rect 240326 313718 240562 313954
rect 240646 313718 240882 313954
rect 240326 313398 240562 313634
rect 240646 313398 240882 313634
rect 240326 277718 240562 277954
rect 240646 277718 240882 277954
rect 240326 277398 240562 277634
rect 240646 277398 240882 277634
rect 240326 241718 240562 241954
rect 240646 241718 240882 241954
rect 240326 241398 240562 241634
rect 240646 241398 240882 241634
rect 240326 205718 240562 205954
rect 240646 205718 240882 205954
rect 240326 205398 240562 205634
rect 240646 205398 240882 205634
rect 240326 169718 240562 169954
rect 240646 169718 240882 169954
rect 240326 169398 240562 169634
rect 240646 169398 240882 169634
rect 240326 133718 240562 133954
rect 240646 133718 240882 133954
rect 240326 133398 240562 133634
rect 240646 133398 240882 133634
rect 240326 97718 240562 97954
rect 240646 97718 240882 97954
rect 240326 97398 240562 97634
rect 240646 97398 240882 97634
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 240326 -5382 240562 -5146
rect 240646 -5382 240882 -5146
rect 240326 -5702 240562 -5466
rect 240646 -5702 240882 -5466
rect 244826 710362 245062 710598
rect 245146 710362 245382 710598
rect 244826 710042 245062 710278
rect 245146 710042 245382 710278
rect 244826 678218 245062 678454
rect 245146 678218 245382 678454
rect 244826 677898 245062 678134
rect 245146 677898 245382 678134
rect 244826 642218 245062 642454
rect 245146 642218 245382 642454
rect 244826 641898 245062 642134
rect 245146 641898 245382 642134
rect 244826 606218 245062 606454
rect 245146 606218 245382 606454
rect 244826 605898 245062 606134
rect 245146 605898 245382 606134
rect 244826 570218 245062 570454
rect 245146 570218 245382 570454
rect 244826 569898 245062 570134
rect 245146 569898 245382 570134
rect 244826 534218 245062 534454
rect 245146 534218 245382 534454
rect 244826 533898 245062 534134
rect 245146 533898 245382 534134
rect 244826 498218 245062 498454
rect 245146 498218 245382 498454
rect 244826 497898 245062 498134
rect 245146 497898 245382 498134
rect 244826 462218 245062 462454
rect 245146 462218 245382 462454
rect 244826 461898 245062 462134
rect 245146 461898 245382 462134
rect 244826 426218 245062 426454
rect 245146 426218 245382 426454
rect 244826 425898 245062 426134
rect 245146 425898 245382 426134
rect 244826 390218 245062 390454
rect 245146 390218 245382 390454
rect 244826 389898 245062 390134
rect 245146 389898 245382 390134
rect 244826 354218 245062 354454
rect 245146 354218 245382 354454
rect 244826 353898 245062 354134
rect 245146 353898 245382 354134
rect 244826 318218 245062 318454
rect 245146 318218 245382 318454
rect 244826 317898 245062 318134
rect 245146 317898 245382 318134
rect 244826 282218 245062 282454
rect 245146 282218 245382 282454
rect 244826 281898 245062 282134
rect 245146 281898 245382 282134
rect 244826 246218 245062 246454
rect 245146 246218 245382 246454
rect 244826 245898 245062 246134
rect 245146 245898 245382 246134
rect 244826 210218 245062 210454
rect 245146 210218 245382 210454
rect 244826 209898 245062 210134
rect 245146 209898 245382 210134
rect 244826 174218 245062 174454
rect 245146 174218 245382 174454
rect 244826 173898 245062 174134
rect 245146 173898 245382 174134
rect 244826 138218 245062 138454
rect 245146 138218 245382 138454
rect 244826 137898 245062 138134
rect 245146 137898 245382 138134
rect 244826 102218 245062 102454
rect 245146 102218 245382 102454
rect 244826 101898 245062 102134
rect 245146 101898 245382 102134
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 244826 30218 245062 30454
rect 245146 30218 245382 30454
rect 244826 29898 245062 30134
rect 245146 29898 245382 30134
rect 244826 -6342 245062 -6106
rect 245146 -6342 245382 -6106
rect 244826 -6662 245062 -6426
rect 245146 -6662 245382 -6426
rect 249326 711322 249562 711558
rect 249646 711322 249882 711558
rect 249326 711002 249562 711238
rect 249646 711002 249882 711238
rect 249326 682718 249562 682954
rect 249646 682718 249882 682954
rect 249326 682398 249562 682634
rect 249646 682398 249882 682634
rect 249326 646718 249562 646954
rect 249646 646718 249882 646954
rect 249326 646398 249562 646634
rect 249646 646398 249882 646634
rect 249326 610718 249562 610954
rect 249646 610718 249882 610954
rect 249326 610398 249562 610634
rect 249646 610398 249882 610634
rect 249326 574718 249562 574954
rect 249646 574718 249882 574954
rect 249326 574398 249562 574634
rect 249646 574398 249882 574634
rect 249326 538718 249562 538954
rect 249646 538718 249882 538954
rect 249326 538398 249562 538634
rect 249646 538398 249882 538634
rect 249326 502718 249562 502954
rect 249646 502718 249882 502954
rect 249326 502398 249562 502634
rect 249646 502398 249882 502634
rect 249326 466718 249562 466954
rect 249646 466718 249882 466954
rect 249326 466398 249562 466634
rect 249646 466398 249882 466634
rect 249326 430718 249562 430954
rect 249646 430718 249882 430954
rect 249326 430398 249562 430634
rect 249646 430398 249882 430634
rect 249326 394718 249562 394954
rect 249646 394718 249882 394954
rect 249326 394398 249562 394634
rect 249646 394398 249882 394634
rect 249326 358718 249562 358954
rect 249646 358718 249882 358954
rect 249326 358398 249562 358634
rect 249646 358398 249882 358634
rect 249326 322718 249562 322954
rect 249646 322718 249882 322954
rect 249326 322398 249562 322634
rect 249646 322398 249882 322634
rect 249326 286718 249562 286954
rect 249646 286718 249882 286954
rect 249326 286398 249562 286634
rect 249646 286398 249882 286634
rect 249326 250718 249562 250954
rect 249646 250718 249882 250954
rect 249326 250398 249562 250634
rect 249646 250398 249882 250634
rect 249326 214718 249562 214954
rect 249646 214718 249882 214954
rect 249326 214398 249562 214634
rect 249646 214398 249882 214634
rect 249326 178718 249562 178954
rect 249646 178718 249882 178954
rect 249326 178398 249562 178634
rect 249646 178398 249882 178634
rect 249326 142718 249562 142954
rect 249646 142718 249882 142954
rect 249326 142398 249562 142634
rect 249646 142398 249882 142634
rect 249326 106718 249562 106954
rect 249646 106718 249882 106954
rect 249326 106398 249562 106634
rect 249646 106398 249882 106634
rect 249326 70718 249562 70954
rect 249646 70718 249882 70954
rect 249326 70398 249562 70634
rect 249646 70398 249882 70634
rect 249326 34718 249562 34954
rect 249646 34718 249882 34954
rect 249326 34398 249562 34634
rect 249646 34398 249882 34634
rect 249326 -7302 249562 -7066
rect 249646 -7302 249882 -7066
rect 249326 -7622 249562 -7386
rect 249646 -7622 249882 -7386
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 258326 705562 258562 705798
rect 258646 705562 258882 705798
rect 258326 705242 258562 705478
rect 258646 705242 258882 705478
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 258326 655718 258562 655954
rect 258646 655718 258882 655954
rect 258326 655398 258562 655634
rect 258646 655398 258882 655634
rect 258326 619718 258562 619954
rect 258646 619718 258882 619954
rect 258326 619398 258562 619634
rect 258646 619398 258882 619634
rect 258326 583718 258562 583954
rect 258646 583718 258882 583954
rect 258326 583398 258562 583634
rect 258646 583398 258882 583634
rect 258326 547718 258562 547954
rect 258646 547718 258882 547954
rect 258326 547398 258562 547634
rect 258646 547398 258882 547634
rect 258326 511718 258562 511954
rect 258646 511718 258882 511954
rect 258326 511398 258562 511634
rect 258646 511398 258882 511634
rect 258326 475718 258562 475954
rect 258646 475718 258882 475954
rect 258326 475398 258562 475634
rect 258646 475398 258882 475634
rect 258326 439718 258562 439954
rect 258646 439718 258882 439954
rect 258326 439398 258562 439634
rect 258646 439398 258882 439634
rect 258326 403718 258562 403954
rect 258646 403718 258882 403954
rect 258326 403398 258562 403634
rect 258646 403398 258882 403634
rect 258326 367718 258562 367954
rect 258646 367718 258882 367954
rect 258326 367398 258562 367634
rect 258646 367398 258882 367634
rect 258326 331718 258562 331954
rect 258646 331718 258882 331954
rect 258326 331398 258562 331634
rect 258646 331398 258882 331634
rect 258326 295718 258562 295954
rect 258646 295718 258882 295954
rect 258326 295398 258562 295634
rect 258646 295398 258882 295634
rect 258326 259718 258562 259954
rect 258646 259718 258882 259954
rect 258326 259398 258562 259634
rect 258646 259398 258882 259634
rect 258326 223718 258562 223954
rect 258646 223718 258882 223954
rect 258326 223398 258562 223634
rect 258646 223398 258882 223634
rect 258326 187718 258562 187954
rect 258646 187718 258882 187954
rect 258326 187398 258562 187634
rect 258646 187398 258882 187634
rect 258326 151718 258562 151954
rect 258646 151718 258882 151954
rect 258326 151398 258562 151634
rect 258646 151398 258882 151634
rect 258326 115718 258562 115954
rect 258646 115718 258882 115954
rect 258326 115398 258562 115634
rect 258646 115398 258882 115634
rect 258326 79718 258562 79954
rect 258646 79718 258882 79954
rect 258326 79398 258562 79634
rect 258646 79398 258882 79634
rect 258326 43718 258562 43954
rect 258646 43718 258882 43954
rect 258326 43398 258562 43634
rect 258646 43398 258882 43634
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 258326 -1542 258562 -1306
rect 258646 -1542 258882 -1306
rect 258326 -1862 258562 -1626
rect 258646 -1862 258882 -1626
rect 262826 706522 263062 706758
rect 263146 706522 263382 706758
rect 262826 706202 263062 706438
rect 263146 706202 263382 706438
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 262826 660218 263062 660454
rect 263146 660218 263382 660454
rect 262826 659898 263062 660134
rect 263146 659898 263382 660134
rect 262826 624218 263062 624454
rect 263146 624218 263382 624454
rect 262826 623898 263062 624134
rect 263146 623898 263382 624134
rect 262826 588218 263062 588454
rect 263146 588218 263382 588454
rect 262826 587898 263062 588134
rect 263146 587898 263382 588134
rect 262826 552218 263062 552454
rect 263146 552218 263382 552454
rect 262826 551898 263062 552134
rect 263146 551898 263382 552134
rect 262826 516218 263062 516454
rect 263146 516218 263382 516454
rect 262826 515898 263062 516134
rect 263146 515898 263382 516134
rect 262826 480218 263062 480454
rect 263146 480218 263382 480454
rect 262826 479898 263062 480134
rect 263146 479898 263382 480134
rect 262826 444218 263062 444454
rect 263146 444218 263382 444454
rect 262826 443898 263062 444134
rect 263146 443898 263382 444134
rect 262826 408218 263062 408454
rect 263146 408218 263382 408454
rect 262826 407898 263062 408134
rect 263146 407898 263382 408134
rect 262826 372218 263062 372454
rect 263146 372218 263382 372454
rect 262826 371898 263062 372134
rect 263146 371898 263382 372134
rect 262826 336218 263062 336454
rect 263146 336218 263382 336454
rect 262826 335898 263062 336134
rect 263146 335898 263382 336134
rect 262826 300218 263062 300454
rect 263146 300218 263382 300454
rect 262826 299898 263062 300134
rect 263146 299898 263382 300134
rect 262826 264218 263062 264454
rect 263146 264218 263382 264454
rect 262826 263898 263062 264134
rect 263146 263898 263382 264134
rect 262826 228218 263062 228454
rect 263146 228218 263382 228454
rect 262826 227898 263062 228134
rect 263146 227898 263382 228134
rect 262826 192218 263062 192454
rect 263146 192218 263382 192454
rect 262826 191898 263062 192134
rect 263146 191898 263382 192134
rect 262826 156218 263062 156454
rect 263146 156218 263382 156454
rect 262826 155898 263062 156134
rect 263146 155898 263382 156134
rect 262826 120218 263062 120454
rect 263146 120218 263382 120454
rect 262826 119898 263062 120134
rect 263146 119898 263382 120134
rect 262826 84218 263062 84454
rect 263146 84218 263382 84454
rect 262826 83898 263062 84134
rect 263146 83898 263382 84134
rect 262826 48218 263062 48454
rect 263146 48218 263382 48454
rect 262826 47898 263062 48134
rect 263146 47898 263382 48134
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 262826 -2502 263062 -2266
rect 263146 -2502 263382 -2266
rect 262826 -2822 263062 -2586
rect 263146 -2822 263382 -2586
rect 267326 707482 267562 707718
rect 267646 707482 267882 707718
rect 267326 707162 267562 707398
rect 267646 707162 267882 707398
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 267326 664718 267562 664954
rect 267646 664718 267882 664954
rect 267326 664398 267562 664634
rect 267646 664398 267882 664634
rect 267326 628718 267562 628954
rect 267646 628718 267882 628954
rect 267326 628398 267562 628634
rect 267646 628398 267882 628634
rect 267326 592718 267562 592954
rect 267646 592718 267882 592954
rect 267326 592398 267562 592634
rect 267646 592398 267882 592634
rect 267326 556718 267562 556954
rect 267646 556718 267882 556954
rect 267326 556398 267562 556634
rect 267646 556398 267882 556634
rect 267326 520718 267562 520954
rect 267646 520718 267882 520954
rect 267326 520398 267562 520634
rect 267646 520398 267882 520634
rect 267326 484718 267562 484954
rect 267646 484718 267882 484954
rect 267326 484398 267562 484634
rect 267646 484398 267882 484634
rect 267326 448718 267562 448954
rect 267646 448718 267882 448954
rect 267326 448398 267562 448634
rect 267646 448398 267882 448634
rect 267326 412718 267562 412954
rect 267646 412718 267882 412954
rect 267326 412398 267562 412634
rect 267646 412398 267882 412634
rect 267326 376718 267562 376954
rect 267646 376718 267882 376954
rect 267326 376398 267562 376634
rect 267646 376398 267882 376634
rect 267326 340718 267562 340954
rect 267646 340718 267882 340954
rect 267326 340398 267562 340634
rect 267646 340398 267882 340634
rect 267326 304718 267562 304954
rect 267646 304718 267882 304954
rect 267326 304398 267562 304634
rect 267646 304398 267882 304634
rect 267326 268718 267562 268954
rect 267646 268718 267882 268954
rect 267326 268398 267562 268634
rect 267646 268398 267882 268634
rect 267326 232718 267562 232954
rect 267646 232718 267882 232954
rect 267326 232398 267562 232634
rect 267646 232398 267882 232634
rect 267326 196718 267562 196954
rect 267646 196718 267882 196954
rect 267326 196398 267562 196634
rect 267646 196398 267882 196634
rect 267326 160718 267562 160954
rect 267646 160718 267882 160954
rect 267326 160398 267562 160634
rect 267646 160398 267882 160634
rect 267326 124718 267562 124954
rect 267646 124718 267882 124954
rect 267326 124398 267562 124634
rect 267646 124398 267882 124634
rect 267326 88718 267562 88954
rect 267646 88718 267882 88954
rect 267326 88398 267562 88634
rect 267646 88398 267882 88634
rect 267326 52718 267562 52954
rect 267646 52718 267882 52954
rect 267326 52398 267562 52634
rect 267646 52398 267882 52634
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3462 267562 -3226
rect 267646 -3462 267882 -3226
rect 267326 -3782 267562 -3546
rect 267646 -3782 267882 -3546
rect 271826 708442 272062 708678
rect 272146 708442 272382 708678
rect 271826 708122 272062 708358
rect 272146 708122 272382 708358
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4422 272062 -4186
rect 272146 -4422 272382 -4186
rect 271826 -4742 272062 -4506
rect 272146 -4742 272382 -4506
rect 276326 709402 276562 709638
rect 276646 709402 276882 709638
rect 276326 709082 276562 709318
rect 276646 709082 276882 709318
rect 276326 673718 276562 673954
rect 276646 673718 276882 673954
rect 276326 673398 276562 673634
rect 276646 673398 276882 673634
rect 276326 637718 276562 637954
rect 276646 637718 276882 637954
rect 276326 637398 276562 637634
rect 276646 637398 276882 637634
rect 276326 601718 276562 601954
rect 276646 601718 276882 601954
rect 276326 601398 276562 601634
rect 276646 601398 276882 601634
rect 276326 565718 276562 565954
rect 276646 565718 276882 565954
rect 276326 565398 276562 565634
rect 276646 565398 276882 565634
rect 276326 529718 276562 529954
rect 276646 529718 276882 529954
rect 276326 529398 276562 529634
rect 276646 529398 276882 529634
rect 276326 493718 276562 493954
rect 276646 493718 276882 493954
rect 276326 493398 276562 493634
rect 276646 493398 276882 493634
rect 276326 457718 276562 457954
rect 276646 457718 276882 457954
rect 276326 457398 276562 457634
rect 276646 457398 276882 457634
rect 276326 421718 276562 421954
rect 276646 421718 276882 421954
rect 276326 421398 276562 421634
rect 276646 421398 276882 421634
rect 276326 385718 276562 385954
rect 276646 385718 276882 385954
rect 276326 385398 276562 385634
rect 276646 385398 276882 385634
rect 276326 349718 276562 349954
rect 276646 349718 276882 349954
rect 276326 349398 276562 349634
rect 276646 349398 276882 349634
rect 276326 313718 276562 313954
rect 276646 313718 276882 313954
rect 276326 313398 276562 313634
rect 276646 313398 276882 313634
rect 276326 277718 276562 277954
rect 276646 277718 276882 277954
rect 276326 277398 276562 277634
rect 276646 277398 276882 277634
rect 276326 241718 276562 241954
rect 276646 241718 276882 241954
rect 276326 241398 276562 241634
rect 276646 241398 276882 241634
rect 276326 205718 276562 205954
rect 276646 205718 276882 205954
rect 276326 205398 276562 205634
rect 276646 205398 276882 205634
rect 276326 169718 276562 169954
rect 276646 169718 276882 169954
rect 276326 169398 276562 169634
rect 276646 169398 276882 169634
rect 276326 133718 276562 133954
rect 276646 133718 276882 133954
rect 276326 133398 276562 133634
rect 276646 133398 276882 133634
rect 276326 97718 276562 97954
rect 276646 97718 276882 97954
rect 276326 97398 276562 97634
rect 276646 97398 276882 97634
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 276326 -5382 276562 -5146
rect 276646 -5382 276882 -5146
rect 276326 -5702 276562 -5466
rect 276646 -5702 276882 -5466
rect 280826 710362 281062 710598
rect 281146 710362 281382 710598
rect 280826 710042 281062 710278
rect 281146 710042 281382 710278
rect 280826 678218 281062 678454
rect 281146 678218 281382 678454
rect 280826 677898 281062 678134
rect 281146 677898 281382 678134
rect 280826 642218 281062 642454
rect 281146 642218 281382 642454
rect 280826 641898 281062 642134
rect 281146 641898 281382 642134
rect 280826 606218 281062 606454
rect 281146 606218 281382 606454
rect 280826 605898 281062 606134
rect 281146 605898 281382 606134
rect 280826 570218 281062 570454
rect 281146 570218 281382 570454
rect 280826 569898 281062 570134
rect 281146 569898 281382 570134
rect 280826 534218 281062 534454
rect 281146 534218 281382 534454
rect 280826 533898 281062 534134
rect 281146 533898 281382 534134
rect 280826 498218 281062 498454
rect 281146 498218 281382 498454
rect 280826 497898 281062 498134
rect 281146 497898 281382 498134
rect 280826 462218 281062 462454
rect 281146 462218 281382 462454
rect 280826 461898 281062 462134
rect 281146 461898 281382 462134
rect 280826 426218 281062 426454
rect 281146 426218 281382 426454
rect 280826 425898 281062 426134
rect 281146 425898 281382 426134
rect 280826 390218 281062 390454
rect 281146 390218 281382 390454
rect 280826 389898 281062 390134
rect 281146 389898 281382 390134
rect 280826 354218 281062 354454
rect 281146 354218 281382 354454
rect 280826 353898 281062 354134
rect 281146 353898 281382 354134
rect 280826 318218 281062 318454
rect 281146 318218 281382 318454
rect 280826 317898 281062 318134
rect 281146 317898 281382 318134
rect 280826 282218 281062 282454
rect 281146 282218 281382 282454
rect 280826 281898 281062 282134
rect 281146 281898 281382 282134
rect 280826 246218 281062 246454
rect 281146 246218 281382 246454
rect 280826 245898 281062 246134
rect 281146 245898 281382 246134
rect 280826 210218 281062 210454
rect 281146 210218 281382 210454
rect 280826 209898 281062 210134
rect 281146 209898 281382 210134
rect 280826 174218 281062 174454
rect 281146 174218 281382 174454
rect 280826 173898 281062 174134
rect 281146 173898 281382 174134
rect 280826 138218 281062 138454
rect 281146 138218 281382 138454
rect 280826 137898 281062 138134
rect 281146 137898 281382 138134
rect 280826 102218 281062 102454
rect 281146 102218 281382 102454
rect 280826 101898 281062 102134
rect 281146 101898 281382 102134
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 280826 30218 281062 30454
rect 281146 30218 281382 30454
rect 280826 29898 281062 30134
rect 281146 29898 281382 30134
rect 280826 -6342 281062 -6106
rect 281146 -6342 281382 -6106
rect 280826 -6662 281062 -6426
rect 281146 -6662 281382 -6426
rect 285326 711322 285562 711558
rect 285646 711322 285882 711558
rect 285326 711002 285562 711238
rect 285646 711002 285882 711238
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 285326 610718 285562 610954
rect 285646 610718 285882 610954
rect 285326 610398 285562 610634
rect 285646 610398 285882 610634
rect 285326 574718 285562 574954
rect 285646 574718 285882 574954
rect 285326 574398 285562 574634
rect 285646 574398 285882 574634
rect 285326 538718 285562 538954
rect 285646 538718 285882 538954
rect 285326 538398 285562 538634
rect 285646 538398 285882 538634
rect 285326 502718 285562 502954
rect 285646 502718 285882 502954
rect 285326 502398 285562 502634
rect 285646 502398 285882 502634
rect 285326 466718 285562 466954
rect 285646 466718 285882 466954
rect 285326 466398 285562 466634
rect 285646 466398 285882 466634
rect 285326 430718 285562 430954
rect 285646 430718 285882 430954
rect 285326 430398 285562 430634
rect 285646 430398 285882 430634
rect 285326 394718 285562 394954
rect 285646 394718 285882 394954
rect 285326 394398 285562 394634
rect 285646 394398 285882 394634
rect 285326 358718 285562 358954
rect 285646 358718 285882 358954
rect 285326 358398 285562 358634
rect 285646 358398 285882 358634
rect 285326 322718 285562 322954
rect 285646 322718 285882 322954
rect 285326 322398 285562 322634
rect 285646 322398 285882 322634
rect 285326 286718 285562 286954
rect 285646 286718 285882 286954
rect 285326 286398 285562 286634
rect 285646 286398 285882 286634
rect 285326 250718 285562 250954
rect 285646 250718 285882 250954
rect 285326 250398 285562 250634
rect 285646 250398 285882 250634
rect 285326 214718 285562 214954
rect 285646 214718 285882 214954
rect 285326 214398 285562 214634
rect 285646 214398 285882 214634
rect 285326 178718 285562 178954
rect 285646 178718 285882 178954
rect 285326 178398 285562 178634
rect 285646 178398 285882 178634
rect 285326 142718 285562 142954
rect 285646 142718 285882 142954
rect 285326 142398 285562 142634
rect 285646 142398 285882 142634
rect 285326 106718 285562 106954
rect 285646 106718 285882 106954
rect 285326 106398 285562 106634
rect 285646 106398 285882 106634
rect 285326 70718 285562 70954
rect 285646 70718 285882 70954
rect 285326 70398 285562 70634
rect 285646 70398 285882 70634
rect 285326 34718 285562 34954
rect 285646 34718 285882 34954
rect 285326 34398 285562 34634
rect 285646 34398 285882 34634
rect 285326 -7302 285562 -7066
rect 285646 -7302 285882 -7066
rect 285326 -7622 285562 -7386
rect 285646 -7622 285882 -7386
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 294326 705562 294562 705798
rect 294646 705562 294882 705798
rect 294326 705242 294562 705478
rect 294646 705242 294882 705478
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 294326 619718 294562 619954
rect 294646 619718 294882 619954
rect 294326 619398 294562 619634
rect 294646 619398 294882 619634
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 294326 547718 294562 547954
rect 294646 547718 294882 547954
rect 294326 547398 294562 547634
rect 294646 547398 294882 547634
rect 294326 511718 294562 511954
rect 294646 511718 294882 511954
rect 294326 511398 294562 511634
rect 294646 511398 294882 511634
rect 294326 475718 294562 475954
rect 294646 475718 294882 475954
rect 294326 475398 294562 475634
rect 294646 475398 294882 475634
rect 294326 439718 294562 439954
rect 294646 439718 294882 439954
rect 294326 439398 294562 439634
rect 294646 439398 294882 439634
rect 294326 403718 294562 403954
rect 294646 403718 294882 403954
rect 294326 403398 294562 403634
rect 294646 403398 294882 403634
rect 294326 367718 294562 367954
rect 294646 367718 294882 367954
rect 294326 367398 294562 367634
rect 294646 367398 294882 367634
rect 294326 331718 294562 331954
rect 294646 331718 294882 331954
rect 294326 331398 294562 331634
rect 294646 331398 294882 331634
rect 294326 295718 294562 295954
rect 294646 295718 294882 295954
rect 294326 295398 294562 295634
rect 294646 295398 294882 295634
rect 294326 259718 294562 259954
rect 294646 259718 294882 259954
rect 294326 259398 294562 259634
rect 294646 259398 294882 259634
rect 294326 223718 294562 223954
rect 294646 223718 294882 223954
rect 294326 223398 294562 223634
rect 294646 223398 294882 223634
rect 294326 187718 294562 187954
rect 294646 187718 294882 187954
rect 294326 187398 294562 187634
rect 294646 187398 294882 187634
rect 294326 151718 294562 151954
rect 294646 151718 294882 151954
rect 294326 151398 294562 151634
rect 294646 151398 294882 151634
rect 294326 115718 294562 115954
rect 294646 115718 294882 115954
rect 294326 115398 294562 115634
rect 294646 115398 294882 115634
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 294326 43718 294562 43954
rect 294646 43718 294882 43954
rect 294326 43398 294562 43634
rect 294646 43398 294882 43634
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 294326 -1542 294562 -1306
rect 294646 -1542 294882 -1306
rect 294326 -1862 294562 -1626
rect 294646 -1862 294882 -1626
rect 298826 706522 299062 706758
rect 299146 706522 299382 706758
rect 298826 706202 299062 706438
rect 299146 706202 299382 706438
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 298826 660218 299062 660454
rect 299146 660218 299382 660454
rect 298826 659898 299062 660134
rect 299146 659898 299382 660134
rect 298826 624218 299062 624454
rect 299146 624218 299382 624454
rect 298826 623898 299062 624134
rect 299146 623898 299382 624134
rect 298826 588218 299062 588454
rect 299146 588218 299382 588454
rect 298826 587898 299062 588134
rect 299146 587898 299382 588134
rect 298826 552218 299062 552454
rect 299146 552218 299382 552454
rect 298826 551898 299062 552134
rect 299146 551898 299382 552134
rect 298826 516218 299062 516454
rect 299146 516218 299382 516454
rect 298826 515898 299062 516134
rect 299146 515898 299382 516134
rect 298826 480218 299062 480454
rect 299146 480218 299382 480454
rect 298826 479898 299062 480134
rect 299146 479898 299382 480134
rect 298826 444218 299062 444454
rect 299146 444218 299382 444454
rect 298826 443898 299062 444134
rect 299146 443898 299382 444134
rect 298826 408218 299062 408454
rect 299146 408218 299382 408454
rect 298826 407898 299062 408134
rect 299146 407898 299382 408134
rect 298826 372218 299062 372454
rect 299146 372218 299382 372454
rect 298826 371898 299062 372134
rect 299146 371898 299382 372134
rect 298826 336218 299062 336454
rect 299146 336218 299382 336454
rect 298826 335898 299062 336134
rect 299146 335898 299382 336134
rect 298826 300218 299062 300454
rect 299146 300218 299382 300454
rect 298826 299898 299062 300134
rect 299146 299898 299382 300134
rect 298826 264218 299062 264454
rect 299146 264218 299382 264454
rect 298826 263898 299062 264134
rect 299146 263898 299382 264134
rect 298826 228218 299062 228454
rect 299146 228218 299382 228454
rect 298826 227898 299062 228134
rect 299146 227898 299382 228134
rect 298826 192218 299062 192454
rect 299146 192218 299382 192454
rect 298826 191898 299062 192134
rect 299146 191898 299382 192134
rect 298826 156218 299062 156454
rect 299146 156218 299382 156454
rect 298826 155898 299062 156134
rect 299146 155898 299382 156134
rect 298826 120218 299062 120454
rect 299146 120218 299382 120454
rect 298826 119898 299062 120134
rect 299146 119898 299382 120134
rect 298826 84218 299062 84454
rect 299146 84218 299382 84454
rect 298826 83898 299062 84134
rect 299146 83898 299382 84134
rect 298826 48218 299062 48454
rect 299146 48218 299382 48454
rect 298826 47898 299062 48134
rect 299146 47898 299382 48134
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 298826 -2502 299062 -2266
rect 299146 -2502 299382 -2266
rect 298826 -2822 299062 -2586
rect 299146 -2822 299382 -2586
rect 303326 707482 303562 707718
rect 303646 707482 303882 707718
rect 303326 707162 303562 707398
rect 303646 707162 303882 707398
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 303326 664718 303562 664954
rect 303646 664718 303882 664954
rect 303326 664398 303562 664634
rect 303646 664398 303882 664634
rect 303326 628718 303562 628954
rect 303646 628718 303882 628954
rect 303326 628398 303562 628634
rect 303646 628398 303882 628634
rect 303326 592718 303562 592954
rect 303646 592718 303882 592954
rect 303326 592398 303562 592634
rect 303646 592398 303882 592634
rect 303326 556718 303562 556954
rect 303646 556718 303882 556954
rect 303326 556398 303562 556634
rect 303646 556398 303882 556634
rect 303326 520718 303562 520954
rect 303646 520718 303882 520954
rect 303326 520398 303562 520634
rect 303646 520398 303882 520634
rect 303326 484718 303562 484954
rect 303646 484718 303882 484954
rect 303326 484398 303562 484634
rect 303646 484398 303882 484634
rect 303326 448718 303562 448954
rect 303646 448718 303882 448954
rect 303326 448398 303562 448634
rect 303646 448398 303882 448634
rect 303326 412718 303562 412954
rect 303646 412718 303882 412954
rect 303326 412398 303562 412634
rect 303646 412398 303882 412634
rect 303326 376718 303562 376954
rect 303646 376718 303882 376954
rect 303326 376398 303562 376634
rect 303646 376398 303882 376634
rect 303326 340718 303562 340954
rect 303646 340718 303882 340954
rect 303326 340398 303562 340634
rect 303646 340398 303882 340634
rect 303326 304718 303562 304954
rect 303646 304718 303882 304954
rect 303326 304398 303562 304634
rect 303646 304398 303882 304634
rect 303326 268718 303562 268954
rect 303646 268718 303882 268954
rect 303326 268398 303562 268634
rect 303646 268398 303882 268634
rect 303326 232718 303562 232954
rect 303646 232718 303882 232954
rect 303326 232398 303562 232634
rect 303646 232398 303882 232634
rect 303326 196718 303562 196954
rect 303646 196718 303882 196954
rect 303326 196398 303562 196634
rect 303646 196398 303882 196634
rect 303326 160718 303562 160954
rect 303646 160718 303882 160954
rect 303326 160398 303562 160634
rect 303646 160398 303882 160634
rect 303326 124718 303562 124954
rect 303646 124718 303882 124954
rect 303326 124398 303562 124634
rect 303646 124398 303882 124634
rect 303326 88718 303562 88954
rect 303646 88718 303882 88954
rect 303326 88398 303562 88634
rect 303646 88398 303882 88634
rect 303326 52718 303562 52954
rect 303646 52718 303882 52954
rect 303326 52398 303562 52634
rect 303646 52398 303882 52634
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 303326 -3462 303562 -3226
rect 303646 -3462 303882 -3226
rect 303326 -3782 303562 -3546
rect 303646 -3782 303882 -3546
rect 307826 708442 308062 708678
rect 308146 708442 308382 708678
rect 307826 708122 308062 708358
rect 308146 708122 308382 708358
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4422 308062 -4186
rect 308146 -4422 308382 -4186
rect 307826 -4742 308062 -4506
rect 308146 -4742 308382 -4506
rect 312326 709402 312562 709638
rect 312646 709402 312882 709638
rect 312326 709082 312562 709318
rect 312646 709082 312882 709318
rect 312326 673718 312562 673954
rect 312646 673718 312882 673954
rect 312326 673398 312562 673634
rect 312646 673398 312882 673634
rect 312326 637718 312562 637954
rect 312646 637718 312882 637954
rect 312326 637398 312562 637634
rect 312646 637398 312882 637634
rect 312326 601718 312562 601954
rect 312646 601718 312882 601954
rect 312326 601398 312562 601634
rect 312646 601398 312882 601634
rect 312326 565718 312562 565954
rect 312646 565718 312882 565954
rect 312326 565398 312562 565634
rect 312646 565398 312882 565634
rect 312326 529718 312562 529954
rect 312646 529718 312882 529954
rect 312326 529398 312562 529634
rect 312646 529398 312882 529634
rect 312326 493718 312562 493954
rect 312646 493718 312882 493954
rect 312326 493398 312562 493634
rect 312646 493398 312882 493634
rect 312326 457718 312562 457954
rect 312646 457718 312882 457954
rect 312326 457398 312562 457634
rect 312646 457398 312882 457634
rect 312326 421718 312562 421954
rect 312646 421718 312882 421954
rect 312326 421398 312562 421634
rect 312646 421398 312882 421634
rect 312326 385718 312562 385954
rect 312646 385718 312882 385954
rect 312326 385398 312562 385634
rect 312646 385398 312882 385634
rect 312326 349718 312562 349954
rect 312646 349718 312882 349954
rect 312326 349398 312562 349634
rect 312646 349398 312882 349634
rect 312326 313718 312562 313954
rect 312646 313718 312882 313954
rect 312326 313398 312562 313634
rect 312646 313398 312882 313634
rect 312326 277718 312562 277954
rect 312646 277718 312882 277954
rect 312326 277398 312562 277634
rect 312646 277398 312882 277634
rect 312326 241718 312562 241954
rect 312646 241718 312882 241954
rect 312326 241398 312562 241634
rect 312646 241398 312882 241634
rect 312326 205718 312562 205954
rect 312646 205718 312882 205954
rect 312326 205398 312562 205634
rect 312646 205398 312882 205634
rect 312326 169718 312562 169954
rect 312646 169718 312882 169954
rect 312326 169398 312562 169634
rect 312646 169398 312882 169634
rect 312326 133718 312562 133954
rect 312646 133718 312882 133954
rect 312326 133398 312562 133634
rect 312646 133398 312882 133634
rect 312326 97718 312562 97954
rect 312646 97718 312882 97954
rect 312326 97398 312562 97634
rect 312646 97398 312882 97634
rect 312326 61718 312562 61954
rect 312646 61718 312882 61954
rect 312326 61398 312562 61634
rect 312646 61398 312882 61634
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 312326 -5382 312562 -5146
rect 312646 -5382 312882 -5146
rect 312326 -5702 312562 -5466
rect 312646 -5702 312882 -5466
rect 316826 710362 317062 710598
rect 317146 710362 317382 710598
rect 316826 710042 317062 710278
rect 317146 710042 317382 710278
rect 316826 678218 317062 678454
rect 317146 678218 317382 678454
rect 316826 677898 317062 678134
rect 317146 677898 317382 678134
rect 316826 642218 317062 642454
rect 317146 642218 317382 642454
rect 316826 641898 317062 642134
rect 317146 641898 317382 642134
rect 316826 606218 317062 606454
rect 317146 606218 317382 606454
rect 316826 605898 317062 606134
rect 317146 605898 317382 606134
rect 316826 570218 317062 570454
rect 317146 570218 317382 570454
rect 316826 569898 317062 570134
rect 317146 569898 317382 570134
rect 316826 534218 317062 534454
rect 317146 534218 317382 534454
rect 316826 533898 317062 534134
rect 317146 533898 317382 534134
rect 316826 498218 317062 498454
rect 317146 498218 317382 498454
rect 316826 497898 317062 498134
rect 317146 497898 317382 498134
rect 316826 462218 317062 462454
rect 317146 462218 317382 462454
rect 316826 461898 317062 462134
rect 317146 461898 317382 462134
rect 316826 426218 317062 426454
rect 317146 426218 317382 426454
rect 316826 425898 317062 426134
rect 317146 425898 317382 426134
rect 316826 390218 317062 390454
rect 317146 390218 317382 390454
rect 316826 389898 317062 390134
rect 317146 389898 317382 390134
rect 316826 354218 317062 354454
rect 317146 354218 317382 354454
rect 316826 353898 317062 354134
rect 317146 353898 317382 354134
rect 316826 318218 317062 318454
rect 317146 318218 317382 318454
rect 316826 317898 317062 318134
rect 317146 317898 317382 318134
rect 316826 282218 317062 282454
rect 317146 282218 317382 282454
rect 316826 281898 317062 282134
rect 317146 281898 317382 282134
rect 316826 246218 317062 246454
rect 317146 246218 317382 246454
rect 316826 245898 317062 246134
rect 317146 245898 317382 246134
rect 316826 210218 317062 210454
rect 317146 210218 317382 210454
rect 316826 209898 317062 210134
rect 317146 209898 317382 210134
rect 316826 174218 317062 174454
rect 317146 174218 317382 174454
rect 316826 173898 317062 174134
rect 317146 173898 317382 174134
rect 316826 138218 317062 138454
rect 317146 138218 317382 138454
rect 316826 137898 317062 138134
rect 317146 137898 317382 138134
rect 316826 102218 317062 102454
rect 317146 102218 317382 102454
rect 316826 101898 317062 102134
rect 317146 101898 317382 102134
rect 316826 66218 317062 66454
rect 317146 66218 317382 66454
rect 316826 65898 317062 66134
rect 317146 65898 317382 66134
rect 316826 30218 317062 30454
rect 317146 30218 317382 30454
rect 316826 29898 317062 30134
rect 317146 29898 317382 30134
rect 316826 -6342 317062 -6106
rect 317146 -6342 317382 -6106
rect 316826 -6662 317062 -6426
rect 317146 -6662 317382 -6426
rect 321326 711322 321562 711558
rect 321646 711322 321882 711558
rect 321326 711002 321562 711238
rect 321646 711002 321882 711238
rect 321326 682718 321562 682954
rect 321646 682718 321882 682954
rect 321326 682398 321562 682634
rect 321646 682398 321882 682634
rect 321326 646718 321562 646954
rect 321646 646718 321882 646954
rect 321326 646398 321562 646634
rect 321646 646398 321882 646634
rect 321326 610718 321562 610954
rect 321646 610718 321882 610954
rect 321326 610398 321562 610634
rect 321646 610398 321882 610634
rect 321326 574718 321562 574954
rect 321646 574718 321882 574954
rect 321326 574398 321562 574634
rect 321646 574398 321882 574634
rect 321326 538718 321562 538954
rect 321646 538718 321882 538954
rect 321326 538398 321562 538634
rect 321646 538398 321882 538634
rect 321326 502718 321562 502954
rect 321646 502718 321882 502954
rect 321326 502398 321562 502634
rect 321646 502398 321882 502634
rect 321326 466718 321562 466954
rect 321646 466718 321882 466954
rect 321326 466398 321562 466634
rect 321646 466398 321882 466634
rect 321326 430718 321562 430954
rect 321646 430718 321882 430954
rect 321326 430398 321562 430634
rect 321646 430398 321882 430634
rect 321326 394718 321562 394954
rect 321646 394718 321882 394954
rect 321326 394398 321562 394634
rect 321646 394398 321882 394634
rect 321326 358718 321562 358954
rect 321646 358718 321882 358954
rect 321326 358398 321562 358634
rect 321646 358398 321882 358634
rect 321326 322718 321562 322954
rect 321646 322718 321882 322954
rect 321326 322398 321562 322634
rect 321646 322398 321882 322634
rect 321326 286718 321562 286954
rect 321646 286718 321882 286954
rect 321326 286398 321562 286634
rect 321646 286398 321882 286634
rect 321326 250718 321562 250954
rect 321646 250718 321882 250954
rect 321326 250398 321562 250634
rect 321646 250398 321882 250634
rect 321326 214718 321562 214954
rect 321646 214718 321882 214954
rect 321326 214398 321562 214634
rect 321646 214398 321882 214634
rect 321326 178718 321562 178954
rect 321646 178718 321882 178954
rect 321326 178398 321562 178634
rect 321646 178398 321882 178634
rect 321326 142718 321562 142954
rect 321646 142718 321882 142954
rect 321326 142398 321562 142634
rect 321646 142398 321882 142634
rect 321326 106718 321562 106954
rect 321646 106718 321882 106954
rect 321326 106398 321562 106634
rect 321646 106398 321882 106634
rect 321326 70718 321562 70954
rect 321646 70718 321882 70954
rect 321326 70398 321562 70634
rect 321646 70398 321882 70634
rect 321326 34718 321562 34954
rect 321646 34718 321882 34954
rect 321326 34398 321562 34634
rect 321646 34398 321882 34634
rect 321326 -7302 321562 -7066
rect 321646 -7302 321882 -7066
rect 321326 -7622 321562 -7386
rect 321646 -7622 321882 -7386
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 330326 705562 330562 705798
rect 330646 705562 330882 705798
rect 330326 705242 330562 705478
rect 330646 705242 330882 705478
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 330326 655718 330562 655954
rect 330646 655718 330882 655954
rect 330326 655398 330562 655634
rect 330646 655398 330882 655634
rect 330326 619718 330562 619954
rect 330646 619718 330882 619954
rect 330326 619398 330562 619634
rect 330646 619398 330882 619634
rect 330326 583718 330562 583954
rect 330646 583718 330882 583954
rect 330326 583398 330562 583634
rect 330646 583398 330882 583634
rect 330326 547718 330562 547954
rect 330646 547718 330882 547954
rect 330326 547398 330562 547634
rect 330646 547398 330882 547634
rect 330326 511718 330562 511954
rect 330646 511718 330882 511954
rect 330326 511398 330562 511634
rect 330646 511398 330882 511634
rect 330326 475718 330562 475954
rect 330646 475718 330882 475954
rect 330326 475398 330562 475634
rect 330646 475398 330882 475634
rect 330326 439718 330562 439954
rect 330646 439718 330882 439954
rect 330326 439398 330562 439634
rect 330646 439398 330882 439634
rect 330326 403718 330562 403954
rect 330646 403718 330882 403954
rect 330326 403398 330562 403634
rect 330646 403398 330882 403634
rect 330326 367718 330562 367954
rect 330646 367718 330882 367954
rect 330326 367398 330562 367634
rect 330646 367398 330882 367634
rect 330326 331718 330562 331954
rect 330646 331718 330882 331954
rect 330326 331398 330562 331634
rect 330646 331398 330882 331634
rect 330326 295718 330562 295954
rect 330646 295718 330882 295954
rect 330326 295398 330562 295634
rect 330646 295398 330882 295634
rect 330326 259718 330562 259954
rect 330646 259718 330882 259954
rect 330326 259398 330562 259634
rect 330646 259398 330882 259634
rect 330326 223718 330562 223954
rect 330646 223718 330882 223954
rect 330326 223398 330562 223634
rect 330646 223398 330882 223634
rect 330326 187718 330562 187954
rect 330646 187718 330882 187954
rect 330326 187398 330562 187634
rect 330646 187398 330882 187634
rect 330326 151718 330562 151954
rect 330646 151718 330882 151954
rect 330326 151398 330562 151634
rect 330646 151398 330882 151634
rect 330326 115718 330562 115954
rect 330646 115718 330882 115954
rect 330326 115398 330562 115634
rect 330646 115398 330882 115634
rect 330326 79718 330562 79954
rect 330646 79718 330882 79954
rect 330326 79398 330562 79634
rect 330646 79398 330882 79634
rect 330326 43718 330562 43954
rect 330646 43718 330882 43954
rect 330326 43398 330562 43634
rect 330646 43398 330882 43634
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1542 330562 -1306
rect 330646 -1542 330882 -1306
rect 330326 -1862 330562 -1626
rect 330646 -1862 330882 -1626
rect 334826 706522 335062 706758
rect 335146 706522 335382 706758
rect 334826 706202 335062 706438
rect 335146 706202 335382 706438
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 334826 660218 335062 660454
rect 335146 660218 335382 660454
rect 334826 659898 335062 660134
rect 335146 659898 335382 660134
rect 334826 624218 335062 624454
rect 335146 624218 335382 624454
rect 334826 623898 335062 624134
rect 335146 623898 335382 624134
rect 334826 588218 335062 588454
rect 335146 588218 335382 588454
rect 334826 587898 335062 588134
rect 335146 587898 335382 588134
rect 334826 552218 335062 552454
rect 335146 552218 335382 552454
rect 334826 551898 335062 552134
rect 335146 551898 335382 552134
rect 334826 516218 335062 516454
rect 335146 516218 335382 516454
rect 334826 515898 335062 516134
rect 335146 515898 335382 516134
rect 334826 480218 335062 480454
rect 335146 480218 335382 480454
rect 334826 479898 335062 480134
rect 335146 479898 335382 480134
rect 334826 444218 335062 444454
rect 335146 444218 335382 444454
rect 334826 443898 335062 444134
rect 335146 443898 335382 444134
rect 334826 408218 335062 408454
rect 335146 408218 335382 408454
rect 334826 407898 335062 408134
rect 335146 407898 335382 408134
rect 334826 372218 335062 372454
rect 335146 372218 335382 372454
rect 334826 371898 335062 372134
rect 335146 371898 335382 372134
rect 334826 336218 335062 336454
rect 335146 336218 335382 336454
rect 334826 335898 335062 336134
rect 335146 335898 335382 336134
rect 334826 300218 335062 300454
rect 335146 300218 335382 300454
rect 334826 299898 335062 300134
rect 335146 299898 335382 300134
rect 334826 264218 335062 264454
rect 335146 264218 335382 264454
rect 334826 263898 335062 264134
rect 335146 263898 335382 264134
rect 334826 228218 335062 228454
rect 335146 228218 335382 228454
rect 334826 227898 335062 228134
rect 335146 227898 335382 228134
rect 334826 192218 335062 192454
rect 335146 192218 335382 192454
rect 334826 191898 335062 192134
rect 335146 191898 335382 192134
rect 334826 156218 335062 156454
rect 335146 156218 335382 156454
rect 334826 155898 335062 156134
rect 335146 155898 335382 156134
rect 334826 120218 335062 120454
rect 335146 120218 335382 120454
rect 334826 119898 335062 120134
rect 335146 119898 335382 120134
rect 334826 84218 335062 84454
rect 335146 84218 335382 84454
rect 334826 83898 335062 84134
rect 335146 83898 335382 84134
rect 334826 48218 335062 48454
rect 335146 48218 335382 48454
rect 334826 47898 335062 48134
rect 335146 47898 335382 48134
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2502 335062 -2266
rect 335146 -2502 335382 -2266
rect 334826 -2822 335062 -2586
rect 335146 -2822 335382 -2586
rect 339326 707482 339562 707718
rect 339646 707482 339882 707718
rect 339326 707162 339562 707398
rect 339646 707162 339882 707398
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 339326 664718 339562 664954
rect 339646 664718 339882 664954
rect 339326 664398 339562 664634
rect 339646 664398 339882 664634
rect 339326 628718 339562 628954
rect 339646 628718 339882 628954
rect 339326 628398 339562 628634
rect 339646 628398 339882 628634
rect 339326 592718 339562 592954
rect 339646 592718 339882 592954
rect 339326 592398 339562 592634
rect 339646 592398 339882 592634
rect 339326 556718 339562 556954
rect 339646 556718 339882 556954
rect 339326 556398 339562 556634
rect 339646 556398 339882 556634
rect 339326 520718 339562 520954
rect 339646 520718 339882 520954
rect 339326 520398 339562 520634
rect 339646 520398 339882 520634
rect 339326 484718 339562 484954
rect 339646 484718 339882 484954
rect 339326 484398 339562 484634
rect 339646 484398 339882 484634
rect 339326 448718 339562 448954
rect 339646 448718 339882 448954
rect 339326 448398 339562 448634
rect 339646 448398 339882 448634
rect 339326 412718 339562 412954
rect 339646 412718 339882 412954
rect 339326 412398 339562 412634
rect 339646 412398 339882 412634
rect 339326 376718 339562 376954
rect 339646 376718 339882 376954
rect 339326 376398 339562 376634
rect 339646 376398 339882 376634
rect 339326 340718 339562 340954
rect 339646 340718 339882 340954
rect 339326 340398 339562 340634
rect 339646 340398 339882 340634
rect 339326 304718 339562 304954
rect 339646 304718 339882 304954
rect 339326 304398 339562 304634
rect 339646 304398 339882 304634
rect 339326 268718 339562 268954
rect 339646 268718 339882 268954
rect 339326 268398 339562 268634
rect 339646 268398 339882 268634
rect 339326 232718 339562 232954
rect 339646 232718 339882 232954
rect 339326 232398 339562 232634
rect 339646 232398 339882 232634
rect 339326 196718 339562 196954
rect 339646 196718 339882 196954
rect 339326 196398 339562 196634
rect 339646 196398 339882 196634
rect 339326 160718 339562 160954
rect 339646 160718 339882 160954
rect 339326 160398 339562 160634
rect 339646 160398 339882 160634
rect 339326 124718 339562 124954
rect 339646 124718 339882 124954
rect 339326 124398 339562 124634
rect 339646 124398 339882 124634
rect 339326 88718 339562 88954
rect 339646 88718 339882 88954
rect 339326 88398 339562 88634
rect 339646 88398 339882 88634
rect 339326 52718 339562 52954
rect 339646 52718 339882 52954
rect 339326 52398 339562 52634
rect 339646 52398 339882 52634
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 339326 -3462 339562 -3226
rect 339646 -3462 339882 -3226
rect 339326 -3782 339562 -3546
rect 339646 -3782 339882 -3546
rect 343826 708442 344062 708678
rect 344146 708442 344382 708678
rect 343826 708122 344062 708358
rect 344146 708122 344382 708358
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -4422 344062 -4186
rect 344146 -4422 344382 -4186
rect 343826 -4742 344062 -4506
rect 344146 -4742 344382 -4506
rect 348326 709402 348562 709638
rect 348646 709402 348882 709638
rect 348326 709082 348562 709318
rect 348646 709082 348882 709318
rect 348326 673718 348562 673954
rect 348646 673718 348882 673954
rect 348326 673398 348562 673634
rect 348646 673398 348882 673634
rect 348326 637718 348562 637954
rect 348646 637718 348882 637954
rect 348326 637398 348562 637634
rect 348646 637398 348882 637634
rect 348326 601718 348562 601954
rect 348646 601718 348882 601954
rect 348326 601398 348562 601634
rect 348646 601398 348882 601634
rect 348326 565718 348562 565954
rect 348646 565718 348882 565954
rect 348326 565398 348562 565634
rect 348646 565398 348882 565634
rect 348326 529718 348562 529954
rect 348646 529718 348882 529954
rect 348326 529398 348562 529634
rect 348646 529398 348882 529634
rect 348326 493718 348562 493954
rect 348646 493718 348882 493954
rect 348326 493398 348562 493634
rect 348646 493398 348882 493634
rect 348326 457718 348562 457954
rect 348646 457718 348882 457954
rect 348326 457398 348562 457634
rect 348646 457398 348882 457634
rect 348326 421718 348562 421954
rect 348646 421718 348882 421954
rect 348326 421398 348562 421634
rect 348646 421398 348882 421634
rect 348326 385718 348562 385954
rect 348646 385718 348882 385954
rect 348326 385398 348562 385634
rect 348646 385398 348882 385634
rect 348326 349718 348562 349954
rect 348646 349718 348882 349954
rect 348326 349398 348562 349634
rect 348646 349398 348882 349634
rect 348326 313718 348562 313954
rect 348646 313718 348882 313954
rect 348326 313398 348562 313634
rect 348646 313398 348882 313634
rect 348326 277718 348562 277954
rect 348646 277718 348882 277954
rect 348326 277398 348562 277634
rect 348646 277398 348882 277634
rect 348326 241718 348562 241954
rect 348646 241718 348882 241954
rect 348326 241398 348562 241634
rect 348646 241398 348882 241634
rect 348326 205718 348562 205954
rect 348646 205718 348882 205954
rect 348326 205398 348562 205634
rect 348646 205398 348882 205634
rect 348326 169718 348562 169954
rect 348646 169718 348882 169954
rect 348326 169398 348562 169634
rect 348646 169398 348882 169634
rect 348326 133718 348562 133954
rect 348646 133718 348882 133954
rect 348326 133398 348562 133634
rect 348646 133398 348882 133634
rect 348326 97718 348562 97954
rect 348646 97718 348882 97954
rect 348326 97398 348562 97634
rect 348646 97398 348882 97634
rect 348326 61718 348562 61954
rect 348646 61718 348882 61954
rect 348326 61398 348562 61634
rect 348646 61398 348882 61634
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 348326 -5382 348562 -5146
rect 348646 -5382 348882 -5146
rect 348326 -5702 348562 -5466
rect 348646 -5702 348882 -5466
rect 352826 710362 353062 710598
rect 353146 710362 353382 710598
rect 352826 710042 353062 710278
rect 353146 710042 353382 710278
rect 352826 678218 353062 678454
rect 353146 678218 353382 678454
rect 352826 677898 353062 678134
rect 353146 677898 353382 678134
rect 352826 642218 353062 642454
rect 353146 642218 353382 642454
rect 352826 641898 353062 642134
rect 353146 641898 353382 642134
rect 352826 606218 353062 606454
rect 353146 606218 353382 606454
rect 352826 605898 353062 606134
rect 353146 605898 353382 606134
rect 352826 570218 353062 570454
rect 353146 570218 353382 570454
rect 352826 569898 353062 570134
rect 353146 569898 353382 570134
rect 352826 534218 353062 534454
rect 353146 534218 353382 534454
rect 352826 533898 353062 534134
rect 353146 533898 353382 534134
rect 352826 498218 353062 498454
rect 353146 498218 353382 498454
rect 352826 497898 353062 498134
rect 353146 497898 353382 498134
rect 352826 462218 353062 462454
rect 353146 462218 353382 462454
rect 352826 461898 353062 462134
rect 353146 461898 353382 462134
rect 352826 426218 353062 426454
rect 353146 426218 353382 426454
rect 352826 425898 353062 426134
rect 353146 425898 353382 426134
rect 352826 390218 353062 390454
rect 353146 390218 353382 390454
rect 352826 389898 353062 390134
rect 353146 389898 353382 390134
rect 352826 354218 353062 354454
rect 353146 354218 353382 354454
rect 352826 353898 353062 354134
rect 353146 353898 353382 354134
rect 352826 318218 353062 318454
rect 353146 318218 353382 318454
rect 352826 317898 353062 318134
rect 353146 317898 353382 318134
rect 352826 282218 353062 282454
rect 353146 282218 353382 282454
rect 352826 281898 353062 282134
rect 353146 281898 353382 282134
rect 352826 246218 353062 246454
rect 353146 246218 353382 246454
rect 352826 245898 353062 246134
rect 353146 245898 353382 246134
rect 352826 210218 353062 210454
rect 353146 210218 353382 210454
rect 352826 209898 353062 210134
rect 353146 209898 353382 210134
rect 352826 174218 353062 174454
rect 353146 174218 353382 174454
rect 352826 173898 353062 174134
rect 353146 173898 353382 174134
rect 352826 138218 353062 138454
rect 353146 138218 353382 138454
rect 352826 137898 353062 138134
rect 353146 137898 353382 138134
rect 352826 102218 353062 102454
rect 353146 102218 353382 102454
rect 352826 101898 353062 102134
rect 353146 101898 353382 102134
rect 352826 66218 353062 66454
rect 353146 66218 353382 66454
rect 352826 65898 353062 66134
rect 353146 65898 353382 66134
rect 352826 30218 353062 30454
rect 353146 30218 353382 30454
rect 352826 29898 353062 30134
rect 353146 29898 353382 30134
rect 352826 -6342 353062 -6106
rect 353146 -6342 353382 -6106
rect 352826 -6662 353062 -6426
rect 353146 -6662 353382 -6426
rect 357326 711322 357562 711558
rect 357646 711322 357882 711558
rect 357326 711002 357562 711238
rect 357646 711002 357882 711238
rect 357326 682718 357562 682954
rect 357646 682718 357882 682954
rect 357326 682398 357562 682634
rect 357646 682398 357882 682634
rect 357326 646718 357562 646954
rect 357646 646718 357882 646954
rect 357326 646398 357562 646634
rect 357646 646398 357882 646634
rect 357326 610718 357562 610954
rect 357646 610718 357882 610954
rect 357326 610398 357562 610634
rect 357646 610398 357882 610634
rect 357326 574718 357562 574954
rect 357646 574718 357882 574954
rect 357326 574398 357562 574634
rect 357646 574398 357882 574634
rect 357326 538718 357562 538954
rect 357646 538718 357882 538954
rect 357326 538398 357562 538634
rect 357646 538398 357882 538634
rect 357326 502718 357562 502954
rect 357646 502718 357882 502954
rect 357326 502398 357562 502634
rect 357646 502398 357882 502634
rect 357326 466718 357562 466954
rect 357646 466718 357882 466954
rect 357326 466398 357562 466634
rect 357646 466398 357882 466634
rect 357326 430718 357562 430954
rect 357646 430718 357882 430954
rect 357326 430398 357562 430634
rect 357646 430398 357882 430634
rect 357326 394718 357562 394954
rect 357646 394718 357882 394954
rect 357326 394398 357562 394634
rect 357646 394398 357882 394634
rect 357326 358718 357562 358954
rect 357646 358718 357882 358954
rect 357326 358398 357562 358634
rect 357646 358398 357882 358634
rect 357326 322718 357562 322954
rect 357646 322718 357882 322954
rect 357326 322398 357562 322634
rect 357646 322398 357882 322634
rect 357326 286718 357562 286954
rect 357646 286718 357882 286954
rect 357326 286398 357562 286634
rect 357646 286398 357882 286634
rect 357326 250718 357562 250954
rect 357646 250718 357882 250954
rect 357326 250398 357562 250634
rect 357646 250398 357882 250634
rect 357326 214718 357562 214954
rect 357646 214718 357882 214954
rect 357326 214398 357562 214634
rect 357646 214398 357882 214634
rect 357326 178718 357562 178954
rect 357646 178718 357882 178954
rect 357326 178398 357562 178634
rect 357646 178398 357882 178634
rect 357326 142718 357562 142954
rect 357646 142718 357882 142954
rect 357326 142398 357562 142634
rect 357646 142398 357882 142634
rect 357326 106718 357562 106954
rect 357646 106718 357882 106954
rect 357326 106398 357562 106634
rect 357646 106398 357882 106634
rect 357326 70718 357562 70954
rect 357646 70718 357882 70954
rect 357326 70398 357562 70634
rect 357646 70398 357882 70634
rect 357326 34718 357562 34954
rect 357646 34718 357882 34954
rect 357326 34398 357562 34634
rect 357646 34398 357882 34634
rect 357326 -7302 357562 -7066
rect 357646 -7302 357882 -7066
rect 357326 -7622 357562 -7386
rect 357646 -7622 357882 -7386
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 366326 705562 366562 705798
rect 366646 705562 366882 705798
rect 366326 705242 366562 705478
rect 366646 705242 366882 705478
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 366326 655718 366562 655954
rect 366646 655718 366882 655954
rect 366326 655398 366562 655634
rect 366646 655398 366882 655634
rect 366326 619718 366562 619954
rect 366646 619718 366882 619954
rect 366326 619398 366562 619634
rect 366646 619398 366882 619634
rect 366326 583718 366562 583954
rect 366646 583718 366882 583954
rect 366326 583398 366562 583634
rect 366646 583398 366882 583634
rect 366326 547718 366562 547954
rect 366646 547718 366882 547954
rect 366326 547398 366562 547634
rect 366646 547398 366882 547634
rect 366326 511718 366562 511954
rect 366646 511718 366882 511954
rect 366326 511398 366562 511634
rect 366646 511398 366882 511634
rect 366326 475718 366562 475954
rect 366646 475718 366882 475954
rect 366326 475398 366562 475634
rect 366646 475398 366882 475634
rect 366326 439718 366562 439954
rect 366646 439718 366882 439954
rect 366326 439398 366562 439634
rect 366646 439398 366882 439634
rect 366326 403718 366562 403954
rect 366646 403718 366882 403954
rect 366326 403398 366562 403634
rect 366646 403398 366882 403634
rect 366326 367718 366562 367954
rect 366646 367718 366882 367954
rect 366326 367398 366562 367634
rect 366646 367398 366882 367634
rect 366326 331718 366562 331954
rect 366646 331718 366882 331954
rect 366326 331398 366562 331634
rect 366646 331398 366882 331634
rect 366326 295718 366562 295954
rect 366646 295718 366882 295954
rect 366326 295398 366562 295634
rect 366646 295398 366882 295634
rect 366326 259718 366562 259954
rect 366646 259718 366882 259954
rect 366326 259398 366562 259634
rect 366646 259398 366882 259634
rect 366326 223718 366562 223954
rect 366646 223718 366882 223954
rect 366326 223398 366562 223634
rect 366646 223398 366882 223634
rect 366326 187718 366562 187954
rect 366646 187718 366882 187954
rect 366326 187398 366562 187634
rect 366646 187398 366882 187634
rect 366326 151718 366562 151954
rect 366646 151718 366882 151954
rect 366326 151398 366562 151634
rect 366646 151398 366882 151634
rect 366326 115718 366562 115954
rect 366646 115718 366882 115954
rect 366326 115398 366562 115634
rect 366646 115398 366882 115634
rect 366326 79718 366562 79954
rect 366646 79718 366882 79954
rect 366326 79398 366562 79634
rect 366646 79398 366882 79634
rect 366326 43718 366562 43954
rect 366646 43718 366882 43954
rect 366326 43398 366562 43634
rect 366646 43398 366882 43634
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 366326 -1542 366562 -1306
rect 366646 -1542 366882 -1306
rect 366326 -1862 366562 -1626
rect 366646 -1862 366882 -1626
rect 370826 706522 371062 706758
rect 371146 706522 371382 706758
rect 370826 706202 371062 706438
rect 371146 706202 371382 706438
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 370826 660218 371062 660454
rect 371146 660218 371382 660454
rect 370826 659898 371062 660134
rect 371146 659898 371382 660134
rect 370826 624218 371062 624454
rect 371146 624218 371382 624454
rect 370826 623898 371062 624134
rect 371146 623898 371382 624134
rect 370826 588218 371062 588454
rect 371146 588218 371382 588454
rect 370826 587898 371062 588134
rect 371146 587898 371382 588134
rect 370826 552218 371062 552454
rect 371146 552218 371382 552454
rect 370826 551898 371062 552134
rect 371146 551898 371382 552134
rect 370826 516218 371062 516454
rect 371146 516218 371382 516454
rect 370826 515898 371062 516134
rect 371146 515898 371382 516134
rect 370826 480218 371062 480454
rect 371146 480218 371382 480454
rect 370826 479898 371062 480134
rect 371146 479898 371382 480134
rect 370826 444218 371062 444454
rect 371146 444218 371382 444454
rect 370826 443898 371062 444134
rect 371146 443898 371382 444134
rect 370826 408218 371062 408454
rect 371146 408218 371382 408454
rect 370826 407898 371062 408134
rect 371146 407898 371382 408134
rect 370826 372218 371062 372454
rect 371146 372218 371382 372454
rect 370826 371898 371062 372134
rect 371146 371898 371382 372134
rect 370826 336218 371062 336454
rect 371146 336218 371382 336454
rect 370826 335898 371062 336134
rect 371146 335898 371382 336134
rect 370826 300218 371062 300454
rect 371146 300218 371382 300454
rect 370826 299898 371062 300134
rect 371146 299898 371382 300134
rect 370826 264218 371062 264454
rect 371146 264218 371382 264454
rect 370826 263898 371062 264134
rect 371146 263898 371382 264134
rect 370826 228218 371062 228454
rect 371146 228218 371382 228454
rect 370826 227898 371062 228134
rect 371146 227898 371382 228134
rect 370826 192218 371062 192454
rect 371146 192218 371382 192454
rect 370826 191898 371062 192134
rect 371146 191898 371382 192134
rect 370826 156218 371062 156454
rect 371146 156218 371382 156454
rect 370826 155898 371062 156134
rect 371146 155898 371382 156134
rect 370826 120218 371062 120454
rect 371146 120218 371382 120454
rect 370826 119898 371062 120134
rect 371146 119898 371382 120134
rect 370826 84218 371062 84454
rect 371146 84218 371382 84454
rect 370826 83898 371062 84134
rect 371146 83898 371382 84134
rect 370826 48218 371062 48454
rect 371146 48218 371382 48454
rect 370826 47898 371062 48134
rect 371146 47898 371382 48134
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -2502 371062 -2266
rect 371146 -2502 371382 -2266
rect 370826 -2822 371062 -2586
rect 371146 -2822 371382 -2586
rect 375326 707482 375562 707718
rect 375646 707482 375882 707718
rect 375326 707162 375562 707398
rect 375646 707162 375882 707398
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 375326 664718 375562 664954
rect 375646 664718 375882 664954
rect 375326 664398 375562 664634
rect 375646 664398 375882 664634
rect 375326 628718 375562 628954
rect 375646 628718 375882 628954
rect 375326 628398 375562 628634
rect 375646 628398 375882 628634
rect 375326 592718 375562 592954
rect 375646 592718 375882 592954
rect 375326 592398 375562 592634
rect 375646 592398 375882 592634
rect 375326 556718 375562 556954
rect 375646 556718 375882 556954
rect 375326 556398 375562 556634
rect 375646 556398 375882 556634
rect 375326 520718 375562 520954
rect 375646 520718 375882 520954
rect 375326 520398 375562 520634
rect 375646 520398 375882 520634
rect 375326 484718 375562 484954
rect 375646 484718 375882 484954
rect 375326 484398 375562 484634
rect 375646 484398 375882 484634
rect 375326 448718 375562 448954
rect 375646 448718 375882 448954
rect 375326 448398 375562 448634
rect 375646 448398 375882 448634
rect 375326 412718 375562 412954
rect 375646 412718 375882 412954
rect 375326 412398 375562 412634
rect 375646 412398 375882 412634
rect 375326 376718 375562 376954
rect 375646 376718 375882 376954
rect 375326 376398 375562 376634
rect 375646 376398 375882 376634
rect 375326 340718 375562 340954
rect 375646 340718 375882 340954
rect 375326 340398 375562 340634
rect 375646 340398 375882 340634
rect 375326 304718 375562 304954
rect 375646 304718 375882 304954
rect 375326 304398 375562 304634
rect 375646 304398 375882 304634
rect 375326 268718 375562 268954
rect 375646 268718 375882 268954
rect 375326 268398 375562 268634
rect 375646 268398 375882 268634
rect 375326 232718 375562 232954
rect 375646 232718 375882 232954
rect 375326 232398 375562 232634
rect 375646 232398 375882 232634
rect 375326 196718 375562 196954
rect 375646 196718 375882 196954
rect 375326 196398 375562 196634
rect 375646 196398 375882 196634
rect 375326 160718 375562 160954
rect 375646 160718 375882 160954
rect 375326 160398 375562 160634
rect 375646 160398 375882 160634
rect 375326 124718 375562 124954
rect 375646 124718 375882 124954
rect 375326 124398 375562 124634
rect 375646 124398 375882 124634
rect 375326 88718 375562 88954
rect 375646 88718 375882 88954
rect 375326 88398 375562 88634
rect 375646 88398 375882 88634
rect 375326 52718 375562 52954
rect 375646 52718 375882 52954
rect 375326 52398 375562 52634
rect 375646 52398 375882 52634
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3462 375562 -3226
rect 375646 -3462 375882 -3226
rect 375326 -3782 375562 -3546
rect 375646 -3782 375882 -3546
rect 379826 708442 380062 708678
rect 380146 708442 380382 708678
rect 379826 708122 380062 708358
rect 380146 708122 380382 708358
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4422 380062 -4186
rect 380146 -4422 380382 -4186
rect 379826 -4742 380062 -4506
rect 380146 -4742 380382 -4506
rect 384326 709402 384562 709638
rect 384646 709402 384882 709638
rect 384326 709082 384562 709318
rect 384646 709082 384882 709318
rect 384326 673718 384562 673954
rect 384646 673718 384882 673954
rect 384326 673398 384562 673634
rect 384646 673398 384882 673634
rect 384326 637718 384562 637954
rect 384646 637718 384882 637954
rect 384326 637398 384562 637634
rect 384646 637398 384882 637634
rect 384326 601718 384562 601954
rect 384646 601718 384882 601954
rect 384326 601398 384562 601634
rect 384646 601398 384882 601634
rect 384326 565718 384562 565954
rect 384646 565718 384882 565954
rect 384326 565398 384562 565634
rect 384646 565398 384882 565634
rect 384326 529718 384562 529954
rect 384646 529718 384882 529954
rect 384326 529398 384562 529634
rect 384646 529398 384882 529634
rect 384326 493718 384562 493954
rect 384646 493718 384882 493954
rect 384326 493398 384562 493634
rect 384646 493398 384882 493634
rect 384326 457718 384562 457954
rect 384646 457718 384882 457954
rect 384326 457398 384562 457634
rect 384646 457398 384882 457634
rect 384326 421718 384562 421954
rect 384646 421718 384882 421954
rect 384326 421398 384562 421634
rect 384646 421398 384882 421634
rect 384326 385718 384562 385954
rect 384646 385718 384882 385954
rect 384326 385398 384562 385634
rect 384646 385398 384882 385634
rect 384326 349718 384562 349954
rect 384646 349718 384882 349954
rect 384326 349398 384562 349634
rect 384646 349398 384882 349634
rect 384326 313718 384562 313954
rect 384646 313718 384882 313954
rect 384326 313398 384562 313634
rect 384646 313398 384882 313634
rect 384326 277718 384562 277954
rect 384646 277718 384882 277954
rect 384326 277398 384562 277634
rect 384646 277398 384882 277634
rect 384326 241718 384562 241954
rect 384646 241718 384882 241954
rect 384326 241398 384562 241634
rect 384646 241398 384882 241634
rect 384326 205718 384562 205954
rect 384646 205718 384882 205954
rect 384326 205398 384562 205634
rect 384646 205398 384882 205634
rect 384326 169718 384562 169954
rect 384646 169718 384882 169954
rect 384326 169398 384562 169634
rect 384646 169398 384882 169634
rect 384326 133718 384562 133954
rect 384646 133718 384882 133954
rect 384326 133398 384562 133634
rect 384646 133398 384882 133634
rect 384326 97718 384562 97954
rect 384646 97718 384882 97954
rect 384326 97398 384562 97634
rect 384646 97398 384882 97634
rect 384326 61718 384562 61954
rect 384646 61718 384882 61954
rect 384326 61398 384562 61634
rect 384646 61398 384882 61634
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 384326 -5382 384562 -5146
rect 384646 -5382 384882 -5146
rect 384326 -5702 384562 -5466
rect 384646 -5702 384882 -5466
rect 388826 710362 389062 710598
rect 389146 710362 389382 710598
rect 388826 710042 389062 710278
rect 389146 710042 389382 710278
rect 388826 678218 389062 678454
rect 389146 678218 389382 678454
rect 388826 677898 389062 678134
rect 389146 677898 389382 678134
rect 388826 642218 389062 642454
rect 389146 642218 389382 642454
rect 388826 641898 389062 642134
rect 389146 641898 389382 642134
rect 388826 606218 389062 606454
rect 389146 606218 389382 606454
rect 388826 605898 389062 606134
rect 389146 605898 389382 606134
rect 388826 570218 389062 570454
rect 389146 570218 389382 570454
rect 388826 569898 389062 570134
rect 389146 569898 389382 570134
rect 388826 534218 389062 534454
rect 389146 534218 389382 534454
rect 388826 533898 389062 534134
rect 389146 533898 389382 534134
rect 388826 498218 389062 498454
rect 389146 498218 389382 498454
rect 388826 497898 389062 498134
rect 389146 497898 389382 498134
rect 388826 462218 389062 462454
rect 389146 462218 389382 462454
rect 388826 461898 389062 462134
rect 389146 461898 389382 462134
rect 388826 426218 389062 426454
rect 389146 426218 389382 426454
rect 388826 425898 389062 426134
rect 389146 425898 389382 426134
rect 388826 390218 389062 390454
rect 389146 390218 389382 390454
rect 388826 389898 389062 390134
rect 389146 389898 389382 390134
rect 388826 354218 389062 354454
rect 389146 354218 389382 354454
rect 388826 353898 389062 354134
rect 389146 353898 389382 354134
rect 388826 318218 389062 318454
rect 389146 318218 389382 318454
rect 388826 317898 389062 318134
rect 389146 317898 389382 318134
rect 388826 282218 389062 282454
rect 389146 282218 389382 282454
rect 388826 281898 389062 282134
rect 389146 281898 389382 282134
rect 388826 246218 389062 246454
rect 389146 246218 389382 246454
rect 388826 245898 389062 246134
rect 389146 245898 389382 246134
rect 388826 210218 389062 210454
rect 389146 210218 389382 210454
rect 388826 209898 389062 210134
rect 389146 209898 389382 210134
rect 388826 174218 389062 174454
rect 389146 174218 389382 174454
rect 388826 173898 389062 174134
rect 389146 173898 389382 174134
rect 388826 138218 389062 138454
rect 389146 138218 389382 138454
rect 388826 137898 389062 138134
rect 389146 137898 389382 138134
rect 388826 102218 389062 102454
rect 389146 102218 389382 102454
rect 388826 101898 389062 102134
rect 389146 101898 389382 102134
rect 388826 66218 389062 66454
rect 389146 66218 389382 66454
rect 388826 65898 389062 66134
rect 389146 65898 389382 66134
rect 388826 30218 389062 30454
rect 389146 30218 389382 30454
rect 388826 29898 389062 30134
rect 389146 29898 389382 30134
rect 388826 -6342 389062 -6106
rect 389146 -6342 389382 -6106
rect 388826 -6662 389062 -6426
rect 389146 -6662 389382 -6426
rect 393326 711322 393562 711558
rect 393646 711322 393882 711558
rect 393326 711002 393562 711238
rect 393646 711002 393882 711238
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 393326 610718 393562 610954
rect 393646 610718 393882 610954
rect 393326 610398 393562 610634
rect 393646 610398 393882 610634
rect 393326 574718 393562 574954
rect 393646 574718 393882 574954
rect 393326 574398 393562 574634
rect 393646 574398 393882 574634
rect 393326 538718 393562 538954
rect 393646 538718 393882 538954
rect 393326 538398 393562 538634
rect 393646 538398 393882 538634
rect 393326 502718 393562 502954
rect 393646 502718 393882 502954
rect 393326 502398 393562 502634
rect 393646 502398 393882 502634
rect 393326 466718 393562 466954
rect 393646 466718 393882 466954
rect 393326 466398 393562 466634
rect 393646 466398 393882 466634
rect 393326 430718 393562 430954
rect 393646 430718 393882 430954
rect 393326 430398 393562 430634
rect 393646 430398 393882 430634
rect 393326 394718 393562 394954
rect 393646 394718 393882 394954
rect 393326 394398 393562 394634
rect 393646 394398 393882 394634
rect 393326 358718 393562 358954
rect 393646 358718 393882 358954
rect 393326 358398 393562 358634
rect 393646 358398 393882 358634
rect 393326 322718 393562 322954
rect 393646 322718 393882 322954
rect 393326 322398 393562 322634
rect 393646 322398 393882 322634
rect 393326 286718 393562 286954
rect 393646 286718 393882 286954
rect 393326 286398 393562 286634
rect 393646 286398 393882 286634
rect 393326 250718 393562 250954
rect 393646 250718 393882 250954
rect 393326 250398 393562 250634
rect 393646 250398 393882 250634
rect 393326 214718 393562 214954
rect 393646 214718 393882 214954
rect 393326 214398 393562 214634
rect 393646 214398 393882 214634
rect 393326 178718 393562 178954
rect 393646 178718 393882 178954
rect 393326 178398 393562 178634
rect 393646 178398 393882 178634
rect 393326 142718 393562 142954
rect 393646 142718 393882 142954
rect 393326 142398 393562 142634
rect 393646 142398 393882 142634
rect 393326 106718 393562 106954
rect 393646 106718 393882 106954
rect 393326 106398 393562 106634
rect 393646 106398 393882 106634
rect 393326 70718 393562 70954
rect 393646 70718 393882 70954
rect 393326 70398 393562 70634
rect 393646 70398 393882 70634
rect 393326 34718 393562 34954
rect 393646 34718 393882 34954
rect 393326 34398 393562 34634
rect 393646 34398 393882 34634
rect 393326 -7302 393562 -7066
rect 393646 -7302 393882 -7066
rect 393326 -7622 393562 -7386
rect 393646 -7622 393882 -7386
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 402326 705562 402562 705798
rect 402646 705562 402882 705798
rect 402326 705242 402562 705478
rect 402646 705242 402882 705478
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 402326 619718 402562 619954
rect 402646 619718 402882 619954
rect 402326 619398 402562 619634
rect 402646 619398 402882 619634
rect 402326 583718 402562 583954
rect 402646 583718 402882 583954
rect 402326 583398 402562 583634
rect 402646 583398 402882 583634
rect 402326 547718 402562 547954
rect 402646 547718 402882 547954
rect 402326 547398 402562 547634
rect 402646 547398 402882 547634
rect 402326 511718 402562 511954
rect 402646 511718 402882 511954
rect 402326 511398 402562 511634
rect 402646 511398 402882 511634
rect 402326 475718 402562 475954
rect 402646 475718 402882 475954
rect 402326 475398 402562 475634
rect 402646 475398 402882 475634
rect 402326 439718 402562 439954
rect 402646 439718 402882 439954
rect 402326 439398 402562 439634
rect 402646 439398 402882 439634
rect 402326 403718 402562 403954
rect 402646 403718 402882 403954
rect 402326 403398 402562 403634
rect 402646 403398 402882 403634
rect 402326 367718 402562 367954
rect 402646 367718 402882 367954
rect 402326 367398 402562 367634
rect 402646 367398 402882 367634
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 402326 295718 402562 295954
rect 402646 295718 402882 295954
rect 402326 295398 402562 295634
rect 402646 295398 402882 295634
rect 402326 259718 402562 259954
rect 402646 259718 402882 259954
rect 402326 259398 402562 259634
rect 402646 259398 402882 259634
rect 402326 223718 402562 223954
rect 402646 223718 402882 223954
rect 402326 223398 402562 223634
rect 402646 223398 402882 223634
rect 402326 187718 402562 187954
rect 402646 187718 402882 187954
rect 402326 187398 402562 187634
rect 402646 187398 402882 187634
rect 402326 151718 402562 151954
rect 402646 151718 402882 151954
rect 402326 151398 402562 151634
rect 402646 151398 402882 151634
rect 402326 115718 402562 115954
rect 402646 115718 402882 115954
rect 402326 115398 402562 115634
rect 402646 115398 402882 115634
rect 402326 79718 402562 79954
rect 402646 79718 402882 79954
rect 402326 79398 402562 79634
rect 402646 79398 402882 79634
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1542 402562 -1306
rect 402646 -1542 402882 -1306
rect 402326 -1862 402562 -1626
rect 402646 -1862 402882 -1626
rect 406826 706522 407062 706758
rect 407146 706522 407382 706758
rect 406826 706202 407062 706438
rect 407146 706202 407382 706438
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 406826 624218 407062 624454
rect 407146 624218 407382 624454
rect 406826 623898 407062 624134
rect 407146 623898 407382 624134
rect 406826 588218 407062 588454
rect 407146 588218 407382 588454
rect 406826 587898 407062 588134
rect 407146 587898 407382 588134
rect 406826 552218 407062 552454
rect 407146 552218 407382 552454
rect 406826 551898 407062 552134
rect 407146 551898 407382 552134
rect 406826 516218 407062 516454
rect 407146 516218 407382 516454
rect 406826 515898 407062 516134
rect 407146 515898 407382 516134
rect 406826 480218 407062 480454
rect 407146 480218 407382 480454
rect 406826 479898 407062 480134
rect 407146 479898 407382 480134
rect 406826 444218 407062 444454
rect 407146 444218 407382 444454
rect 406826 443898 407062 444134
rect 407146 443898 407382 444134
rect 406826 408218 407062 408454
rect 407146 408218 407382 408454
rect 406826 407898 407062 408134
rect 407146 407898 407382 408134
rect 406826 372218 407062 372454
rect 407146 372218 407382 372454
rect 406826 371898 407062 372134
rect 407146 371898 407382 372134
rect 406826 336218 407062 336454
rect 407146 336218 407382 336454
rect 406826 335898 407062 336134
rect 407146 335898 407382 336134
rect 406826 300218 407062 300454
rect 407146 300218 407382 300454
rect 406826 299898 407062 300134
rect 407146 299898 407382 300134
rect 406826 264218 407062 264454
rect 407146 264218 407382 264454
rect 406826 263898 407062 264134
rect 407146 263898 407382 264134
rect 406826 228218 407062 228454
rect 407146 228218 407382 228454
rect 406826 227898 407062 228134
rect 407146 227898 407382 228134
rect 406826 192218 407062 192454
rect 407146 192218 407382 192454
rect 406826 191898 407062 192134
rect 407146 191898 407382 192134
rect 406826 156218 407062 156454
rect 407146 156218 407382 156454
rect 406826 155898 407062 156134
rect 407146 155898 407382 156134
rect 406826 120218 407062 120454
rect 407146 120218 407382 120454
rect 406826 119898 407062 120134
rect 407146 119898 407382 120134
rect 406826 84218 407062 84454
rect 407146 84218 407382 84454
rect 406826 83898 407062 84134
rect 407146 83898 407382 84134
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2502 407062 -2266
rect 407146 -2502 407382 -2266
rect 406826 -2822 407062 -2586
rect 407146 -2822 407382 -2586
rect 411326 707482 411562 707718
rect 411646 707482 411882 707718
rect 411326 707162 411562 707398
rect 411646 707162 411882 707398
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 411326 664718 411562 664954
rect 411646 664718 411882 664954
rect 411326 664398 411562 664634
rect 411646 664398 411882 664634
rect 411326 628718 411562 628954
rect 411646 628718 411882 628954
rect 411326 628398 411562 628634
rect 411646 628398 411882 628634
rect 411326 592718 411562 592954
rect 411646 592718 411882 592954
rect 411326 592398 411562 592634
rect 411646 592398 411882 592634
rect 411326 556718 411562 556954
rect 411646 556718 411882 556954
rect 411326 556398 411562 556634
rect 411646 556398 411882 556634
rect 411326 520718 411562 520954
rect 411646 520718 411882 520954
rect 411326 520398 411562 520634
rect 411646 520398 411882 520634
rect 411326 484718 411562 484954
rect 411646 484718 411882 484954
rect 411326 484398 411562 484634
rect 411646 484398 411882 484634
rect 411326 448718 411562 448954
rect 411646 448718 411882 448954
rect 411326 448398 411562 448634
rect 411646 448398 411882 448634
rect 411326 412718 411562 412954
rect 411646 412718 411882 412954
rect 411326 412398 411562 412634
rect 411646 412398 411882 412634
rect 411326 376718 411562 376954
rect 411646 376718 411882 376954
rect 411326 376398 411562 376634
rect 411646 376398 411882 376634
rect 411326 340718 411562 340954
rect 411646 340718 411882 340954
rect 411326 340398 411562 340634
rect 411646 340398 411882 340634
rect 411326 304718 411562 304954
rect 411646 304718 411882 304954
rect 411326 304398 411562 304634
rect 411646 304398 411882 304634
rect 411326 268718 411562 268954
rect 411646 268718 411882 268954
rect 411326 268398 411562 268634
rect 411646 268398 411882 268634
rect 411326 232718 411562 232954
rect 411646 232718 411882 232954
rect 411326 232398 411562 232634
rect 411646 232398 411882 232634
rect 411326 196718 411562 196954
rect 411646 196718 411882 196954
rect 411326 196398 411562 196634
rect 411646 196398 411882 196634
rect 411326 160718 411562 160954
rect 411646 160718 411882 160954
rect 411326 160398 411562 160634
rect 411646 160398 411882 160634
rect 411326 124718 411562 124954
rect 411646 124718 411882 124954
rect 411326 124398 411562 124634
rect 411646 124398 411882 124634
rect 411326 88718 411562 88954
rect 411646 88718 411882 88954
rect 411326 88398 411562 88634
rect 411646 88398 411882 88634
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3462 411562 -3226
rect 411646 -3462 411882 -3226
rect 411326 -3782 411562 -3546
rect 411646 -3782 411882 -3546
rect 415826 708442 416062 708678
rect 416146 708442 416382 708678
rect 415826 708122 416062 708358
rect 416146 708122 416382 708358
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4422 416062 -4186
rect 416146 -4422 416382 -4186
rect 415826 -4742 416062 -4506
rect 416146 -4742 416382 -4506
rect 420326 709402 420562 709638
rect 420646 709402 420882 709638
rect 420326 709082 420562 709318
rect 420646 709082 420882 709318
rect 420326 673718 420562 673954
rect 420646 673718 420882 673954
rect 420326 673398 420562 673634
rect 420646 673398 420882 673634
rect 420326 637718 420562 637954
rect 420646 637718 420882 637954
rect 420326 637398 420562 637634
rect 420646 637398 420882 637634
rect 420326 601718 420562 601954
rect 420646 601718 420882 601954
rect 420326 601398 420562 601634
rect 420646 601398 420882 601634
rect 420326 565718 420562 565954
rect 420646 565718 420882 565954
rect 420326 565398 420562 565634
rect 420646 565398 420882 565634
rect 420326 529718 420562 529954
rect 420646 529718 420882 529954
rect 420326 529398 420562 529634
rect 420646 529398 420882 529634
rect 420326 493718 420562 493954
rect 420646 493718 420882 493954
rect 420326 493398 420562 493634
rect 420646 493398 420882 493634
rect 420326 457718 420562 457954
rect 420646 457718 420882 457954
rect 420326 457398 420562 457634
rect 420646 457398 420882 457634
rect 420326 421718 420562 421954
rect 420646 421718 420882 421954
rect 420326 421398 420562 421634
rect 420646 421398 420882 421634
rect 420326 385718 420562 385954
rect 420646 385718 420882 385954
rect 420326 385398 420562 385634
rect 420646 385398 420882 385634
rect 420326 349718 420562 349954
rect 420646 349718 420882 349954
rect 420326 349398 420562 349634
rect 420646 349398 420882 349634
rect 420326 313718 420562 313954
rect 420646 313718 420882 313954
rect 420326 313398 420562 313634
rect 420646 313398 420882 313634
rect 420326 277718 420562 277954
rect 420646 277718 420882 277954
rect 420326 277398 420562 277634
rect 420646 277398 420882 277634
rect 420326 241718 420562 241954
rect 420646 241718 420882 241954
rect 420326 241398 420562 241634
rect 420646 241398 420882 241634
rect 420326 205718 420562 205954
rect 420646 205718 420882 205954
rect 420326 205398 420562 205634
rect 420646 205398 420882 205634
rect 420326 169718 420562 169954
rect 420646 169718 420882 169954
rect 420326 169398 420562 169634
rect 420646 169398 420882 169634
rect 420326 133718 420562 133954
rect 420646 133718 420882 133954
rect 420326 133398 420562 133634
rect 420646 133398 420882 133634
rect 420326 97718 420562 97954
rect 420646 97718 420882 97954
rect 420326 97398 420562 97634
rect 420646 97398 420882 97634
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5382 420562 -5146
rect 420646 -5382 420882 -5146
rect 420326 -5702 420562 -5466
rect 420646 -5702 420882 -5466
rect 424826 710362 425062 710598
rect 425146 710362 425382 710598
rect 424826 710042 425062 710278
rect 425146 710042 425382 710278
rect 424826 678218 425062 678454
rect 425146 678218 425382 678454
rect 424826 677898 425062 678134
rect 425146 677898 425382 678134
rect 424826 642218 425062 642454
rect 425146 642218 425382 642454
rect 424826 641898 425062 642134
rect 425146 641898 425382 642134
rect 424826 606218 425062 606454
rect 425146 606218 425382 606454
rect 424826 605898 425062 606134
rect 425146 605898 425382 606134
rect 424826 570218 425062 570454
rect 425146 570218 425382 570454
rect 424826 569898 425062 570134
rect 425146 569898 425382 570134
rect 424826 534218 425062 534454
rect 425146 534218 425382 534454
rect 424826 533898 425062 534134
rect 425146 533898 425382 534134
rect 424826 498218 425062 498454
rect 425146 498218 425382 498454
rect 424826 497898 425062 498134
rect 425146 497898 425382 498134
rect 424826 462218 425062 462454
rect 425146 462218 425382 462454
rect 424826 461898 425062 462134
rect 425146 461898 425382 462134
rect 424826 426218 425062 426454
rect 425146 426218 425382 426454
rect 424826 425898 425062 426134
rect 425146 425898 425382 426134
rect 424826 390218 425062 390454
rect 425146 390218 425382 390454
rect 424826 389898 425062 390134
rect 425146 389898 425382 390134
rect 424826 354218 425062 354454
rect 425146 354218 425382 354454
rect 424826 353898 425062 354134
rect 425146 353898 425382 354134
rect 424826 318218 425062 318454
rect 425146 318218 425382 318454
rect 424826 317898 425062 318134
rect 425146 317898 425382 318134
rect 424826 282218 425062 282454
rect 425146 282218 425382 282454
rect 424826 281898 425062 282134
rect 425146 281898 425382 282134
rect 424826 246218 425062 246454
rect 425146 246218 425382 246454
rect 424826 245898 425062 246134
rect 425146 245898 425382 246134
rect 424826 210218 425062 210454
rect 425146 210218 425382 210454
rect 424826 209898 425062 210134
rect 425146 209898 425382 210134
rect 424826 174218 425062 174454
rect 425146 174218 425382 174454
rect 424826 173898 425062 174134
rect 425146 173898 425382 174134
rect 424826 138218 425062 138454
rect 425146 138218 425382 138454
rect 424826 137898 425062 138134
rect 425146 137898 425382 138134
rect 424826 102218 425062 102454
rect 425146 102218 425382 102454
rect 424826 101898 425062 102134
rect 425146 101898 425382 102134
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6342 425062 -6106
rect 425146 -6342 425382 -6106
rect 424826 -6662 425062 -6426
rect 425146 -6662 425382 -6426
rect 429326 711322 429562 711558
rect 429646 711322 429882 711558
rect 429326 711002 429562 711238
rect 429646 711002 429882 711238
rect 429326 682718 429562 682954
rect 429646 682718 429882 682954
rect 429326 682398 429562 682634
rect 429646 682398 429882 682634
rect 429326 646718 429562 646954
rect 429646 646718 429882 646954
rect 429326 646398 429562 646634
rect 429646 646398 429882 646634
rect 429326 610718 429562 610954
rect 429646 610718 429882 610954
rect 429326 610398 429562 610634
rect 429646 610398 429882 610634
rect 429326 574718 429562 574954
rect 429646 574718 429882 574954
rect 429326 574398 429562 574634
rect 429646 574398 429882 574634
rect 429326 538718 429562 538954
rect 429646 538718 429882 538954
rect 429326 538398 429562 538634
rect 429646 538398 429882 538634
rect 429326 502718 429562 502954
rect 429646 502718 429882 502954
rect 429326 502398 429562 502634
rect 429646 502398 429882 502634
rect 429326 466718 429562 466954
rect 429646 466718 429882 466954
rect 429326 466398 429562 466634
rect 429646 466398 429882 466634
rect 429326 430718 429562 430954
rect 429646 430718 429882 430954
rect 429326 430398 429562 430634
rect 429646 430398 429882 430634
rect 429326 394718 429562 394954
rect 429646 394718 429882 394954
rect 429326 394398 429562 394634
rect 429646 394398 429882 394634
rect 429326 358718 429562 358954
rect 429646 358718 429882 358954
rect 429326 358398 429562 358634
rect 429646 358398 429882 358634
rect 429326 322718 429562 322954
rect 429646 322718 429882 322954
rect 429326 322398 429562 322634
rect 429646 322398 429882 322634
rect 429326 286718 429562 286954
rect 429646 286718 429882 286954
rect 429326 286398 429562 286634
rect 429646 286398 429882 286634
rect 429326 250718 429562 250954
rect 429646 250718 429882 250954
rect 429326 250398 429562 250634
rect 429646 250398 429882 250634
rect 429326 214718 429562 214954
rect 429646 214718 429882 214954
rect 429326 214398 429562 214634
rect 429646 214398 429882 214634
rect 429326 178718 429562 178954
rect 429646 178718 429882 178954
rect 429326 178398 429562 178634
rect 429646 178398 429882 178634
rect 429326 142718 429562 142954
rect 429646 142718 429882 142954
rect 429326 142398 429562 142634
rect 429646 142398 429882 142634
rect 429326 106718 429562 106954
rect 429646 106718 429882 106954
rect 429326 106398 429562 106634
rect 429646 106398 429882 106634
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7302 429562 -7066
rect 429646 -7302 429882 -7066
rect 429326 -7622 429562 -7386
rect 429646 -7622 429882 -7386
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 438326 705562 438562 705798
rect 438646 705562 438882 705798
rect 438326 705242 438562 705478
rect 438646 705242 438882 705478
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 438326 655718 438562 655954
rect 438646 655718 438882 655954
rect 438326 655398 438562 655634
rect 438646 655398 438882 655634
rect 438326 619718 438562 619954
rect 438646 619718 438882 619954
rect 438326 619398 438562 619634
rect 438646 619398 438882 619634
rect 438326 583718 438562 583954
rect 438646 583718 438882 583954
rect 438326 583398 438562 583634
rect 438646 583398 438882 583634
rect 438326 547718 438562 547954
rect 438646 547718 438882 547954
rect 438326 547398 438562 547634
rect 438646 547398 438882 547634
rect 438326 511718 438562 511954
rect 438646 511718 438882 511954
rect 438326 511398 438562 511634
rect 438646 511398 438882 511634
rect 438326 475718 438562 475954
rect 438646 475718 438882 475954
rect 438326 475398 438562 475634
rect 438646 475398 438882 475634
rect 438326 439718 438562 439954
rect 438646 439718 438882 439954
rect 438326 439398 438562 439634
rect 438646 439398 438882 439634
rect 438326 403718 438562 403954
rect 438646 403718 438882 403954
rect 438326 403398 438562 403634
rect 438646 403398 438882 403634
rect 438326 367718 438562 367954
rect 438646 367718 438882 367954
rect 438326 367398 438562 367634
rect 438646 367398 438882 367634
rect 438326 331718 438562 331954
rect 438646 331718 438882 331954
rect 438326 331398 438562 331634
rect 438646 331398 438882 331634
rect 438326 295718 438562 295954
rect 438646 295718 438882 295954
rect 438326 295398 438562 295634
rect 438646 295398 438882 295634
rect 438326 259718 438562 259954
rect 438646 259718 438882 259954
rect 438326 259398 438562 259634
rect 438646 259398 438882 259634
rect 438326 223718 438562 223954
rect 438646 223718 438882 223954
rect 438326 223398 438562 223634
rect 438646 223398 438882 223634
rect 438326 187718 438562 187954
rect 438646 187718 438882 187954
rect 438326 187398 438562 187634
rect 438646 187398 438882 187634
rect 438326 151718 438562 151954
rect 438646 151718 438882 151954
rect 438326 151398 438562 151634
rect 438646 151398 438882 151634
rect 438326 115718 438562 115954
rect 438646 115718 438882 115954
rect 438326 115398 438562 115634
rect 438646 115398 438882 115634
rect 438326 79718 438562 79954
rect 438646 79718 438882 79954
rect 438326 79398 438562 79634
rect 438646 79398 438882 79634
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1542 438562 -1306
rect 438646 -1542 438882 -1306
rect 438326 -1862 438562 -1626
rect 438646 -1862 438882 -1626
rect 442826 706522 443062 706758
rect 443146 706522 443382 706758
rect 442826 706202 443062 706438
rect 443146 706202 443382 706438
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 442826 660218 443062 660454
rect 443146 660218 443382 660454
rect 442826 659898 443062 660134
rect 443146 659898 443382 660134
rect 442826 624218 443062 624454
rect 443146 624218 443382 624454
rect 442826 623898 443062 624134
rect 443146 623898 443382 624134
rect 442826 588218 443062 588454
rect 443146 588218 443382 588454
rect 442826 587898 443062 588134
rect 443146 587898 443382 588134
rect 442826 552218 443062 552454
rect 443146 552218 443382 552454
rect 442826 551898 443062 552134
rect 443146 551898 443382 552134
rect 442826 516218 443062 516454
rect 443146 516218 443382 516454
rect 442826 515898 443062 516134
rect 443146 515898 443382 516134
rect 442826 480218 443062 480454
rect 443146 480218 443382 480454
rect 442826 479898 443062 480134
rect 443146 479898 443382 480134
rect 442826 444218 443062 444454
rect 443146 444218 443382 444454
rect 442826 443898 443062 444134
rect 443146 443898 443382 444134
rect 442826 408218 443062 408454
rect 443146 408218 443382 408454
rect 442826 407898 443062 408134
rect 443146 407898 443382 408134
rect 442826 372218 443062 372454
rect 443146 372218 443382 372454
rect 442826 371898 443062 372134
rect 443146 371898 443382 372134
rect 442826 336218 443062 336454
rect 443146 336218 443382 336454
rect 442826 335898 443062 336134
rect 443146 335898 443382 336134
rect 442826 300218 443062 300454
rect 443146 300218 443382 300454
rect 442826 299898 443062 300134
rect 443146 299898 443382 300134
rect 442826 264218 443062 264454
rect 443146 264218 443382 264454
rect 442826 263898 443062 264134
rect 443146 263898 443382 264134
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 442826 192218 443062 192454
rect 443146 192218 443382 192454
rect 442826 191898 443062 192134
rect 443146 191898 443382 192134
rect 442826 156218 443062 156454
rect 443146 156218 443382 156454
rect 442826 155898 443062 156134
rect 443146 155898 443382 156134
rect 442826 120218 443062 120454
rect 443146 120218 443382 120454
rect 442826 119898 443062 120134
rect 443146 119898 443382 120134
rect 442826 84218 443062 84454
rect 443146 84218 443382 84454
rect 442826 83898 443062 84134
rect 443146 83898 443382 84134
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2502 443062 -2266
rect 443146 -2502 443382 -2266
rect 442826 -2822 443062 -2586
rect 443146 -2822 443382 -2586
rect 447326 707482 447562 707718
rect 447646 707482 447882 707718
rect 447326 707162 447562 707398
rect 447646 707162 447882 707398
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 447326 664718 447562 664954
rect 447646 664718 447882 664954
rect 447326 664398 447562 664634
rect 447646 664398 447882 664634
rect 447326 628718 447562 628954
rect 447646 628718 447882 628954
rect 447326 628398 447562 628634
rect 447646 628398 447882 628634
rect 447326 592718 447562 592954
rect 447646 592718 447882 592954
rect 447326 592398 447562 592634
rect 447646 592398 447882 592634
rect 447326 556718 447562 556954
rect 447646 556718 447882 556954
rect 447326 556398 447562 556634
rect 447646 556398 447882 556634
rect 447326 520718 447562 520954
rect 447646 520718 447882 520954
rect 447326 520398 447562 520634
rect 447646 520398 447882 520634
rect 447326 484718 447562 484954
rect 447646 484718 447882 484954
rect 447326 484398 447562 484634
rect 447646 484398 447882 484634
rect 447326 448718 447562 448954
rect 447646 448718 447882 448954
rect 447326 448398 447562 448634
rect 447646 448398 447882 448634
rect 447326 412718 447562 412954
rect 447646 412718 447882 412954
rect 447326 412398 447562 412634
rect 447646 412398 447882 412634
rect 447326 376718 447562 376954
rect 447646 376718 447882 376954
rect 447326 376398 447562 376634
rect 447646 376398 447882 376634
rect 447326 340718 447562 340954
rect 447646 340718 447882 340954
rect 447326 340398 447562 340634
rect 447646 340398 447882 340634
rect 447326 304718 447562 304954
rect 447646 304718 447882 304954
rect 447326 304398 447562 304634
rect 447646 304398 447882 304634
rect 447326 268718 447562 268954
rect 447646 268718 447882 268954
rect 447326 268398 447562 268634
rect 447646 268398 447882 268634
rect 447326 232718 447562 232954
rect 447646 232718 447882 232954
rect 447326 232398 447562 232634
rect 447646 232398 447882 232634
rect 447326 196718 447562 196954
rect 447646 196718 447882 196954
rect 447326 196398 447562 196634
rect 447646 196398 447882 196634
rect 447326 160718 447562 160954
rect 447646 160718 447882 160954
rect 447326 160398 447562 160634
rect 447646 160398 447882 160634
rect 447326 124718 447562 124954
rect 447646 124718 447882 124954
rect 447326 124398 447562 124634
rect 447646 124398 447882 124634
rect 447326 88718 447562 88954
rect 447646 88718 447882 88954
rect 447326 88398 447562 88634
rect 447646 88398 447882 88634
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3462 447562 -3226
rect 447646 -3462 447882 -3226
rect 447326 -3782 447562 -3546
rect 447646 -3782 447882 -3546
rect 451826 708442 452062 708678
rect 452146 708442 452382 708678
rect 451826 708122 452062 708358
rect 452146 708122 452382 708358
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4422 452062 -4186
rect 452146 -4422 452382 -4186
rect 451826 -4742 452062 -4506
rect 452146 -4742 452382 -4506
rect 456326 709402 456562 709638
rect 456646 709402 456882 709638
rect 456326 709082 456562 709318
rect 456646 709082 456882 709318
rect 456326 673718 456562 673954
rect 456646 673718 456882 673954
rect 456326 673398 456562 673634
rect 456646 673398 456882 673634
rect 456326 637718 456562 637954
rect 456646 637718 456882 637954
rect 456326 637398 456562 637634
rect 456646 637398 456882 637634
rect 456326 601718 456562 601954
rect 456646 601718 456882 601954
rect 456326 601398 456562 601634
rect 456646 601398 456882 601634
rect 456326 565718 456562 565954
rect 456646 565718 456882 565954
rect 456326 565398 456562 565634
rect 456646 565398 456882 565634
rect 456326 529718 456562 529954
rect 456646 529718 456882 529954
rect 456326 529398 456562 529634
rect 456646 529398 456882 529634
rect 456326 493718 456562 493954
rect 456646 493718 456882 493954
rect 456326 493398 456562 493634
rect 456646 493398 456882 493634
rect 456326 457718 456562 457954
rect 456646 457718 456882 457954
rect 456326 457398 456562 457634
rect 456646 457398 456882 457634
rect 456326 421718 456562 421954
rect 456646 421718 456882 421954
rect 456326 421398 456562 421634
rect 456646 421398 456882 421634
rect 456326 385718 456562 385954
rect 456646 385718 456882 385954
rect 456326 385398 456562 385634
rect 456646 385398 456882 385634
rect 456326 349718 456562 349954
rect 456646 349718 456882 349954
rect 456326 349398 456562 349634
rect 456646 349398 456882 349634
rect 456326 313718 456562 313954
rect 456646 313718 456882 313954
rect 456326 313398 456562 313634
rect 456646 313398 456882 313634
rect 456326 277718 456562 277954
rect 456646 277718 456882 277954
rect 456326 277398 456562 277634
rect 456646 277398 456882 277634
rect 456326 241718 456562 241954
rect 456646 241718 456882 241954
rect 456326 241398 456562 241634
rect 456646 241398 456882 241634
rect 456326 205718 456562 205954
rect 456646 205718 456882 205954
rect 456326 205398 456562 205634
rect 456646 205398 456882 205634
rect 456326 169718 456562 169954
rect 456646 169718 456882 169954
rect 456326 169398 456562 169634
rect 456646 169398 456882 169634
rect 456326 133718 456562 133954
rect 456646 133718 456882 133954
rect 456326 133398 456562 133634
rect 456646 133398 456882 133634
rect 456326 97718 456562 97954
rect 456646 97718 456882 97954
rect 456326 97398 456562 97634
rect 456646 97398 456882 97634
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5382 456562 -5146
rect 456646 -5382 456882 -5146
rect 456326 -5702 456562 -5466
rect 456646 -5702 456882 -5466
rect 460826 710362 461062 710598
rect 461146 710362 461382 710598
rect 460826 710042 461062 710278
rect 461146 710042 461382 710278
rect 460826 678218 461062 678454
rect 461146 678218 461382 678454
rect 460826 677898 461062 678134
rect 461146 677898 461382 678134
rect 460826 642218 461062 642454
rect 461146 642218 461382 642454
rect 460826 641898 461062 642134
rect 461146 641898 461382 642134
rect 460826 606218 461062 606454
rect 461146 606218 461382 606454
rect 460826 605898 461062 606134
rect 461146 605898 461382 606134
rect 460826 570218 461062 570454
rect 461146 570218 461382 570454
rect 460826 569898 461062 570134
rect 461146 569898 461382 570134
rect 460826 534218 461062 534454
rect 461146 534218 461382 534454
rect 460826 533898 461062 534134
rect 461146 533898 461382 534134
rect 460826 498218 461062 498454
rect 461146 498218 461382 498454
rect 460826 497898 461062 498134
rect 461146 497898 461382 498134
rect 460826 462218 461062 462454
rect 461146 462218 461382 462454
rect 460826 461898 461062 462134
rect 461146 461898 461382 462134
rect 460826 426218 461062 426454
rect 461146 426218 461382 426454
rect 460826 425898 461062 426134
rect 461146 425898 461382 426134
rect 460826 390218 461062 390454
rect 461146 390218 461382 390454
rect 460826 389898 461062 390134
rect 461146 389898 461382 390134
rect 460826 354218 461062 354454
rect 461146 354218 461382 354454
rect 460826 353898 461062 354134
rect 461146 353898 461382 354134
rect 460826 318218 461062 318454
rect 461146 318218 461382 318454
rect 460826 317898 461062 318134
rect 461146 317898 461382 318134
rect 460826 282218 461062 282454
rect 461146 282218 461382 282454
rect 460826 281898 461062 282134
rect 461146 281898 461382 282134
rect 460826 246218 461062 246454
rect 461146 246218 461382 246454
rect 460826 245898 461062 246134
rect 461146 245898 461382 246134
rect 460826 210218 461062 210454
rect 461146 210218 461382 210454
rect 460826 209898 461062 210134
rect 461146 209898 461382 210134
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 460826 138218 461062 138454
rect 461146 138218 461382 138454
rect 460826 137898 461062 138134
rect 461146 137898 461382 138134
rect 460826 102218 461062 102454
rect 461146 102218 461382 102454
rect 460826 101898 461062 102134
rect 461146 101898 461382 102134
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6342 461062 -6106
rect 461146 -6342 461382 -6106
rect 460826 -6662 461062 -6426
rect 461146 -6662 461382 -6426
rect 465326 711322 465562 711558
rect 465646 711322 465882 711558
rect 465326 711002 465562 711238
rect 465646 711002 465882 711238
rect 465326 682718 465562 682954
rect 465646 682718 465882 682954
rect 465326 682398 465562 682634
rect 465646 682398 465882 682634
rect 465326 646718 465562 646954
rect 465646 646718 465882 646954
rect 465326 646398 465562 646634
rect 465646 646398 465882 646634
rect 465326 610718 465562 610954
rect 465646 610718 465882 610954
rect 465326 610398 465562 610634
rect 465646 610398 465882 610634
rect 465326 574718 465562 574954
rect 465646 574718 465882 574954
rect 465326 574398 465562 574634
rect 465646 574398 465882 574634
rect 465326 538718 465562 538954
rect 465646 538718 465882 538954
rect 465326 538398 465562 538634
rect 465646 538398 465882 538634
rect 465326 502718 465562 502954
rect 465646 502718 465882 502954
rect 465326 502398 465562 502634
rect 465646 502398 465882 502634
rect 465326 466718 465562 466954
rect 465646 466718 465882 466954
rect 465326 466398 465562 466634
rect 465646 466398 465882 466634
rect 465326 430718 465562 430954
rect 465646 430718 465882 430954
rect 465326 430398 465562 430634
rect 465646 430398 465882 430634
rect 465326 394718 465562 394954
rect 465646 394718 465882 394954
rect 465326 394398 465562 394634
rect 465646 394398 465882 394634
rect 465326 358718 465562 358954
rect 465646 358718 465882 358954
rect 465326 358398 465562 358634
rect 465646 358398 465882 358634
rect 465326 322718 465562 322954
rect 465646 322718 465882 322954
rect 465326 322398 465562 322634
rect 465646 322398 465882 322634
rect 465326 286718 465562 286954
rect 465646 286718 465882 286954
rect 465326 286398 465562 286634
rect 465646 286398 465882 286634
rect 465326 250718 465562 250954
rect 465646 250718 465882 250954
rect 465326 250398 465562 250634
rect 465646 250398 465882 250634
rect 465326 214718 465562 214954
rect 465646 214718 465882 214954
rect 465326 214398 465562 214634
rect 465646 214398 465882 214634
rect 465326 178718 465562 178954
rect 465646 178718 465882 178954
rect 465326 178398 465562 178634
rect 465646 178398 465882 178634
rect 465326 142718 465562 142954
rect 465646 142718 465882 142954
rect 465326 142398 465562 142634
rect 465646 142398 465882 142634
rect 465326 106718 465562 106954
rect 465646 106718 465882 106954
rect 465326 106398 465562 106634
rect 465646 106398 465882 106634
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7302 465562 -7066
rect 465646 -7302 465882 -7066
rect 465326 -7622 465562 -7386
rect 465646 -7622 465882 -7386
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 474326 705562 474562 705798
rect 474646 705562 474882 705798
rect 474326 705242 474562 705478
rect 474646 705242 474882 705478
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 474326 655718 474562 655954
rect 474646 655718 474882 655954
rect 474326 655398 474562 655634
rect 474646 655398 474882 655634
rect 474326 619718 474562 619954
rect 474646 619718 474882 619954
rect 474326 619398 474562 619634
rect 474646 619398 474882 619634
rect 474326 583718 474562 583954
rect 474646 583718 474882 583954
rect 474326 583398 474562 583634
rect 474646 583398 474882 583634
rect 474326 547718 474562 547954
rect 474646 547718 474882 547954
rect 474326 547398 474562 547634
rect 474646 547398 474882 547634
rect 474326 511718 474562 511954
rect 474646 511718 474882 511954
rect 474326 511398 474562 511634
rect 474646 511398 474882 511634
rect 474326 475718 474562 475954
rect 474646 475718 474882 475954
rect 474326 475398 474562 475634
rect 474646 475398 474882 475634
rect 474326 439718 474562 439954
rect 474646 439718 474882 439954
rect 474326 439398 474562 439634
rect 474646 439398 474882 439634
rect 474326 403718 474562 403954
rect 474646 403718 474882 403954
rect 474326 403398 474562 403634
rect 474646 403398 474882 403634
rect 474326 367718 474562 367954
rect 474646 367718 474882 367954
rect 474326 367398 474562 367634
rect 474646 367398 474882 367634
rect 474326 331718 474562 331954
rect 474646 331718 474882 331954
rect 474326 331398 474562 331634
rect 474646 331398 474882 331634
rect 474326 295718 474562 295954
rect 474646 295718 474882 295954
rect 474326 295398 474562 295634
rect 474646 295398 474882 295634
rect 474326 259718 474562 259954
rect 474646 259718 474882 259954
rect 474326 259398 474562 259634
rect 474646 259398 474882 259634
rect 474326 223718 474562 223954
rect 474646 223718 474882 223954
rect 474326 223398 474562 223634
rect 474646 223398 474882 223634
rect 474326 187718 474562 187954
rect 474646 187718 474882 187954
rect 474326 187398 474562 187634
rect 474646 187398 474882 187634
rect 474326 151718 474562 151954
rect 474646 151718 474882 151954
rect 474326 151398 474562 151634
rect 474646 151398 474882 151634
rect 474326 115718 474562 115954
rect 474646 115718 474882 115954
rect 474326 115398 474562 115634
rect 474646 115398 474882 115634
rect 474326 79718 474562 79954
rect 474646 79718 474882 79954
rect 474326 79398 474562 79634
rect 474646 79398 474882 79634
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1542 474562 -1306
rect 474646 -1542 474882 -1306
rect 474326 -1862 474562 -1626
rect 474646 -1862 474882 -1626
rect 478826 706522 479062 706758
rect 479146 706522 479382 706758
rect 478826 706202 479062 706438
rect 479146 706202 479382 706438
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 478826 660218 479062 660454
rect 479146 660218 479382 660454
rect 478826 659898 479062 660134
rect 479146 659898 479382 660134
rect 478826 624218 479062 624454
rect 479146 624218 479382 624454
rect 478826 623898 479062 624134
rect 479146 623898 479382 624134
rect 478826 588218 479062 588454
rect 479146 588218 479382 588454
rect 478826 587898 479062 588134
rect 479146 587898 479382 588134
rect 478826 552218 479062 552454
rect 479146 552218 479382 552454
rect 478826 551898 479062 552134
rect 479146 551898 479382 552134
rect 478826 516218 479062 516454
rect 479146 516218 479382 516454
rect 478826 515898 479062 516134
rect 479146 515898 479382 516134
rect 478826 480218 479062 480454
rect 479146 480218 479382 480454
rect 478826 479898 479062 480134
rect 479146 479898 479382 480134
rect 478826 444218 479062 444454
rect 479146 444218 479382 444454
rect 478826 443898 479062 444134
rect 479146 443898 479382 444134
rect 478826 408218 479062 408454
rect 479146 408218 479382 408454
rect 478826 407898 479062 408134
rect 479146 407898 479382 408134
rect 478826 372218 479062 372454
rect 479146 372218 479382 372454
rect 478826 371898 479062 372134
rect 479146 371898 479382 372134
rect 478826 336218 479062 336454
rect 479146 336218 479382 336454
rect 478826 335898 479062 336134
rect 479146 335898 479382 336134
rect 478826 300218 479062 300454
rect 479146 300218 479382 300454
rect 478826 299898 479062 300134
rect 479146 299898 479382 300134
rect 478826 264218 479062 264454
rect 479146 264218 479382 264454
rect 478826 263898 479062 264134
rect 479146 263898 479382 264134
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 478826 192218 479062 192454
rect 479146 192218 479382 192454
rect 478826 191898 479062 192134
rect 479146 191898 479382 192134
rect 478826 156218 479062 156454
rect 479146 156218 479382 156454
rect 478826 155898 479062 156134
rect 479146 155898 479382 156134
rect 478826 120218 479062 120454
rect 479146 120218 479382 120454
rect 478826 119898 479062 120134
rect 479146 119898 479382 120134
rect 478826 84218 479062 84454
rect 479146 84218 479382 84454
rect 478826 83898 479062 84134
rect 479146 83898 479382 84134
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2502 479062 -2266
rect 479146 -2502 479382 -2266
rect 478826 -2822 479062 -2586
rect 479146 -2822 479382 -2586
rect 483326 707482 483562 707718
rect 483646 707482 483882 707718
rect 483326 707162 483562 707398
rect 483646 707162 483882 707398
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 483326 664718 483562 664954
rect 483646 664718 483882 664954
rect 483326 664398 483562 664634
rect 483646 664398 483882 664634
rect 483326 628718 483562 628954
rect 483646 628718 483882 628954
rect 483326 628398 483562 628634
rect 483646 628398 483882 628634
rect 483326 592718 483562 592954
rect 483646 592718 483882 592954
rect 483326 592398 483562 592634
rect 483646 592398 483882 592634
rect 483326 556718 483562 556954
rect 483646 556718 483882 556954
rect 483326 556398 483562 556634
rect 483646 556398 483882 556634
rect 483326 520718 483562 520954
rect 483646 520718 483882 520954
rect 483326 520398 483562 520634
rect 483646 520398 483882 520634
rect 483326 484718 483562 484954
rect 483646 484718 483882 484954
rect 483326 484398 483562 484634
rect 483646 484398 483882 484634
rect 483326 448718 483562 448954
rect 483646 448718 483882 448954
rect 483326 448398 483562 448634
rect 483646 448398 483882 448634
rect 483326 412718 483562 412954
rect 483646 412718 483882 412954
rect 483326 412398 483562 412634
rect 483646 412398 483882 412634
rect 483326 376718 483562 376954
rect 483646 376718 483882 376954
rect 483326 376398 483562 376634
rect 483646 376398 483882 376634
rect 483326 340718 483562 340954
rect 483646 340718 483882 340954
rect 483326 340398 483562 340634
rect 483646 340398 483882 340634
rect 483326 304718 483562 304954
rect 483646 304718 483882 304954
rect 483326 304398 483562 304634
rect 483646 304398 483882 304634
rect 483326 268718 483562 268954
rect 483646 268718 483882 268954
rect 483326 268398 483562 268634
rect 483646 268398 483882 268634
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 483326 124718 483562 124954
rect 483646 124718 483882 124954
rect 483326 124398 483562 124634
rect 483646 124398 483882 124634
rect 483326 88718 483562 88954
rect 483646 88718 483882 88954
rect 483326 88398 483562 88634
rect 483646 88398 483882 88634
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3462 483562 -3226
rect 483646 -3462 483882 -3226
rect 483326 -3782 483562 -3546
rect 483646 -3782 483882 -3546
rect 487826 708442 488062 708678
rect 488146 708442 488382 708678
rect 487826 708122 488062 708358
rect 488146 708122 488382 708358
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4422 488062 -4186
rect 488146 -4422 488382 -4186
rect 487826 -4742 488062 -4506
rect 488146 -4742 488382 -4506
rect 492326 709402 492562 709638
rect 492646 709402 492882 709638
rect 492326 709082 492562 709318
rect 492646 709082 492882 709318
rect 492326 673718 492562 673954
rect 492646 673718 492882 673954
rect 492326 673398 492562 673634
rect 492646 673398 492882 673634
rect 492326 637718 492562 637954
rect 492646 637718 492882 637954
rect 492326 637398 492562 637634
rect 492646 637398 492882 637634
rect 492326 601718 492562 601954
rect 492646 601718 492882 601954
rect 492326 601398 492562 601634
rect 492646 601398 492882 601634
rect 492326 565718 492562 565954
rect 492646 565718 492882 565954
rect 492326 565398 492562 565634
rect 492646 565398 492882 565634
rect 492326 529718 492562 529954
rect 492646 529718 492882 529954
rect 492326 529398 492562 529634
rect 492646 529398 492882 529634
rect 492326 493718 492562 493954
rect 492646 493718 492882 493954
rect 492326 493398 492562 493634
rect 492646 493398 492882 493634
rect 492326 457718 492562 457954
rect 492646 457718 492882 457954
rect 492326 457398 492562 457634
rect 492646 457398 492882 457634
rect 492326 421718 492562 421954
rect 492646 421718 492882 421954
rect 492326 421398 492562 421634
rect 492646 421398 492882 421634
rect 492326 385718 492562 385954
rect 492646 385718 492882 385954
rect 492326 385398 492562 385634
rect 492646 385398 492882 385634
rect 492326 349718 492562 349954
rect 492646 349718 492882 349954
rect 492326 349398 492562 349634
rect 492646 349398 492882 349634
rect 492326 313718 492562 313954
rect 492646 313718 492882 313954
rect 492326 313398 492562 313634
rect 492646 313398 492882 313634
rect 492326 277718 492562 277954
rect 492646 277718 492882 277954
rect 492326 277398 492562 277634
rect 492646 277398 492882 277634
rect 492326 241718 492562 241954
rect 492646 241718 492882 241954
rect 492326 241398 492562 241634
rect 492646 241398 492882 241634
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 492326 133718 492562 133954
rect 492646 133718 492882 133954
rect 492326 133398 492562 133634
rect 492646 133398 492882 133634
rect 492326 97718 492562 97954
rect 492646 97718 492882 97954
rect 492326 97398 492562 97634
rect 492646 97398 492882 97634
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5382 492562 -5146
rect 492646 -5382 492882 -5146
rect 492326 -5702 492562 -5466
rect 492646 -5702 492882 -5466
rect 496826 710362 497062 710598
rect 497146 710362 497382 710598
rect 496826 710042 497062 710278
rect 497146 710042 497382 710278
rect 496826 678218 497062 678454
rect 497146 678218 497382 678454
rect 496826 677898 497062 678134
rect 497146 677898 497382 678134
rect 496826 642218 497062 642454
rect 497146 642218 497382 642454
rect 496826 641898 497062 642134
rect 497146 641898 497382 642134
rect 496826 606218 497062 606454
rect 497146 606218 497382 606454
rect 496826 605898 497062 606134
rect 497146 605898 497382 606134
rect 496826 570218 497062 570454
rect 497146 570218 497382 570454
rect 496826 569898 497062 570134
rect 497146 569898 497382 570134
rect 496826 534218 497062 534454
rect 497146 534218 497382 534454
rect 496826 533898 497062 534134
rect 497146 533898 497382 534134
rect 496826 498218 497062 498454
rect 497146 498218 497382 498454
rect 496826 497898 497062 498134
rect 497146 497898 497382 498134
rect 496826 462218 497062 462454
rect 497146 462218 497382 462454
rect 496826 461898 497062 462134
rect 497146 461898 497382 462134
rect 496826 426218 497062 426454
rect 497146 426218 497382 426454
rect 496826 425898 497062 426134
rect 497146 425898 497382 426134
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 496826 354218 497062 354454
rect 497146 354218 497382 354454
rect 496826 353898 497062 354134
rect 497146 353898 497382 354134
rect 496826 318218 497062 318454
rect 497146 318218 497382 318454
rect 496826 317898 497062 318134
rect 497146 317898 497382 318134
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 496826 246218 497062 246454
rect 497146 246218 497382 246454
rect 496826 245898 497062 246134
rect 497146 245898 497382 246134
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 496826 138218 497062 138454
rect 497146 138218 497382 138454
rect 496826 137898 497062 138134
rect 497146 137898 497382 138134
rect 496826 102218 497062 102454
rect 497146 102218 497382 102454
rect 496826 101898 497062 102134
rect 497146 101898 497382 102134
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6342 497062 -6106
rect 497146 -6342 497382 -6106
rect 496826 -6662 497062 -6426
rect 497146 -6662 497382 -6426
rect 501326 711322 501562 711558
rect 501646 711322 501882 711558
rect 501326 711002 501562 711238
rect 501646 711002 501882 711238
rect 501326 682718 501562 682954
rect 501646 682718 501882 682954
rect 501326 682398 501562 682634
rect 501646 682398 501882 682634
rect 501326 646718 501562 646954
rect 501646 646718 501882 646954
rect 501326 646398 501562 646634
rect 501646 646398 501882 646634
rect 501326 610718 501562 610954
rect 501646 610718 501882 610954
rect 501326 610398 501562 610634
rect 501646 610398 501882 610634
rect 501326 574718 501562 574954
rect 501646 574718 501882 574954
rect 501326 574398 501562 574634
rect 501646 574398 501882 574634
rect 501326 538718 501562 538954
rect 501646 538718 501882 538954
rect 501326 538398 501562 538634
rect 501646 538398 501882 538634
rect 501326 502718 501562 502954
rect 501646 502718 501882 502954
rect 501326 502398 501562 502634
rect 501646 502398 501882 502634
rect 501326 466718 501562 466954
rect 501646 466718 501882 466954
rect 501326 466398 501562 466634
rect 501646 466398 501882 466634
rect 501326 430718 501562 430954
rect 501646 430718 501882 430954
rect 501326 430398 501562 430634
rect 501646 430398 501882 430634
rect 501326 394718 501562 394954
rect 501646 394718 501882 394954
rect 501326 394398 501562 394634
rect 501646 394398 501882 394634
rect 501326 358718 501562 358954
rect 501646 358718 501882 358954
rect 501326 358398 501562 358634
rect 501646 358398 501882 358634
rect 501326 322718 501562 322954
rect 501646 322718 501882 322954
rect 501326 322398 501562 322634
rect 501646 322398 501882 322634
rect 501326 286718 501562 286954
rect 501646 286718 501882 286954
rect 501326 286398 501562 286634
rect 501646 286398 501882 286634
rect 501326 250718 501562 250954
rect 501646 250718 501882 250954
rect 501326 250398 501562 250634
rect 501646 250398 501882 250634
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 501326 142718 501562 142954
rect 501646 142718 501882 142954
rect 501326 142398 501562 142634
rect 501646 142398 501882 142634
rect 501326 106718 501562 106954
rect 501646 106718 501882 106954
rect 501326 106398 501562 106634
rect 501646 106398 501882 106634
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7302 501562 -7066
rect 501646 -7302 501882 -7066
rect 501326 -7622 501562 -7386
rect 501646 -7622 501882 -7386
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 510326 705562 510562 705798
rect 510646 705562 510882 705798
rect 510326 705242 510562 705478
rect 510646 705242 510882 705478
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 510326 619718 510562 619954
rect 510646 619718 510882 619954
rect 510326 619398 510562 619634
rect 510646 619398 510882 619634
rect 510326 583718 510562 583954
rect 510646 583718 510882 583954
rect 510326 583398 510562 583634
rect 510646 583398 510882 583634
rect 510326 547718 510562 547954
rect 510646 547718 510882 547954
rect 510326 547398 510562 547634
rect 510646 547398 510882 547634
rect 510326 511718 510562 511954
rect 510646 511718 510882 511954
rect 510326 511398 510562 511634
rect 510646 511398 510882 511634
rect 510326 475718 510562 475954
rect 510646 475718 510882 475954
rect 510326 475398 510562 475634
rect 510646 475398 510882 475634
rect 510326 439718 510562 439954
rect 510646 439718 510882 439954
rect 510326 439398 510562 439634
rect 510646 439398 510882 439634
rect 510326 403718 510562 403954
rect 510646 403718 510882 403954
rect 510326 403398 510562 403634
rect 510646 403398 510882 403634
rect 510326 367718 510562 367954
rect 510646 367718 510882 367954
rect 510326 367398 510562 367634
rect 510646 367398 510882 367634
rect 510326 331718 510562 331954
rect 510646 331718 510882 331954
rect 510326 331398 510562 331634
rect 510646 331398 510882 331634
rect 510326 295718 510562 295954
rect 510646 295718 510882 295954
rect 510326 295398 510562 295634
rect 510646 295398 510882 295634
rect 510326 259718 510562 259954
rect 510646 259718 510882 259954
rect 510326 259398 510562 259634
rect 510646 259398 510882 259634
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 510326 151718 510562 151954
rect 510646 151718 510882 151954
rect 510326 151398 510562 151634
rect 510646 151398 510882 151634
rect 510326 115718 510562 115954
rect 510646 115718 510882 115954
rect 510326 115398 510562 115634
rect 510646 115398 510882 115634
rect 510326 79718 510562 79954
rect 510646 79718 510882 79954
rect 510326 79398 510562 79634
rect 510646 79398 510882 79634
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1542 510562 -1306
rect 510646 -1542 510882 -1306
rect 510326 -1862 510562 -1626
rect 510646 -1862 510882 -1626
rect 514826 706522 515062 706758
rect 515146 706522 515382 706758
rect 514826 706202 515062 706438
rect 515146 706202 515382 706438
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 514826 624218 515062 624454
rect 515146 624218 515382 624454
rect 514826 623898 515062 624134
rect 515146 623898 515382 624134
rect 514826 588218 515062 588454
rect 515146 588218 515382 588454
rect 514826 587898 515062 588134
rect 515146 587898 515382 588134
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 514826 516218 515062 516454
rect 515146 516218 515382 516454
rect 514826 515898 515062 516134
rect 515146 515898 515382 516134
rect 514826 480218 515062 480454
rect 515146 480218 515382 480454
rect 514826 479898 515062 480134
rect 515146 479898 515382 480134
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 514826 408218 515062 408454
rect 515146 408218 515382 408454
rect 514826 407898 515062 408134
rect 515146 407898 515382 408134
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 514826 264218 515062 264454
rect 515146 264218 515382 264454
rect 514826 263898 515062 264134
rect 515146 263898 515382 264134
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2502 515062 -2266
rect 515146 -2502 515382 -2266
rect 514826 -2822 515062 -2586
rect 515146 -2822 515382 -2586
rect 519326 707482 519562 707718
rect 519646 707482 519882 707718
rect 519326 707162 519562 707398
rect 519646 707162 519882 707398
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 519326 628718 519562 628954
rect 519646 628718 519882 628954
rect 519326 628398 519562 628634
rect 519646 628398 519882 628634
rect 519326 592718 519562 592954
rect 519646 592718 519882 592954
rect 519326 592398 519562 592634
rect 519646 592398 519882 592634
rect 519326 556718 519562 556954
rect 519646 556718 519882 556954
rect 519326 556398 519562 556634
rect 519646 556398 519882 556634
rect 519326 520718 519562 520954
rect 519646 520718 519882 520954
rect 519326 520398 519562 520634
rect 519646 520398 519882 520634
rect 519326 484718 519562 484954
rect 519646 484718 519882 484954
rect 519326 484398 519562 484634
rect 519646 484398 519882 484634
rect 519326 448718 519562 448954
rect 519646 448718 519882 448954
rect 519326 448398 519562 448634
rect 519646 448398 519882 448634
rect 519326 412718 519562 412954
rect 519646 412718 519882 412954
rect 519326 412398 519562 412634
rect 519646 412398 519882 412634
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 519326 268718 519562 268954
rect 519646 268718 519882 268954
rect 519326 268398 519562 268634
rect 519646 268398 519882 268634
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 519326 124718 519562 124954
rect 519646 124718 519882 124954
rect 519326 124398 519562 124634
rect 519646 124398 519882 124634
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3462 519562 -3226
rect 519646 -3462 519882 -3226
rect 519326 -3782 519562 -3546
rect 519646 -3782 519882 -3546
rect 523826 708442 524062 708678
rect 524146 708442 524382 708678
rect 523826 708122 524062 708358
rect 524146 708122 524382 708358
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4422 524062 -4186
rect 524146 -4422 524382 -4186
rect 523826 -4742 524062 -4506
rect 524146 -4742 524382 -4506
rect 528326 709402 528562 709638
rect 528646 709402 528882 709638
rect 528326 709082 528562 709318
rect 528646 709082 528882 709318
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 528326 565718 528562 565954
rect 528646 565718 528882 565954
rect 528326 565398 528562 565634
rect 528646 565398 528882 565634
rect 528326 529718 528562 529954
rect 528646 529718 528882 529954
rect 528326 529398 528562 529634
rect 528646 529398 528882 529634
rect 528326 493718 528562 493954
rect 528646 493718 528882 493954
rect 528326 493398 528562 493634
rect 528646 493398 528882 493634
rect 528326 457718 528562 457954
rect 528646 457718 528882 457954
rect 528326 457398 528562 457634
rect 528646 457398 528882 457634
rect 528326 421718 528562 421954
rect 528646 421718 528882 421954
rect 528326 421398 528562 421634
rect 528646 421398 528882 421634
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 528326 277718 528562 277954
rect 528646 277718 528882 277954
rect 528326 277398 528562 277634
rect 528646 277398 528882 277634
rect 528326 241718 528562 241954
rect 528646 241718 528882 241954
rect 528326 241398 528562 241634
rect 528646 241398 528882 241634
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 528326 133718 528562 133954
rect 528646 133718 528882 133954
rect 528326 133398 528562 133634
rect 528646 133398 528882 133634
rect 528326 97718 528562 97954
rect 528646 97718 528882 97954
rect 528326 97398 528562 97634
rect 528646 97398 528882 97634
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5382 528562 -5146
rect 528646 -5382 528882 -5146
rect 528326 -5702 528562 -5466
rect 528646 -5702 528882 -5466
rect 532826 710362 533062 710598
rect 533146 710362 533382 710598
rect 532826 710042 533062 710278
rect 533146 710042 533382 710278
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 532826 570218 533062 570454
rect 533146 570218 533382 570454
rect 532826 569898 533062 570134
rect 533146 569898 533382 570134
rect 532826 534218 533062 534454
rect 533146 534218 533382 534454
rect 532826 533898 533062 534134
rect 533146 533898 533382 534134
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 532826 462218 533062 462454
rect 533146 462218 533382 462454
rect 532826 461898 533062 462134
rect 533146 461898 533382 462134
rect 532826 426218 533062 426454
rect 533146 426218 533382 426454
rect 532826 425898 533062 426134
rect 533146 425898 533382 426134
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 532826 246218 533062 246454
rect 533146 246218 533382 246454
rect 532826 245898 533062 246134
rect 533146 245898 533382 246134
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 532826 138218 533062 138454
rect 533146 138218 533382 138454
rect 532826 137898 533062 138134
rect 533146 137898 533382 138134
rect 532826 102218 533062 102454
rect 533146 102218 533382 102454
rect 532826 101898 533062 102134
rect 533146 101898 533382 102134
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6342 533062 -6106
rect 533146 -6342 533382 -6106
rect 532826 -6662 533062 -6426
rect 533146 -6662 533382 -6426
rect 537326 711322 537562 711558
rect 537646 711322 537882 711558
rect 537326 711002 537562 711238
rect 537646 711002 537882 711238
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 537326 250718 537562 250954
rect 537646 250718 537882 250954
rect 537326 250398 537562 250634
rect 537646 250398 537882 250634
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 537326 142718 537562 142954
rect 537646 142718 537882 142954
rect 537326 142398 537562 142634
rect 537646 142398 537882 142634
rect 537326 106718 537562 106954
rect 537646 106718 537882 106954
rect 537326 106398 537562 106634
rect 537646 106398 537882 106634
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7302 537562 -7066
rect 537646 -7302 537882 -7066
rect 537326 -7622 537562 -7386
rect 537646 -7622 537882 -7386
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 546326 705562 546562 705798
rect 546646 705562 546882 705798
rect 546326 705242 546562 705478
rect 546646 705242 546882 705478
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 546326 259718 546562 259954
rect 546646 259718 546882 259954
rect 546326 259398 546562 259634
rect 546646 259398 546882 259634
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1542 546562 -1306
rect 546646 -1542 546882 -1306
rect 546326 -1862 546562 -1626
rect 546646 -1862 546882 -1626
rect 550826 706522 551062 706758
rect 551146 706522 551382 706758
rect 550826 706202 551062 706438
rect 551146 706202 551382 706438
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 550826 300218 551062 300454
rect 551146 300218 551382 300454
rect 550826 299898 551062 300134
rect 551146 299898 551382 300134
rect 550826 264218 551062 264454
rect 551146 264218 551382 264454
rect 550826 263898 551062 264134
rect 551146 263898 551382 264134
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2502 551062 -2266
rect 551146 -2502 551382 -2266
rect 550826 -2822 551062 -2586
rect 551146 -2822 551382 -2586
rect 555326 707482 555562 707718
rect 555646 707482 555882 707718
rect 555326 707162 555562 707398
rect 555646 707162 555882 707398
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3462 555562 -3226
rect 555646 -3462 555882 -3226
rect 555326 -3782 555562 -3546
rect 555646 -3782 555882 -3546
rect 559826 708442 560062 708678
rect 560146 708442 560382 708678
rect 559826 708122 560062 708358
rect 560146 708122 560382 708358
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4422 560062 -4186
rect 560146 -4422 560382 -4186
rect 559826 -4742 560062 -4506
rect 560146 -4742 560382 -4506
rect 564326 709402 564562 709638
rect 564646 709402 564882 709638
rect 564326 709082 564562 709318
rect 564646 709082 564882 709318
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5382 564562 -5146
rect 564646 -5382 564882 -5146
rect 564326 -5702 564562 -5466
rect 564646 -5702 564882 -5466
rect 568826 710362 569062 710598
rect 569146 710362 569382 710598
rect 568826 710042 569062 710278
rect 569146 710042 569382 710278
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6342 569062 -6106
rect 569146 -6342 569382 -6106
rect 568826 -6662 569062 -6426
rect 569146 -6662 569382 -6426
rect 573326 711322 573562 711558
rect 573646 711322 573882 711558
rect 573326 711002 573562 711238
rect 573646 711002 573882 711238
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7302 573562 -7066
rect 573646 -7302 573882 -7066
rect 573326 -7622 573562 -7386
rect 573646 -7622 573882 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 691718 586538 691954
rect 586622 691718 586858 691954
rect 586302 691398 586538 691634
rect 586622 691398 586858 691634
rect 586302 655718 586538 655954
rect 586622 655718 586858 655954
rect 586302 655398 586538 655634
rect 586622 655398 586858 655634
rect 586302 619718 586538 619954
rect 586622 619718 586858 619954
rect 586302 619398 586538 619634
rect 586622 619398 586858 619634
rect 586302 583718 586538 583954
rect 586622 583718 586858 583954
rect 586302 583398 586538 583634
rect 586622 583398 586858 583634
rect 586302 547718 586538 547954
rect 586622 547718 586858 547954
rect 586302 547398 586538 547634
rect 586622 547398 586858 547634
rect 586302 511718 586538 511954
rect 586622 511718 586858 511954
rect 586302 511398 586538 511634
rect 586622 511398 586858 511634
rect 586302 475718 586538 475954
rect 586622 475718 586858 475954
rect 586302 475398 586538 475634
rect 586622 475398 586858 475634
rect 586302 439718 586538 439954
rect 586622 439718 586858 439954
rect 586302 439398 586538 439634
rect 586622 439398 586858 439634
rect 586302 403718 586538 403954
rect 586622 403718 586858 403954
rect 586302 403398 586538 403634
rect 586622 403398 586858 403634
rect 586302 367718 586538 367954
rect 586622 367718 586858 367954
rect 586302 367398 586538 367634
rect 586622 367398 586858 367634
rect 586302 331718 586538 331954
rect 586622 331718 586858 331954
rect 586302 331398 586538 331634
rect 586622 331398 586858 331634
rect 586302 295718 586538 295954
rect 586622 295718 586858 295954
rect 586302 295398 586538 295634
rect 586622 295398 586858 295634
rect 586302 259718 586538 259954
rect 586622 259718 586858 259954
rect 586302 259398 586538 259634
rect 586622 259398 586858 259634
rect 586302 223718 586538 223954
rect 586622 223718 586858 223954
rect 586302 223398 586538 223634
rect 586622 223398 586858 223634
rect 586302 187718 586538 187954
rect 586622 187718 586858 187954
rect 586302 187398 586538 187634
rect 586622 187398 586858 187634
rect 586302 151718 586538 151954
rect 586622 151718 586858 151954
rect 586302 151398 586538 151634
rect 586622 151398 586858 151634
rect 586302 115718 586538 115954
rect 586622 115718 586858 115954
rect 586302 115398 586538 115634
rect 586622 115398 586858 115634
rect 586302 79718 586538 79954
rect 586622 79718 586858 79954
rect 586302 79398 586538 79634
rect 586622 79398 586858 79634
rect 586302 43718 586538 43954
rect 586622 43718 586858 43954
rect 586302 43398 586538 43634
rect 586622 43398 586858 43634
rect 586302 7718 586538 7954
rect 586622 7718 586858 7954
rect 586302 7398 586538 7634
rect 586622 7398 586858 7634
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 696218 587498 696454
rect 587582 696218 587818 696454
rect 587262 695898 587498 696134
rect 587582 695898 587818 696134
rect 587262 660218 587498 660454
rect 587582 660218 587818 660454
rect 587262 659898 587498 660134
rect 587582 659898 587818 660134
rect 587262 624218 587498 624454
rect 587582 624218 587818 624454
rect 587262 623898 587498 624134
rect 587582 623898 587818 624134
rect 587262 588218 587498 588454
rect 587582 588218 587818 588454
rect 587262 587898 587498 588134
rect 587582 587898 587818 588134
rect 587262 552218 587498 552454
rect 587582 552218 587818 552454
rect 587262 551898 587498 552134
rect 587582 551898 587818 552134
rect 587262 516218 587498 516454
rect 587582 516218 587818 516454
rect 587262 515898 587498 516134
rect 587582 515898 587818 516134
rect 587262 480218 587498 480454
rect 587582 480218 587818 480454
rect 587262 479898 587498 480134
rect 587582 479898 587818 480134
rect 587262 444218 587498 444454
rect 587582 444218 587818 444454
rect 587262 443898 587498 444134
rect 587582 443898 587818 444134
rect 587262 408218 587498 408454
rect 587582 408218 587818 408454
rect 587262 407898 587498 408134
rect 587582 407898 587818 408134
rect 587262 372218 587498 372454
rect 587582 372218 587818 372454
rect 587262 371898 587498 372134
rect 587582 371898 587818 372134
rect 587262 336218 587498 336454
rect 587582 336218 587818 336454
rect 587262 335898 587498 336134
rect 587582 335898 587818 336134
rect 587262 300218 587498 300454
rect 587582 300218 587818 300454
rect 587262 299898 587498 300134
rect 587582 299898 587818 300134
rect 587262 264218 587498 264454
rect 587582 264218 587818 264454
rect 587262 263898 587498 264134
rect 587582 263898 587818 264134
rect 587262 228218 587498 228454
rect 587582 228218 587818 228454
rect 587262 227898 587498 228134
rect 587582 227898 587818 228134
rect 587262 192218 587498 192454
rect 587582 192218 587818 192454
rect 587262 191898 587498 192134
rect 587582 191898 587818 192134
rect 587262 156218 587498 156454
rect 587582 156218 587818 156454
rect 587262 155898 587498 156134
rect 587582 155898 587818 156134
rect 587262 120218 587498 120454
rect 587582 120218 587818 120454
rect 587262 119898 587498 120134
rect 587582 119898 587818 120134
rect 587262 84218 587498 84454
rect 587582 84218 587818 84454
rect 587262 83898 587498 84134
rect 587582 83898 587818 84134
rect 587262 48218 587498 48454
rect 587582 48218 587818 48454
rect 587262 47898 587498 48134
rect 587582 47898 587818 48134
rect 587262 12218 587498 12454
rect 587582 12218 587818 12454
rect 587262 11898 587498 12134
rect 587582 11898 587818 12134
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 700718 588458 700954
rect 588542 700718 588778 700954
rect 588222 700398 588458 700634
rect 588542 700398 588778 700634
rect 588222 664718 588458 664954
rect 588542 664718 588778 664954
rect 588222 664398 588458 664634
rect 588542 664398 588778 664634
rect 588222 628718 588458 628954
rect 588542 628718 588778 628954
rect 588222 628398 588458 628634
rect 588542 628398 588778 628634
rect 588222 592718 588458 592954
rect 588542 592718 588778 592954
rect 588222 592398 588458 592634
rect 588542 592398 588778 592634
rect 588222 556718 588458 556954
rect 588542 556718 588778 556954
rect 588222 556398 588458 556634
rect 588542 556398 588778 556634
rect 588222 520718 588458 520954
rect 588542 520718 588778 520954
rect 588222 520398 588458 520634
rect 588542 520398 588778 520634
rect 588222 484718 588458 484954
rect 588542 484718 588778 484954
rect 588222 484398 588458 484634
rect 588542 484398 588778 484634
rect 588222 448718 588458 448954
rect 588542 448718 588778 448954
rect 588222 448398 588458 448634
rect 588542 448398 588778 448634
rect 588222 412718 588458 412954
rect 588542 412718 588778 412954
rect 588222 412398 588458 412634
rect 588542 412398 588778 412634
rect 588222 376718 588458 376954
rect 588542 376718 588778 376954
rect 588222 376398 588458 376634
rect 588542 376398 588778 376634
rect 588222 340718 588458 340954
rect 588542 340718 588778 340954
rect 588222 340398 588458 340634
rect 588542 340398 588778 340634
rect 588222 304718 588458 304954
rect 588542 304718 588778 304954
rect 588222 304398 588458 304634
rect 588542 304398 588778 304634
rect 588222 268718 588458 268954
rect 588542 268718 588778 268954
rect 588222 268398 588458 268634
rect 588542 268398 588778 268634
rect 588222 232718 588458 232954
rect 588542 232718 588778 232954
rect 588222 232398 588458 232634
rect 588542 232398 588778 232634
rect 588222 196718 588458 196954
rect 588542 196718 588778 196954
rect 588222 196398 588458 196634
rect 588542 196398 588778 196634
rect 588222 160718 588458 160954
rect 588542 160718 588778 160954
rect 588222 160398 588458 160634
rect 588542 160398 588778 160634
rect 588222 124718 588458 124954
rect 588542 124718 588778 124954
rect 588222 124398 588458 124634
rect 588542 124398 588778 124634
rect 588222 88718 588458 88954
rect 588542 88718 588778 88954
rect 588222 88398 588458 88634
rect 588542 88398 588778 88634
rect 588222 52718 588458 52954
rect 588542 52718 588778 52954
rect 588222 52398 588458 52634
rect 588542 52398 588778 52634
rect 588222 16718 588458 16954
rect 588542 16718 588778 16954
rect 588222 16398 588458 16634
rect 588542 16398 588778 16634
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 669218 589418 669454
rect 589502 669218 589738 669454
rect 589182 668898 589418 669134
rect 589502 668898 589738 669134
rect 589182 633218 589418 633454
rect 589502 633218 589738 633454
rect 589182 632898 589418 633134
rect 589502 632898 589738 633134
rect 589182 597218 589418 597454
rect 589502 597218 589738 597454
rect 589182 596898 589418 597134
rect 589502 596898 589738 597134
rect 589182 561218 589418 561454
rect 589502 561218 589738 561454
rect 589182 560898 589418 561134
rect 589502 560898 589738 561134
rect 589182 525218 589418 525454
rect 589502 525218 589738 525454
rect 589182 524898 589418 525134
rect 589502 524898 589738 525134
rect 589182 489218 589418 489454
rect 589502 489218 589738 489454
rect 589182 488898 589418 489134
rect 589502 488898 589738 489134
rect 589182 453218 589418 453454
rect 589502 453218 589738 453454
rect 589182 452898 589418 453134
rect 589502 452898 589738 453134
rect 589182 417218 589418 417454
rect 589502 417218 589738 417454
rect 589182 416898 589418 417134
rect 589502 416898 589738 417134
rect 589182 381218 589418 381454
rect 589502 381218 589738 381454
rect 589182 380898 589418 381134
rect 589502 380898 589738 381134
rect 589182 345218 589418 345454
rect 589502 345218 589738 345454
rect 589182 344898 589418 345134
rect 589502 344898 589738 345134
rect 589182 309218 589418 309454
rect 589502 309218 589738 309454
rect 589182 308898 589418 309134
rect 589502 308898 589738 309134
rect 589182 273218 589418 273454
rect 589502 273218 589738 273454
rect 589182 272898 589418 273134
rect 589502 272898 589738 273134
rect 589182 237218 589418 237454
rect 589502 237218 589738 237454
rect 589182 236898 589418 237134
rect 589502 236898 589738 237134
rect 589182 201218 589418 201454
rect 589502 201218 589738 201454
rect 589182 200898 589418 201134
rect 589502 200898 589738 201134
rect 589182 165218 589418 165454
rect 589502 165218 589738 165454
rect 589182 164898 589418 165134
rect 589502 164898 589738 165134
rect 589182 129218 589418 129454
rect 589502 129218 589738 129454
rect 589182 128898 589418 129134
rect 589502 128898 589738 129134
rect 589182 93218 589418 93454
rect 589502 93218 589738 93454
rect 589182 92898 589418 93134
rect 589502 92898 589738 93134
rect 589182 57218 589418 57454
rect 589502 57218 589738 57454
rect 589182 56898 589418 57134
rect 589502 56898 589738 57134
rect 589182 21218 589418 21454
rect 589502 21218 589738 21454
rect 589182 20898 589418 21134
rect 589502 20898 589738 21134
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 673718 590378 673954
rect 590462 673718 590698 673954
rect 590142 673398 590378 673634
rect 590462 673398 590698 673634
rect 590142 637718 590378 637954
rect 590462 637718 590698 637954
rect 590142 637398 590378 637634
rect 590462 637398 590698 637634
rect 590142 601718 590378 601954
rect 590462 601718 590698 601954
rect 590142 601398 590378 601634
rect 590462 601398 590698 601634
rect 590142 565718 590378 565954
rect 590462 565718 590698 565954
rect 590142 565398 590378 565634
rect 590462 565398 590698 565634
rect 590142 529718 590378 529954
rect 590462 529718 590698 529954
rect 590142 529398 590378 529634
rect 590462 529398 590698 529634
rect 590142 493718 590378 493954
rect 590462 493718 590698 493954
rect 590142 493398 590378 493634
rect 590462 493398 590698 493634
rect 590142 457718 590378 457954
rect 590462 457718 590698 457954
rect 590142 457398 590378 457634
rect 590462 457398 590698 457634
rect 590142 421718 590378 421954
rect 590462 421718 590698 421954
rect 590142 421398 590378 421634
rect 590462 421398 590698 421634
rect 590142 385718 590378 385954
rect 590462 385718 590698 385954
rect 590142 385398 590378 385634
rect 590462 385398 590698 385634
rect 590142 349718 590378 349954
rect 590462 349718 590698 349954
rect 590142 349398 590378 349634
rect 590462 349398 590698 349634
rect 590142 313718 590378 313954
rect 590462 313718 590698 313954
rect 590142 313398 590378 313634
rect 590462 313398 590698 313634
rect 590142 277718 590378 277954
rect 590462 277718 590698 277954
rect 590142 277398 590378 277634
rect 590462 277398 590698 277634
rect 590142 241718 590378 241954
rect 590462 241718 590698 241954
rect 590142 241398 590378 241634
rect 590462 241398 590698 241634
rect 590142 205718 590378 205954
rect 590462 205718 590698 205954
rect 590142 205398 590378 205634
rect 590462 205398 590698 205634
rect 590142 169718 590378 169954
rect 590462 169718 590698 169954
rect 590142 169398 590378 169634
rect 590462 169398 590698 169634
rect 590142 133718 590378 133954
rect 590462 133718 590698 133954
rect 590142 133398 590378 133634
rect 590462 133398 590698 133634
rect 590142 97718 590378 97954
rect 590462 97718 590698 97954
rect 590142 97398 590378 97634
rect 590462 97398 590698 97634
rect 590142 61718 590378 61954
rect 590462 61718 590698 61954
rect 590142 61398 590378 61634
rect 590462 61398 590698 61634
rect 590142 25718 590378 25954
rect 590462 25718 590698 25954
rect 590142 25398 590378 25634
rect 590462 25398 590698 25634
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 678218 591338 678454
rect 591422 678218 591658 678454
rect 591102 677898 591338 678134
rect 591422 677898 591658 678134
rect 591102 642218 591338 642454
rect 591422 642218 591658 642454
rect 591102 641898 591338 642134
rect 591422 641898 591658 642134
rect 591102 606218 591338 606454
rect 591422 606218 591658 606454
rect 591102 605898 591338 606134
rect 591422 605898 591658 606134
rect 591102 570218 591338 570454
rect 591422 570218 591658 570454
rect 591102 569898 591338 570134
rect 591422 569898 591658 570134
rect 591102 534218 591338 534454
rect 591422 534218 591658 534454
rect 591102 533898 591338 534134
rect 591422 533898 591658 534134
rect 591102 498218 591338 498454
rect 591422 498218 591658 498454
rect 591102 497898 591338 498134
rect 591422 497898 591658 498134
rect 591102 462218 591338 462454
rect 591422 462218 591658 462454
rect 591102 461898 591338 462134
rect 591422 461898 591658 462134
rect 591102 426218 591338 426454
rect 591422 426218 591658 426454
rect 591102 425898 591338 426134
rect 591422 425898 591658 426134
rect 591102 390218 591338 390454
rect 591422 390218 591658 390454
rect 591102 389898 591338 390134
rect 591422 389898 591658 390134
rect 591102 354218 591338 354454
rect 591422 354218 591658 354454
rect 591102 353898 591338 354134
rect 591422 353898 591658 354134
rect 591102 318218 591338 318454
rect 591422 318218 591658 318454
rect 591102 317898 591338 318134
rect 591422 317898 591658 318134
rect 591102 282218 591338 282454
rect 591422 282218 591658 282454
rect 591102 281898 591338 282134
rect 591422 281898 591658 282134
rect 591102 246218 591338 246454
rect 591422 246218 591658 246454
rect 591102 245898 591338 246134
rect 591422 245898 591658 246134
rect 591102 210218 591338 210454
rect 591422 210218 591658 210454
rect 591102 209898 591338 210134
rect 591422 209898 591658 210134
rect 591102 174218 591338 174454
rect 591422 174218 591658 174454
rect 591102 173898 591338 174134
rect 591422 173898 591658 174134
rect 591102 138218 591338 138454
rect 591422 138218 591658 138454
rect 591102 137898 591338 138134
rect 591422 137898 591658 138134
rect 591102 102218 591338 102454
rect 591422 102218 591658 102454
rect 591102 101898 591338 102134
rect 591422 101898 591658 102134
rect 591102 66218 591338 66454
rect 591422 66218 591658 66454
rect 591102 65898 591338 66134
rect 591422 65898 591658 66134
rect 591102 30218 591338 30454
rect 591422 30218 591658 30454
rect 591102 29898 591338 30134
rect 591422 29898 591658 30134
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 682718 592298 682954
rect 592382 682718 592618 682954
rect 592062 682398 592298 682634
rect 592382 682398 592618 682634
rect 592062 646718 592298 646954
rect 592382 646718 592618 646954
rect 592062 646398 592298 646634
rect 592382 646398 592618 646634
rect 592062 610718 592298 610954
rect 592382 610718 592618 610954
rect 592062 610398 592298 610634
rect 592382 610398 592618 610634
rect 592062 574718 592298 574954
rect 592382 574718 592618 574954
rect 592062 574398 592298 574634
rect 592382 574398 592618 574634
rect 592062 538718 592298 538954
rect 592382 538718 592618 538954
rect 592062 538398 592298 538634
rect 592382 538398 592618 538634
rect 592062 502718 592298 502954
rect 592382 502718 592618 502954
rect 592062 502398 592298 502634
rect 592382 502398 592618 502634
rect 592062 466718 592298 466954
rect 592382 466718 592618 466954
rect 592062 466398 592298 466634
rect 592382 466398 592618 466634
rect 592062 430718 592298 430954
rect 592382 430718 592618 430954
rect 592062 430398 592298 430634
rect 592382 430398 592618 430634
rect 592062 394718 592298 394954
rect 592382 394718 592618 394954
rect 592062 394398 592298 394634
rect 592382 394398 592618 394634
rect 592062 358718 592298 358954
rect 592382 358718 592618 358954
rect 592062 358398 592298 358634
rect 592382 358398 592618 358634
rect 592062 322718 592298 322954
rect 592382 322718 592618 322954
rect 592062 322398 592298 322634
rect 592382 322398 592618 322634
rect 592062 286718 592298 286954
rect 592382 286718 592618 286954
rect 592062 286398 592298 286634
rect 592382 286398 592618 286634
rect 592062 250718 592298 250954
rect 592382 250718 592618 250954
rect 592062 250398 592298 250634
rect 592382 250398 592618 250634
rect 592062 214718 592298 214954
rect 592382 214718 592618 214954
rect 592062 214398 592298 214634
rect 592382 214398 592618 214634
rect 592062 178718 592298 178954
rect 592382 178718 592618 178954
rect 592062 178398 592298 178634
rect 592382 178398 592618 178634
rect 592062 142718 592298 142954
rect 592382 142718 592618 142954
rect 592062 142398 592298 142634
rect 592382 142398 592618 142634
rect 592062 106718 592298 106954
rect 592382 106718 592618 106954
rect 592062 106398 592298 106634
rect 592382 106398 592618 106634
rect 592062 70718 592298 70954
rect 592382 70718 592618 70954
rect 592062 70398 592298 70634
rect 592382 70398 592618 70634
rect 592062 34718 592298 34954
rect 592382 34718 592618 34954
rect 592062 34398 592298 34634
rect 592382 34398 592618 34634
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700954 592650 700986
rect -8726 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 592650 700954
rect -8726 700634 592650 700718
rect -8726 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 592650 700634
rect -8726 700366 592650 700398
rect -8726 696454 592650 696486
rect -8726 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 691954 592650 691986
rect -8726 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 592650 691954
rect -8726 691634 592650 691718
rect -8726 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 592650 691634
rect -8726 691366 592650 691398
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 682954 592650 682986
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect -8726 682634 592650 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect -8726 682366 592650 682398
rect -8726 678454 592650 678486
rect -8726 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 592650 678454
rect -8726 678134 592650 678218
rect -8726 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 592650 678134
rect -8726 677866 592650 677898
rect -8726 673954 592650 673986
rect -8726 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 592650 673954
rect -8726 673634 592650 673718
rect -8726 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 592650 673634
rect -8726 673366 592650 673398
rect -8726 669454 592650 669486
rect -8726 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 592650 669454
rect -8726 669134 592650 669218
rect -8726 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 592650 669134
rect -8726 668866 592650 668898
rect -8726 664954 592650 664986
rect -8726 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 592650 664954
rect -8726 664634 592650 664718
rect -8726 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 592650 664634
rect -8726 664366 592650 664398
rect -8726 660454 592650 660486
rect -8726 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 655954 592650 655986
rect -8726 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 592650 655954
rect -8726 655634 592650 655718
rect -8726 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 592650 655634
rect -8726 655366 592650 655398
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 646954 592650 646986
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect -8726 646634 592650 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect -8726 646366 592650 646398
rect -8726 642454 592650 642486
rect -8726 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 592650 642454
rect -8726 642134 592650 642218
rect -8726 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 592650 642134
rect -8726 641866 592650 641898
rect -8726 637954 592650 637986
rect -8726 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 592650 637954
rect -8726 637634 592650 637718
rect -8726 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 592650 637634
rect -8726 637366 592650 637398
rect -8726 633454 592650 633486
rect -8726 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 592650 633454
rect -8726 633134 592650 633218
rect -8726 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 592650 633134
rect -8726 632866 592650 632898
rect -8726 628954 592650 628986
rect -8726 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 592650 628954
rect -8726 628634 592650 628718
rect -8726 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 592650 628634
rect -8726 628366 592650 628398
rect -8726 624454 592650 624486
rect -8726 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 619954 592650 619986
rect -8726 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 592650 619954
rect -8726 619634 592650 619718
rect -8726 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 592650 619634
rect -8726 619366 592650 619398
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 610954 592650 610986
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect -8726 610634 592650 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect -8726 610366 592650 610398
rect -8726 606454 592650 606486
rect -8726 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 592650 606454
rect -8726 606134 592650 606218
rect -8726 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 592650 606134
rect -8726 605866 592650 605898
rect -8726 601954 592650 601986
rect -8726 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 592650 601954
rect -8726 601634 592650 601718
rect -8726 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 592650 601634
rect -8726 601366 592650 601398
rect -8726 597454 592650 597486
rect -8726 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 592650 597454
rect -8726 597134 592650 597218
rect -8726 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 592650 597134
rect -8726 596866 592650 596898
rect -8726 592954 592650 592986
rect -8726 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 592650 592954
rect -8726 592634 592650 592718
rect -8726 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 592650 592634
rect -8726 592366 592650 592398
rect -8726 588454 592650 588486
rect -8726 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 583954 592650 583986
rect -8726 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 592650 583954
rect -8726 583634 592650 583718
rect -8726 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 592650 583634
rect -8726 583366 592650 583398
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 574954 592650 574986
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect -8726 574634 592650 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect -8726 574366 592650 574398
rect -8726 570454 592650 570486
rect -8726 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 592650 570454
rect -8726 570134 592650 570218
rect -8726 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 592650 570134
rect -8726 569866 592650 569898
rect -8726 565954 592650 565986
rect -8726 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 592650 565954
rect -8726 565634 592650 565718
rect -8726 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 592650 565634
rect -8726 565366 592650 565398
rect -8726 561454 592650 561486
rect -8726 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 592650 561454
rect -8726 561134 592650 561218
rect -8726 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 592650 561134
rect -8726 560866 592650 560898
rect -8726 556954 592650 556986
rect -8726 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 592650 556954
rect -8726 556634 592650 556718
rect -8726 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 592650 556634
rect -8726 556366 592650 556398
rect -8726 552454 592650 552486
rect -8726 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 592650 552454
rect -8726 552134 592650 552218
rect -8726 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 547954 592650 547986
rect -8726 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 592650 547954
rect -8726 547634 592650 547718
rect -8726 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 592650 547634
rect -8726 547366 592650 547398
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 538954 592650 538986
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect -8726 538634 592650 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect -8726 538366 592650 538398
rect -8726 534454 592650 534486
rect -8726 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 529954 592650 529986
rect -8726 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 592650 529954
rect -8726 529634 592650 529718
rect -8726 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 592650 529634
rect -8726 529366 592650 529398
rect -8726 525454 592650 525486
rect -8726 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 592650 525454
rect -8726 525134 592650 525218
rect -8726 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 592650 525134
rect -8726 524866 592650 524898
rect -8726 520954 592650 520986
rect -8726 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 592650 520954
rect -8726 520634 592650 520718
rect -8726 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 592650 520634
rect -8726 520366 592650 520398
rect -8726 516454 592650 516486
rect -8726 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 511954 592650 511986
rect -8726 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 592650 511954
rect -8726 511634 592650 511718
rect -8726 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 592650 511634
rect -8726 511366 592650 511398
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 502954 592650 502986
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect -8726 502634 592650 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect -8726 502366 592650 502398
rect -8726 498454 592650 498486
rect -8726 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 592650 498454
rect -8726 498134 592650 498218
rect -8726 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 592650 498134
rect -8726 497866 592650 497898
rect -8726 493954 592650 493986
rect -8726 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 592650 493954
rect -8726 493634 592650 493718
rect -8726 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 592650 493634
rect -8726 493366 592650 493398
rect -8726 489454 592650 489486
rect -8726 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 592650 489454
rect -8726 489134 592650 489218
rect -8726 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 592650 489134
rect -8726 488866 592650 488898
rect -8726 484954 592650 484986
rect -8726 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 592650 484954
rect -8726 484634 592650 484718
rect -8726 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 592650 484634
rect -8726 484366 592650 484398
rect -8726 480454 592650 480486
rect -8726 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 475954 592650 475986
rect -8726 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 592650 475954
rect -8726 475634 592650 475718
rect -8726 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 592650 475634
rect -8726 475366 592650 475398
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 466954 592650 466986
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect -8726 466634 592650 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect -8726 466366 592650 466398
rect -8726 462454 592650 462486
rect -8726 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 592650 462454
rect -8726 462134 592650 462218
rect -8726 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 592650 462134
rect -8726 461866 592650 461898
rect -8726 457954 592650 457986
rect -8726 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 592650 457954
rect -8726 457634 592650 457718
rect -8726 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 592650 457634
rect -8726 457366 592650 457398
rect -8726 453454 592650 453486
rect -8726 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 592650 453454
rect -8726 453134 592650 453218
rect -8726 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 592650 453134
rect -8726 452866 592650 452898
rect -8726 448954 592650 448986
rect -8726 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 592650 448954
rect -8726 448634 592650 448718
rect -8726 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 592650 448634
rect -8726 448366 592650 448398
rect -8726 444454 592650 444486
rect -8726 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 439954 592650 439986
rect -8726 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 592650 439954
rect -8726 439634 592650 439718
rect -8726 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 592650 439634
rect -8726 439366 592650 439398
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 430954 592650 430986
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect -8726 430634 592650 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect -8726 430366 592650 430398
rect -8726 426454 592650 426486
rect -8726 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 592650 426454
rect -8726 426134 592650 426218
rect -8726 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 592650 426134
rect -8726 425866 592650 425898
rect -8726 421954 592650 421986
rect -8726 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 592650 421954
rect -8726 421634 592650 421718
rect -8726 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 592650 421634
rect -8726 421366 592650 421398
rect -8726 417454 592650 417486
rect -8726 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 592650 417454
rect -8726 417134 592650 417218
rect -8726 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 592650 417134
rect -8726 416866 592650 416898
rect -8726 412954 592650 412986
rect -8726 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 592650 412954
rect -8726 412634 592650 412718
rect -8726 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 592650 412634
rect -8726 412366 592650 412398
rect -8726 408454 592650 408486
rect -8726 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 403954 592650 403986
rect -8726 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 592650 403954
rect -8726 403634 592650 403718
rect -8726 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 592650 403634
rect -8726 403366 592650 403398
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 394954 592650 394986
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect -8726 394634 592650 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect -8726 394366 592650 394398
rect -8726 390454 592650 390486
rect -8726 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 592650 390454
rect -8726 390134 592650 390218
rect -8726 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 592650 390134
rect -8726 389866 592650 389898
rect -8726 385954 592650 385986
rect -8726 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 592650 385954
rect -8726 385634 592650 385718
rect -8726 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 592650 385634
rect -8726 385366 592650 385398
rect -8726 381454 592650 381486
rect -8726 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 592650 381454
rect -8726 381134 592650 381218
rect -8726 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 592650 381134
rect -8726 380866 592650 380898
rect -8726 376954 592650 376986
rect -8726 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 592650 376954
rect -8726 376634 592650 376718
rect -8726 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 592650 376634
rect -8726 376366 592650 376398
rect -8726 372454 592650 372486
rect -8726 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 367954 592650 367986
rect -8726 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 592650 367954
rect -8726 367634 592650 367718
rect -8726 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 592650 367634
rect -8726 367366 592650 367398
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 358954 592650 358986
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect -8726 358634 592650 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect -8726 358366 592650 358398
rect -8726 354454 592650 354486
rect -8726 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 349954 592650 349986
rect -8726 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 592650 349954
rect -8726 349634 592650 349718
rect -8726 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 592650 349634
rect -8726 349366 592650 349398
rect -8726 345454 592650 345486
rect -8726 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 592650 345454
rect -8726 345134 592650 345218
rect -8726 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 592650 345134
rect -8726 344866 592650 344898
rect -8726 340954 592650 340986
rect -8726 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 592650 340954
rect -8726 340634 592650 340718
rect -8726 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 592650 340634
rect -8726 340366 592650 340398
rect -8726 336454 592650 336486
rect -8726 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 331954 592650 331986
rect -8726 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 592650 331954
rect -8726 331634 592650 331718
rect -8726 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 592650 331634
rect -8726 331366 592650 331398
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 322954 592650 322986
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect -8726 322634 592650 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect -8726 322366 592650 322398
rect -8726 318454 592650 318486
rect -8726 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 592650 318454
rect -8726 318134 592650 318218
rect -8726 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 592650 318134
rect -8726 317866 592650 317898
rect -8726 313954 592650 313986
rect -8726 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 592650 313954
rect -8726 313634 592650 313718
rect -8726 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 592650 313634
rect -8726 313366 592650 313398
rect -8726 309454 592650 309486
rect -8726 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 592650 309454
rect -8726 309134 592650 309218
rect -8726 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 592650 309134
rect -8726 308866 592650 308898
rect -8726 304954 592650 304986
rect -8726 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 592650 304954
rect -8726 304634 592650 304718
rect -8726 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 592650 304634
rect -8726 304366 592650 304398
rect -8726 300454 592650 300486
rect -8726 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 295954 592650 295986
rect -8726 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 592650 295954
rect -8726 295634 592650 295718
rect -8726 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 592650 295634
rect -8726 295366 592650 295398
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 286954 592650 286986
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect -8726 286634 592650 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect -8726 286366 592650 286398
rect -8726 282454 592650 282486
rect -8726 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 592650 282454
rect -8726 282134 592650 282218
rect -8726 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 592650 282134
rect -8726 281866 592650 281898
rect -8726 277954 592650 277986
rect -8726 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 592650 277954
rect -8726 277634 592650 277718
rect -8726 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 592650 277634
rect -8726 277366 592650 277398
rect -8726 273454 592650 273486
rect -8726 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 592650 273454
rect -8726 273134 592650 273218
rect -8726 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 592650 273134
rect -8726 272866 592650 272898
rect -8726 268954 592650 268986
rect -8726 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 592650 268954
rect -8726 268634 592650 268718
rect -8726 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 592650 268634
rect -8726 268366 592650 268398
rect -8726 264454 592650 264486
rect -8726 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 259954 592650 259986
rect -8726 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 592650 259954
rect -8726 259634 592650 259718
rect -8726 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 592650 259634
rect -8726 259366 592650 259398
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 124250 255454
rect 124486 255218 154970 255454
rect 155206 255218 185690 255454
rect 185926 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 124250 255134
rect 124486 254898 154970 255134
rect 155206 254898 185690 255134
rect 185926 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 250954 592650 250986
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect -8726 250634 592650 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect -8726 250366 592650 250398
rect -8726 246454 592650 246486
rect -8726 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 592650 246454
rect -8726 246134 592650 246218
rect -8726 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 592650 246134
rect -8726 245866 592650 245898
rect -8726 241954 592650 241986
rect -8726 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 592650 241954
rect -8726 241634 592650 241718
rect -8726 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 592650 241634
rect -8726 241366 592650 241398
rect -8726 237454 592650 237486
rect -8726 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 592650 237454
rect -8726 237134 592650 237218
rect -8726 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 592650 237134
rect -8726 236866 592650 236898
rect -8726 232954 592650 232986
rect -8726 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 592650 232954
rect -8726 232634 592650 232718
rect -8726 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 592650 232634
rect -8726 232366 592650 232398
rect -8726 228454 592650 228486
rect -8726 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 592650 228454
rect -8726 228134 592650 228218
rect -8726 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 592650 228134
rect -8726 227866 592650 227898
rect -8726 223954 592650 223986
rect -8726 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 139610 223954
rect 139846 223718 170330 223954
rect 170566 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 592650 223954
rect -8726 223634 592650 223718
rect -8726 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 139610 223634
rect 139846 223398 170330 223634
rect 170566 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 592650 223634
rect -8726 223366 592650 223398
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 124250 219454
rect 124486 219218 154970 219454
rect 155206 219218 185690 219454
rect 185926 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 124250 219134
rect 124486 218898 154970 219134
rect 155206 218898 185690 219134
rect 185926 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 214954 592650 214986
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect -8726 214634 592650 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect -8726 214366 592650 214398
rect -8726 210454 592650 210486
rect -8726 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 592650 210454
rect -8726 210134 592650 210218
rect -8726 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 592650 210134
rect -8726 209866 592650 209898
rect -8726 205954 592650 205986
rect -8726 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 592650 205954
rect -8726 205634 592650 205718
rect -8726 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 592650 205634
rect -8726 205366 592650 205398
rect -8726 201454 592650 201486
rect -8726 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 592650 201454
rect -8726 201134 592650 201218
rect -8726 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 592650 201134
rect -8726 200866 592650 200898
rect -8726 196954 592650 196986
rect -8726 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 592650 196954
rect -8726 196634 592650 196718
rect -8726 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 592650 196634
rect -8726 196366 592650 196398
rect -8726 192454 592650 192486
rect -8726 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 187954 592650 187986
rect -8726 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 592650 187954
rect -8726 187634 592650 187718
rect -8726 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 592650 187634
rect -8726 187366 592650 187398
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 178954 592650 178986
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect -8726 178634 592650 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect -8726 178366 592650 178398
rect -8726 174454 592650 174486
rect -8726 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 169954 592650 169986
rect -8726 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 592650 169954
rect -8726 169634 592650 169718
rect -8726 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 592650 169634
rect -8726 169366 592650 169398
rect -8726 165454 592650 165486
rect -8726 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 592650 165454
rect -8726 165134 592650 165218
rect -8726 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 592650 165134
rect -8726 164866 592650 164898
rect -8726 160954 592650 160986
rect -8726 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 592650 160954
rect -8726 160634 592650 160718
rect -8726 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 592650 160634
rect -8726 160366 592650 160398
rect -8726 156454 592650 156486
rect -8726 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 151954 592650 151986
rect -8726 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 592650 151954
rect -8726 151634 592650 151718
rect -8726 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 592650 151634
rect -8726 151366 592650 151398
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 142954 592650 142986
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect -8726 142634 592650 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect -8726 142366 592650 142398
rect -8726 138454 592650 138486
rect -8726 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 592650 138454
rect -8726 138134 592650 138218
rect -8726 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 592650 138134
rect -8726 137866 592650 137898
rect -8726 133954 592650 133986
rect -8726 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 592650 133954
rect -8726 133634 592650 133718
rect -8726 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 592650 133634
rect -8726 133366 592650 133398
rect -8726 129454 592650 129486
rect -8726 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 592650 129454
rect -8726 129134 592650 129218
rect -8726 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 592650 129134
rect -8726 128866 592650 128898
rect -8726 124954 592650 124986
rect -8726 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 592650 124954
rect -8726 124634 592650 124718
rect -8726 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 592650 124634
rect -8726 124366 592650 124398
rect -8726 120454 592650 120486
rect -8726 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 115954 592650 115986
rect -8726 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 139610 115954
rect 139846 115718 170330 115954
rect 170566 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 592650 115954
rect -8726 115634 592650 115718
rect -8726 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 139610 115634
rect 139846 115398 170330 115634
rect 170566 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 592650 115634
rect -8726 115366 592650 115398
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 124250 111454
rect 124486 111218 154970 111454
rect 155206 111218 185690 111454
rect 185926 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 124250 111134
rect 124486 110898 154970 111134
rect 155206 110898 185690 111134
rect 185926 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 106954 592650 106986
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect -8726 106634 592650 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect -8726 106366 592650 106398
rect -8726 102454 592650 102486
rect -8726 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 592650 102454
rect -8726 102134 592650 102218
rect -8726 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 592650 102134
rect -8726 101866 592650 101898
rect -8726 97954 592650 97986
rect -8726 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 592650 97954
rect -8726 97634 592650 97718
rect -8726 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 592650 97634
rect -8726 97366 592650 97398
rect -8726 93454 592650 93486
rect -8726 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 592650 93454
rect -8726 93134 592650 93218
rect -8726 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 592650 93134
rect -8726 92866 592650 92898
rect -8726 88954 592650 88986
rect -8726 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 592650 88954
rect -8726 88634 592650 88718
rect -8726 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 592650 88634
rect -8726 88366 592650 88398
rect -8726 84454 592650 84486
rect -8726 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 79954 592650 79986
rect -8726 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 592650 79954
rect -8726 79634 592650 79718
rect -8726 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 592650 79634
rect -8726 79366 592650 79398
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 70954 592650 70986
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect -8726 70634 592650 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect -8726 70366 592650 70398
rect -8726 66454 592650 66486
rect -8726 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 592650 66454
rect -8726 66134 592650 66218
rect -8726 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 592650 66134
rect -8726 65866 592650 65898
rect -8726 61954 592650 61986
rect -8726 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 592650 61954
rect -8726 61634 592650 61718
rect -8726 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 592650 61634
rect -8726 61366 592650 61398
rect -8726 57454 592650 57486
rect -8726 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 592650 57454
rect -8726 57134 592650 57218
rect -8726 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 592650 57134
rect -8726 56866 592650 56898
rect -8726 52954 592650 52986
rect -8726 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 592650 52954
rect -8726 52634 592650 52718
rect -8726 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 592650 52634
rect -8726 52366 592650 52398
rect -8726 48454 592650 48486
rect -8726 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 43954 592650 43986
rect -8726 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 592650 43954
rect -8726 43634 592650 43718
rect -8726 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 592650 43634
rect -8726 43366 592650 43398
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 34954 592650 34986
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect -8726 34634 592650 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect -8726 34366 592650 34398
rect -8726 30454 592650 30486
rect -8726 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 592650 30454
rect -8726 30134 592650 30218
rect -8726 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 592650 30134
rect -8726 29866 592650 29898
rect -8726 25954 592650 25986
rect -8726 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 592650 25954
rect -8726 25634 592650 25718
rect -8726 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 592650 25634
rect -8726 25366 592650 25398
rect -8726 21454 592650 21486
rect -8726 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 592650 21454
rect -8726 21134 592650 21218
rect -8726 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 592650 21134
rect -8726 20866 592650 20898
rect -8726 16954 592650 16986
rect -8726 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 592650 16954
rect -8726 16634 592650 16718
rect -8726 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 592650 16634
rect -8726 16366 592650 16398
rect -8726 12454 592650 12486
rect -8726 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 592650 12134
rect -8726 11866 592650 11898
rect -8726 7954 592650 7986
rect -8726 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 592650 7954
rect -8726 7634 592650 7718
rect -8726 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 592650 7634
rect -8726 7366 592650 7398
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use pixel_macro  pixel_macro0
timestamp 0
transform 1 0 120000 0 1 200000
box 1066 0 68854 60000
use rlbp_macro  rlbp_macro0
timestamp 0
transform 1 0 120000 0 1 80000
box 1066 0 68854 60000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 78000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 142000 146414 198000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 262000 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 78000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 142000 182414 198000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 262000 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 10794 -7654 11414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 -7654 47414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 -7654 83414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 -7654 119414 78000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 142000 119414 198000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 262000 119414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 -7654 155414 78000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 142000 155414 198000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 262000 155414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 -7654 191414 78000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 142000 191414 198000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 262000 191414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 -7654 227414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 -7654 263414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 -7654 299414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 -7654 335414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 -7654 371414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 -7654 407414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 -7654 443414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 -7654 479414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 -7654 515414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 550794 -7654 551414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 11866 592650 12486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 47866 592650 48486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 83866 592650 84486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 119866 592650 120486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 155866 592650 156486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 191866 592650 192486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 227866 592650 228486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 263866 592650 264486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 299866 592650 300486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 335866 592650 336486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 371866 592650 372486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 407866 592650 408486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 443866 592650 444486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 479866 592650 480486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 515866 592650 516486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 551866 592650 552486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 587866 592650 588486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 623866 592650 624486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 659866 592650 660486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 695866 592650 696486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 19794 -7654 20414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 -7654 56414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 -7654 92414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 -7654 128414 78000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 262000 128414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 -7654 164414 78000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 262000 164414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 -7654 200414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 -7654 236414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 -7654 272414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 -7654 308414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 -7654 344414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 -7654 380414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 -7654 416414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 451794 -7654 452414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 -7654 488414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 523794 -7654 524414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 559794 -7654 560414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 20866 592650 21486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 56866 592650 57486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 92866 592650 93486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 128866 592650 129486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 164866 592650 165486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 200866 592650 201486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 236866 592650 237486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 272866 592650 273486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 308866 592650 309486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 344866 592650 345486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 380866 592650 381486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 416866 592650 417486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 452866 592650 453486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 488866 592650 489486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 524866 592650 525486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 560866 592650 561486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 596866 592650 597486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 632866 592650 633486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 668866 592650 669486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 28794 -7654 29414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 -7654 65414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 -7654 101414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 -7654 137414 78000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 262000 137414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 -7654 173414 78000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 262000 173414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 -7654 209414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 -7654 245414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 -7654 281414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 -7654 317414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 -7654 353414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 -7654 389414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 424794 -7654 425414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 460794 -7654 461414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 496794 -7654 497414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 532794 -7654 533414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 568794 -7654 569414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 29866 592650 30486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 65866 592650 66486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 101866 592650 102486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 137866 592650 138486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 173866 592650 174486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 209866 592650 210486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 245866 592650 246486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 281866 592650 282486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 317866 592650 318486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 353866 592650 354486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 389866 592650 390486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 425866 592650 426486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 461866 592650 462486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 497866 592650 498486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 533866 592650 534486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 569866 592650 570486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 605866 592650 606486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 641866 592650 642486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 677866 592650 678486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 24294 -7654 24914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 -7654 60914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 -7654 96914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 -7654 132914 78000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 262000 132914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 -7654 168914 78000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 262000 168914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 -7654 204914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 -7654 240914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 -7654 276914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 -7654 312914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 -7654 348914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 -7654 384914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 -7654 420914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 456294 -7654 456914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 492294 -7654 492914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 528294 -7654 528914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 564294 -7654 564914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 25366 592650 25986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 61366 592650 61986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 97366 592650 97986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 133366 592650 133986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 169366 592650 169986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 205366 592650 205986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 241366 592650 241986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 277366 592650 277986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 313366 592650 313986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 349366 592650 349986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 385366 592650 385986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 421366 592650 421986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 457366 592650 457986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 493366 592650 493986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 529366 592650 529986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 565366 592650 565986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 601366 592650 601986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 637366 592650 637986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 673366 592650 673986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 33294 -7654 33914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 -7654 69914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 -7654 105914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 -7654 141914 78000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 142000 141914 198000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 262000 141914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 -7654 177914 78000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 142000 177914 198000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 262000 177914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 -7654 213914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 -7654 249914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 -7654 285914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 -7654 321914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 -7654 357914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 -7654 393914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 -7654 429914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 465294 -7654 465914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 -7654 501914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 537294 -7654 537914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 573294 -7654 573914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 34366 592650 34986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 70366 592650 70986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 106366 592650 106986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 142366 592650 142986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 178366 592650 178986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 214366 592650 214986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 250366 592650 250986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 286366 592650 286986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 322366 592650 322986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 358366 592650 358986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 394366 592650 394986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 430366 592650 430986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 466366 592650 466986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 502366 592650 502986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 538366 592650 538986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 574366 592650 574986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 610366 592650 610986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 646366 592650 646986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 682366 592650 682986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 6294 -7654 6914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 42294 -7654 42914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 -7654 78914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 -7654 114914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 -7654 150914 78000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 142000 150914 198000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 262000 150914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 -7654 186914 78000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 142000 186914 198000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 262000 186914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 -7654 222914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 -7654 258914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 -7654 294914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 -7654 330914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 -7654 366914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 -7654 402914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 -7654 438914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 -7654 474914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 -7654 510914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 546294 -7654 546914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 582294 -7654 582914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 7366 592650 7986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 43366 592650 43986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 79366 592650 79986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 115366 592650 115986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 151366 592650 151986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 187366 592650 187986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 223366 592650 223986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 259366 592650 259986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 295366 592650 295986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 331366 592650 331986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 367366 592650 367986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 403366 592650 403986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 439366 592650 439986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 475366 592650 475986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 511366 592650 511986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 547366 592650 547986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 583366 592650 583986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 619366 592650 619986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 655366 592650 655986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 691366 592650 691986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 15294 -7654 15914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 -7654 51914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 -7654 87914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 -7654 123914 78000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 142000 123914 198000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 262000 123914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 -7654 159914 78000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 142000 159914 198000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 262000 159914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 -7654 195914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 -7654 231914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 -7654 267914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 -7654 303914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 -7654 339914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 -7654 375914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 -7654 411914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 -7654 447914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 -7654 483914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 -7654 519914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 555294 -7654 555914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 16366 592650 16986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 52366 592650 52986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 88366 592650 88986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 124366 592650 124986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 160366 592650 160986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 196366 592650 196986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 232366 592650 232986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 268366 592650 268986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 304366 592650 304986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 340366 592650 340986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 376366 592650 376986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 412366 592650 412986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 448366 592650 448986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 484366 592650 484986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 520366 592650 520986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 556366 592650 556986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 592366 592650 592986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 628366 592650 628986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 664366 592650 664986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 700366 592650 700986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
