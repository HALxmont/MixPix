* NGSPICE file created from rlbp_macro.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtn_1 abstract view
.subckt sky130_fd_sc_hd__dlxtn_1 D GATE_N VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtn_2 abstract view
.subckt sky130_fd_sc_hd__dlxtn_2 D GATE_N VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_1 abstract view
.subckt sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
.ends

.subckt rlbp_macro CLR CMP CMP_out_c OTA_out_c OTA_sh_c Pd10_a Pd10_b Pd11_a Pd11_b
+ Pd12_a Pd12_b Pd1_a Pd1_b Pd2_a Pd2_b Pd3_a Pd3_b Pd4_a Pd4_b Pd5_a Pd5_b Pd6_a
+ Pd6_b Pd7_a Pd7_b Pd8_a Pd8_b Pd9_a Pd9_b SH_out_c Sh Sh_cmp Sh_rst Sw1 Sw2 Vd1
+ Vd2 Vref_cmp_c Vref_sel_c io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ irq[0] irq[1] irq[2] la_data_in[0] la_data_in[100] la_data_in[101] la_data_in[102]
+ la_data_in[103] la_data_in[104] la_data_in[105] la_data_in[106] la_data_in[107]
+ la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111] la_data_in[112]
+ la_data_in[113] la_data_in[114] la_data_in[115] la_data_in[116] la_data_in[117]
+ la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122]
+ la_data_in[123] la_data_in[124] la_data_in[125] la_data_in[126] la_data_in[127]
+ la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16] la_data_in[17]
+ la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21] la_data_in[22]
+ la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27] la_data_in[28]
+ la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32] la_data_in[33]
+ la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38] la_data_in[39]
+ la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43] la_data_in[44]
+ la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49] la_data_in[4]
+ la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54] la_data_in[55]
+ la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5] la_data_in[60]
+ la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64] la_data_in[65] la_data_in[66]
+ la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6] la_data_in[70] la_data_in[71]
+ la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76] la_data_in[77]
+ la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80] la_data_in[81] la_data_in[82]
+ la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86] la_data_in[87] la_data_in[88]
+ la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91] la_data_in[92] la_data_in[93]
+ la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98] la_data_in[99]
+ la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89]
+ la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110]
+ la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117]
+ la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123]
+ la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65]
+ la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71]
+ la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78]
+ la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84]
+ la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90]
+ la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97]
+ la_oenb[98] la_oenb[99] la_oenb[9] vccd1 vssd1 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i
XFILLER_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3140__A1 _3343_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3155_ _3155_/A _3155_/B vssd1 vssd1 vccd1 vccd1 _3155_/X sky130_fd_sc_hd__or2_1
XFILLER_82_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2106_ _3362_/Q _2106_/B vssd1 vssd1 vccd1 vccd1 _2153_/B sky130_fd_sc_hd__xnor2_1
XFILLER_54_214 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3086_ _3482_/Q _3074_/X _3085_/X _3031_/X vssd1 vssd1 vccd1 vccd1 _3482_/D sky130_fd_sc_hd__o211a_1
XFILLER_39_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2037_ _3352_/Q _2037_/B vssd1 vssd1 vccd1 vccd1 _2091_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__2455__A _2576_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2939_ _2971_/A vssd1 vssd1 vccd1 vccd1 _2939_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2190__A _3395_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2706__A1 _3391_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1709__A hold5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_376 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_320 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2724_ _2762_/A _2726_/B vssd1 vssd1 vccd1 vccd1 _2724_/X sky130_fd_sc_hd__or2_1
X_2655_ _3373_/Q _2642_/X _2653_/X _2654_/X vssd1 vssd1 vccd1 vccd1 _3373_/D sky130_fd_sc_hd__o211a_1
XFILLER_8_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2586_ _2586_/A _2586_/B vssd1 vssd1 vccd1 vccd1 _2586_/X sky130_fd_sc_hd__or2_1
XFILLER_101_403 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3113__A1 _3389_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3207_ _3207_/A vssd1 vssd1 vccd1 vccd1 _3207_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1675__A1 _3509_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3138_ _3415_/Q _2754_/B _3134_/X _3137_/X vssd1 vssd1 vccd1 vccd1 _3138_/X sky130_fd_sc_hd__a211o_1
XFILLER_82_342 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_375 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3069_ _3337_/Q _2516_/A _2640_/A _3373_/Q _3068_/X vssd1 vssd1 vccd1 vccd1 _3070_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_35_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2913__A _2951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_464 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3104__B2 _3528_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_567 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2823__A _3183_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2918__A1 _3454_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2440_ _3236_/A vssd1 vssd1 vccd1 vccd1 _2568_/A sky130_fd_sc_hd__buf_2
XFILLER_96_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2371_ hold1/X vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__buf_2
XFILLER_96_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_12_net107_A clkbuf_2_3__f_net107/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2303__C1 _3467_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2733__A _2771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2707_ _2782_/A _2707_/B vssd1 vssd1 vccd1 vccd1 _2707_/X sky130_fd_sc_hd__or2_1
X_2638_ _2943_/A _2709_/B vssd1 vssd1 vccd1 vccd1 _2997_/A sky130_fd_sc_hd__nor2_1
XFILLER_99_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2569_ _3349_/Q _2556_/X _2568_/X _2566_/X vssd1 vssd1 vccd1 vccd1 _3349_/D sky130_fd_sc_hd__o211a_1
XFILLER_59_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2643__A _2679_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_24 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1706__B _3262_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input55_A wbs_dat_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1722__A _3490_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2818__A _2968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_534 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_515 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1940_ _3316_/Q _3304_/Q vssd1 vssd1 vccd1 vccd1 _1941_/B sky130_fd_sc_hd__and2b_1
X_1871_ _3417_/Q _2046_/B vssd1 vssd1 vccd1 vccd1 _1901_/C sky130_fd_sc_hd__or2_1
XANTENNA__2272__B _2407_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3541_ _3541_/D _2360_/X vssd1 vssd1 vccd1 vccd1 _3543_/D sky130_fd_sc_hd__dlxtn_1
X_3472_ _3474_/CLK _3472_/D vssd1 vssd1 vccd1 vccd1 _3472_/Q sky130_fd_sc_hd__dfxtp_1
X_2423_ _2834_/A vssd1 vssd1 vccd1 vccd1 _3225_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_69_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2354_ _3560_/D _2352_/X _2353_/X vssd1 vssd1 vccd1 vccd1 _3562_/D sky130_fd_sc_hd__a21bo_1
XFILLER_96_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2285_ _3472_/Q _2285_/B vssd1 vssd1 vccd1 vccd1 _2286_/B sky130_fd_sc_hd__and2b_1
XFILLER_37_353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_47 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_231 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3808_ _3808_/A vssd1 vssd1 vccd1 vccd1 _3808_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrlbp_macro_203 vssd1 vssd1 vccd1 vccd1 rlbp_macro_203/HI la_data_out[5] sky130_fd_sc_hd__conb_1
Xrlbp_macro_214 vssd1 vssd1 vccd1 vccd1 rlbp_macro_214/HI la_data_out[16] sky130_fd_sc_hd__conb_1
Xrlbp_macro_225 vssd1 vssd1 vccd1 vccd1 rlbp_macro_225/HI la_data_out[27] sky130_fd_sc_hd__conb_1
Xrlbp_macro_236 vssd1 vssd1 vccd1 vccd1 rlbp_macro_236/HI la_data_out[38] sky130_fd_sc_hd__conb_1
Xrlbp_macro_247 vssd1 vssd1 vccd1 vccd1 rlbp_macro_247/HI la_data_out[49] sky130_fd_sc_hd__conb_1
Xrlbp_macro_258 vssd1 vssd1 vccd1 vccd1 rlbp_macro_258/HI la_data_out[60] sky130_fd_sc_hd__conb_1
XFILLER_0_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_231 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrlbp_macro_269 vssd1 vssd1 vccd1 vccd1 rlbp_macro_269/HI la_data_out[71] sky130_fd_sc_hd__conb_1
XFILLER_87_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2638__A _2943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2373__A _2373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2070_ _2068_/A _2068_/B _2059_/X vssd1 vssd1 vccd1 vccd1 _2072_/A sky130_fd_sc_hd__a21bo_1
XFILLER_19_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2972_ _3473_/Q _2962_/X _2970_/X _2971_/X vssd1 vssd1 vccd1 vccd1 _3473_/D sky130_fd_sc_hd__o211a_1
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1923_ _1921_/Y _1922_/X _1851_/A vssd1 vssd1 vccd1 vccd1 _1923_/X sky130_fd_sc_hd__o21a_1
X_1854_ _1854_/A _1900_/A _1901_/B _1854_/D vssd1 vssd1 vccd1 vccd1 _1873_/A sky130_fd_sc_hd__and4_1
X_1785_ _1785_/A _1785_/B _1837_/A _1785_/D vssd1 vssd1 vccd1 vccd1 _1786_/B sky130_fd_sc_hd__nand4_1
X_3524_ _3528_/CLK _3524_/D vssd1 vssd1 vccd1 vccd1 _3524_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3455_ _3464_/CLK _3455_/D vssd1 vssd1 vccd1 vccd1 _3455_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2406_ _2404_/Y _2402_/Y _2407_/B _3808_/A _2381_/B vssd1 vssd1 vccd1 vccd1 _3304_/D
+ sky130_fd_sc_hd__a2111oi_2
X_3386_ _3387_/CLK _3386_/D vssd1 vssd1 vccd1 vccd1 _3386_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2337_ _3454_/Q _2329_/Y _2332_/Y _2334_/Y _2336_/Y vssd1 vssd1 vccd1 vccd1 _2338_/D
+ sky130_fd_sc_hd__o2111ai_1
XANTENNA__2458__A _2578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2268_ _3391_/Q _2268_/B vssd1 vssd1 vccd1 vccd1 _2269_/D sky130_fd_sc_hd__xnor2_1
XFILLER_84_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2199_ _3404_/Q _2294_/B vssd1 vssd1 vccd1 vccd1 _2233_/B sky130_fd_sc_hd__xnor2_1
XFILLER_65_492 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2193__A _3394_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_518 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2921__A _2957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1711__B1 _1657_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input18_A la_data_in[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3199__A _3199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2831__A _3199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3240_ _3526_/Q _3224_/A _3238_/X _3239_/X vssd1 vssd1 vccd1 vccd1 _3518_/D sky130_fd_sc_hd__o211a_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3171_ _3184_/A vssd1 vssd1 vccd1 vccd1 _3171_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2122_ _2169_/A _2150_/B vssd1 vssd1 vccd1 vccd1 _2132_/A sky130_fd_sc_hd__and2_1
XFILLER_66_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2053_ _2073_/A _2074_/B _2052_/X vssd1 vssd1 vccd1 vccd1 _2080_/B sky130_fd_sc_hd__a21o_1
XFILLER_47_492 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_495 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2955_ _2955_/A _2960_/B vssd1 vssd1 vccd1 vccd1 _2955_/X sky130_fd_sc_hd__or2_1
XANTENNA__2741__A _2780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1906_ _1906_/A _1906_/B vssd1 vssd1 vccd1 vccd1 _1906_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__2430__A1 _3309_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2886_ _2960_/A _2886_/B vssd1 vssd1 vccd1 vccd1 _2886_/X sky130_fd_sc_hd__or2_1
X_1837_ _1837_/A _1837_/B vssd1 vssd1 vccd1 vccd1 _1838_/B sky130_fd_sc_hd__xor2_1
X_1768_ _3304_/Q vssd1 vssd1 vccd1 vccd1 _2145_/A sky130_fd_sc_hd__clkbuf_2
X_3507_ _3507_/CLK _3507_/D vssd1 vssd1 vccd1 vccd1 _3507_/Q sky130_fd_sc_hd__dfxtp_1
X_1699_ _3297_/Q vssd1 vssd1 vccd1 vccd1 _2389_/C sky130_fd_sc_hd__buf_2
X_3438_ _3450_/CLK _3438_/D vssd1 vssd1 vccd1 vccd1 _3438_/Q sky130_fd_sc_hd__dfxtp_1
X_3369_ _3377_/CLK _3369_/D vssd1 vssd1 vccd1 vccd1 _3369_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3143__C1 _3142_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_15_net107 clkbuf_2_3__f_net107/X vssd1 vssd1 vccd1 vccd1 _3392_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_38_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_602 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2406__D1 _2381_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2651__A _2762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput75 _3784_/X vssd1 vssd1 vccd1 vccd1 Pd12_a sky130_fd_sc_hd__buf_2
Xoutput97 _3295_/Q vssd1 vssd1 vccd1 vccd1 Sh_cmp sky130_fd_sc_hd__buf_2
Xoutput86 _3795_/X vssd1 vssd1 vccd1 vccd1 Pd5_b sky130_fd_sc_hd__buf_2
XFILLER_95_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2098__A _3343_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2488__A1 _3323_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2826__A _3186_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_37_net107_A _3494_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2740_ _3402_/Q _2728_/X _2739_/X _2731_/X vssd1 vssd1 vccd1 vccd1 _3402_/D sky130_fd_sc_hd__o211a_1
XANTENNA__2561__A _2561_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2671_ _3379_/Q _2656_/A _2670_/X _2668_/X vssd1 vssd1 vccd1 vccd1 _3379_/D sky130_fd_sc_hd__o211a_1
XFILLER_75_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3223_ _3223_/A _3225_/B vssd1 vssd1 vccd1 vccd1 _3224_/A sky130_fd_sc_hd__and2_1
XFILLER_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3140__A2 _2516_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3154_ _3320_/Q _2988_/A _3146_/X _3153_/X vssd1 vssd1 vccd1 vccd1 _3155_/B sky130_fd_sc_hd__a211o_1
X_2105_ _3361_/Q _2105_/B vssd1 vssd1 vccd1 vccd1 _2155_/A sky130_fd_sc_hd__xnor2_1
XFILLER_54_226 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3085_ _3121_/A _3085_/B vssd1 vssd1 vccd1 vccd1 _3085_/X sky130_fd_sc_hd__or2_1
XFILLER_82_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2036_ _2068_/A _2071_/B vssd1 vssd1 vccd1 vccd1 _2041_/A sky130_fd_sc_hd__and2_1
XFILLER_35_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2938_ _2975_/A _2941_/B vssd1 vssd1 vccd1 vccd1 _2938_/X sky130_fd_sc_hd__or2_1
XANTENNA__2471__A _3160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2190__B _2190_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2869_ _3440_/Q _2853_/A _2868_/X _2864_/X vssd1 vssd1 vccd1 vccd1 _3440_/D sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_2_net107 _3494_/CLK vssd1 vssd1 vccd1 vccd1 _3308_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_2_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_535 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2381__A _3808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1725__A _3498_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2275__B _2301_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2291__A _3475_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2723_ _3395_/Q _2713_/X _2722_/X _2718_/X vssd1 vssd1 vccd1 vccd1 _3395_/D sky130_fd_sc_hd__o211a_1
X_2654_ _2654_/A vssd1 vssd1 vccd1 vccd1 _2654_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2585_ _3355_/Q _2570_/A _2584_/X _2580_/X vssd1 vssd1 vccd1 vccd1 _3355_/D sky130_fd_sc_hd__o211a_1
XFILLER_101_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3113__A2 _3053_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3206_ _2568_/A _3191_/X _3205_/Y _3200_/X vssd1 vssd1 vccd1 vccd1 _3505_/D sky130_fd_sc_hd__o211a_1
XFILLER_55_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1675__A2 _2313_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3137_ _3355_/Q _2554_/A _3135_/X _3136_/X vssd1 vssd1 vccd1 vccd1 _3137_/X sky130_fd_sc_hd__a211o_1
XFILLER_82_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_387 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3068_ _3385_/Q _3053_/X _3033_/A _3525_/Q vssd1 vssd1 vccd1 vccd1 _3068_/X sky130_fd_sc_hd__a22o_1
XFILLER_42_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2019_ _3332_/Q _2019_/B vssd1 vssd1 vccd1 vccd1 _2020_/B sky130_fd_sc_hd__xor2_1
XFILLER_23_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_476 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_347 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3104__A2 _3053_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2376__A _3282_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3040__A1 _3323_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3040__B2 _3407_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2370_ _2742_/A vssd1 vssd1 vccd1 vccd1 _2370_/X sky130_fd_sc_hd__buf_2
XANTENNA__2054__A_N _3347_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2303__B1 _1678_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2706_ _3391_/Q _2692_/A _2705_/X _2699_/X vssd1 vssd1 vccd1 vccd1 _3391_/D sky130_fd_sc_hd__o211a_1
X_2637_ _3160_/A vssd1 vssd1 vccd1 vccd1 _2788_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_99_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2568_ _2568_/A _2568_/B vssd1 vssd1 vccd1 vccd1 _2568_/X sky130_fd_sc_hd__or2_1
XFILLER_101_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2499_ _2576_/A _2505_/B vssd1 vssd1 vccd1 vccd1 _2499_/X sky130_fd_sc_hd__or2_1
XFILLER_101_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_267 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2845__A1 _3430_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2643__B _2643_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3022__A1 _3346_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3022__B2 _3430_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_36 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input48_A wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3089__B2 _3527_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_546 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3261__A1 _3527_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1870_ _1870_/A _1870_/B vssd1 vssd1 vccd1 vccd1 _1928_/A sky130_fd_sc_hd__nor2_1
X_3540_ _3540_/D _2360_/X vssd1 vssd1 vccd1 vccd1 _3540_/Q sky130_fd_sc_hd__dlxtn_2
X_3471_ _3474_/CLK _3471_/D vssd1 vssd1 vccd1 vccd1 _3471_/Q sky130_fd_sc_hd__dfxtp_1
X_2422_ _2470_/A vssd1 vssd1 vccd1 vccd1 _2834_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_43_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2353_ _2353_/A _3564_/Q _3563_/Q vssd1 vssd1 vccd1 vccd1 _2353_/X sky130_fd_sc_hd__or3b_1
XFILLER_96_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2284_ _2285_/B _3472_/Q vssd1 vssd1 vccd1 vccd1 _2286_/A sky130_fd_sc_hd__and2b_1
XFILLER_37_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_538 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2055__A2 _1698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_59 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3807_ _3807_/A vssd1 vssd1 vccd1 vccd1 _3807_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3004__A1 _3393_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1999_ _1999_/A _1999_/B vssd1 vssd1 vccd1 vccd1 _2000_/B sky130_fd_sc_hd__xnor2_1
Xrlbp_macro_215 vssd1 vssd1 vccd1 vccd1 rlbp_macro_215/HI la_data_out[17] sky130_fd_sc_hd__conb_1
Xrlbp_macro_204 vssd1 vssd1 vccd1 vccd1 rlbp_macro_204/HI la_data_out[6] sky130_fd_sc_hd__conb_1
Xrlbp_macro_226 vssd1 vssd1 vccd1 vccd1 rlbp_macro_226/HI la_data_out[28] sky130_fd_sc_hd__conb_1
Xrlbp_macro_237 vssd1 vssd1 vccd1 vccd1 rlbp_macro_237/HI la_data_out[39] sky130_fd_sc_hd__conb_1
Xrlbp_macro_248 vssd1 vssd1 vccd1 vccd1 rlbp_macro_248/HI la_data_out[50] sky130_fd_sc_hd__conb_1
XANTENNA__2919__A _2955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_243 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrlbp_macro_259 vssd1 vssd1 vccd1 vccd1 rlbp_macro_259/HI la_data_out[61] sky130_fd_sc_hd__conb_1
XANTENNA__1937__A_N _2288_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2638__B _2709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2829__A _3188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_276 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2971_ _2971_/A vssd1 vssd1 vccd1 vccd1 _2971_/X sky130_fd_sc_hd__buf_2
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1922_ _1922_/A vssd1 vssd1 vccd1 vccd1 _1922_/X sky130_fd_sc_hd__clkbuf_4
X_1853_ _1911_/A _1893_/B vssd1 vssd1 vccd1 vccd1 _1854_/D sky130_fd_sc_hd__and2_1
XANTENNA__1908__A _3407_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1784_ _3294_/Q _3293_/Q _1840_/B _1813_/C vssd1 vssd1 vccd1 vccd1 _1785_/D sky130_fd_sc_hd__and4b_1
X_3523_ _3528_/CLK _3523_/D vssd1 vssd1 vccd1 vccd1 _3523_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_6_291 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3454_ _3464_/CLK _3454_/D vssd1 vssd1 vccd1 vccd1 _3454_/Q sky130_fd_sc_hd__dfxtp_1
X_2405_ _2405_/A _2405_/B _2405_/C vssd1 vssd1 vccd1 vccd1 _2407_/B sky130_fd_sc_hd__and3_1
XFILLER_97_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3385_ _3387_/CLK _3385_/D vssd1 vssd1 vccd1 vccd1 _3385_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2739__A _2778_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2336_ _3455_/Q _2336_/B vssd1 vssd1 vccd1 vccd1 _2336_/Y sky130_fd_sc_hd__xnor2_1
X_2267_ _2267_/A _2267_/B vssd1 vssd1 vccd1 vccd1 _2268_/B sky130_fd_sc_hd__xnor2_1
XFILLER_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2198_ _2249_/A _2251_/B _2198_/C vssd1 vssd1 vccd1 vccd1 _2213_/B sky130_fd_sc_hd__and3_1
XFILLER_25_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2433__C1 _2370_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_38_net107 _3494_/CLK vssd1 vssd1 vccd1 vccd1 _3332_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_96_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2649__A _2760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1711__A1 _3499_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1711__B2 _3492_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3216__A1 _2578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output79_A _3788_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2559__A _2559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2278__B _3300_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3170_ _3236_/A _3170_/B vssd1 vssd1 vccd1 vccd1 _3170_/X sky130_fd_sc_hd__or2_1
XFILLER_39_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2121_ _3366_/Q _2121_/B vssd1 vssd1 vccd1 vccd1 _2150_/B sky130_fd_sc_hd__xnor2_1
XFILLER_39_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2052_ _3346_/Q _2052_/B vssd1 vssd1 vccd1 vccd1 _2052_/X sky130_fd_sc_hd__and2b_1
XFILLER_81_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2954_ _3466_/Q _2948_/X _2953_/X _2939_/X vssd1 vssd1 vccd1 vccd1 _3466_/D sky130_fd_sc_hd__o211a_1
X_1905_ _3408_/Q _1905_/B vssd1 vssd1 vccd1 vccd1 _1906_/B sky130_fd_sc_hd__xnor2_1
X_2885_ _3444_/Q _2874_/X _2884_/X _2882_/X vssd1 vssd1 vccd1 vccd1 _3444_/D sky130_fd_sc_hd__o211a_1
X_1836_ _1833_/Y _1834_/X _1762_/D _1827_/B _1835_/X vssd1 vssd1 vccd1 vccd1 _1837_/B
+ sky130_fd_sc_hd__a221o_1
X_1767_ _1810_/A _1808_/B vssd1 vssd1 vccd1 vccd1 _1776_/A sky130_fd_sc_hd__and2_1
X_3506_ _3511_/CLK _3506_/D vssd1 vssd1 vccd1 vccd1 _3506_/Q sky130_fd_sc_hd__dfxtp_1
X_1698_ _1698_/A vssd1 vssd1 vccd1 vccd1 _2395_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_89_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3437_ _3450_/CLK _3437_/D vssd1 vssd1 vccd1 vccd1 _3437_/Q sky130_fd_sc_hd__dfxtp_1
X_3368_ _3404_/CLK _3368_/D vssd1 vssd1 vccd1 vccd1 _3368_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2319_ _2339_/A _2339_/B _2313_/Y vssd1 vssd1 vccd1 vccd1 _2321_/A sky130_fd_sc_hd__a21o_1
XFILLER_57_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3299_ _3308_/CLK _3299_/D vssd1 vssd1 vccd1 vccd1 _3299_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_45_408 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2406__C1 _3808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2932__A _2968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput76 _3785_/X vssd1 vssd1 vccd1 vccd1 Pd12_b sky130_fd_sc_hd__buf_2
XFILLER_0_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput98 _3560_/Q vssd1 vssd1 vccd1 vccd1 Sh_rst sky130_fd_sc_hd__buf_2
Xoutput87 _3796_/X vssd1 vssd1 vccd1 vccd1 Pd6_a sky130_fd_sc_hd__buf_2
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input30_A la_data_in[33] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1730__B _2378_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2842__A _2951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2670_ _2780_/A _2672_/B vssd1 vssd1 vccd1 vccd1 _2670_/X sky130_fd_sc_hd__or2_1
XFILLER_8_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2280__C _2330_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_21_net107 _3436_/CLK vssd1 vssd1 vccd1 vccd1 _3427_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_4_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3222_ _2586_/A _3202_/B _3221_/X _3213_/X vssd1 vssd1 vccd1 vccd1 _3512_/D sky130_fd_sc_hd__o211a_1
XFILLER_79_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3153_ _3153_/A _3153_/B _3153_/C _3153_/D vssd1 vssd1 vccd1 vccd1 _3153_/X sky130_fd_sc_hd__or4_2
X_2104_ _3553_/Q _3554_/Q vssd1 vssd1 vccd1 vccd1 _2134_/A sky130_fd_sc_hd__or2b_1
XFILLER_39_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3084_ _3314_/Q _2993_/X _3076_/X _3083_/X vssd1 vssd1 vccd1 vccd1 _3085_/B sky130_fd_sc_hd__a211o_1
XFILLER_82_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2035_ _3350_/Q _2106_/B vssd1 vssd1 vccd1 vccd1 _2071_/B sky130_fd_sc_hd__xnor2_1
XFILLER_54_238 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2752__A _2788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2937_ _3462_/Q _2925_/X _2936_/X _2928_/X vssd1 vssd1 vccd1 vccd1 _3462_/D sky130_fd_sc_hd__o211a_1
X_2868_ _2977_/A _2868_/B vssd1 vssd1 vccd1 vccd1 _2868_/X sky130_fd_sc_hd__or2_1
X_1819_ _3432_/Q _1819_/B vssd1 vssd1 vccd1 vccd1 _1820_/B sky130_fd_sc_hd__xnor2_1
X_2799_ _3232_/A vssd1 vssd1 vccd1 vccd1 _2955_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_89_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2927__A _2964_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_547 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2662__A _2773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2381__B _2381_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2158__A1 _3359_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3107__B1 _3195_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2572__A _2572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2291__B _2291_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2722_ _2760_/A _2726_/B vssd1 vssd1 vccd1 vccd1 _2722_/X sky130_fd_sc_hd__or2_1
X_2653_ _2765_/A _2653_/B vssd1 vssd1 vccd1 vccd1 _2653_/X sky130_fd_sc_hd__or2_1
XANTENNA__1916__A _3411_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2584_ _2584_/A _2586_/B vssd1 vssd1 vccd1 vccd1 _2584_/X sky130_fd_sc_hd__or2_1
XFILLER_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3205_ _3205_/A _3219_/B vssd1 vssd1 vccd1 vccd1 _3205_/Y sky130_fd_sc_hd__nand2_1
X_3136_ _3331_/Q _2476_/A _3017_/X _3451_/Q vssd1 vssd1 vccd1 vccd1 _3136_/X sky130_fd_sc_hd__a22o_1
XFILLER_55_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3067_ _3397_/Q _3041_/X _3056_/A _3505_/Q _3066_/X vssd1 vssd1 vccd1 vccd1 _3070_/B
+ sky130_fd_sc_hd__a221o_1
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2018_ _1983_/A _1983_/B _1934_/A vssd1 vssd1 vccd1 vccd1 _2020_/A sky130_fd_sc_hd__o21ai_1
XFILLER_82_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2482__A _2559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_488 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1826__A _3435_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2560__A1 _3345_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2392__A _2395_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1814__B1 _3429_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_21_net107_A _3436_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2705_ _2780_/A _2707_/B vssd1 vssd1 vccd1 vccd1 _2705_/X sky130_fd_sc_hd__or2_1
X_2636_ _3368_/Q _2612_/A _2634_/X _2635_/X vssd1 vssd1 vccd1 vccd1 _3368_/D sky130_fd_sc_hd__o211a_1
X_2567_ _3348_/Q _2556_/X _2565_/X _2566_/X vssd1 vssd1 vccd1 vccd1 _3348_/D sky130_fd_sc_hd__o211a_1
XFILLER_87_436 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2498_ _3327_/Q _2493_/X _2497_/X _2487_/X vssd1 vssd1 vccd1 vccd1 _3327_/D sky130_fd_sc_hd__o211a_1
XFILLER_101_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2196__B _3306_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3274__A_N _2378_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3119_ _3119_/A _3119_/B _3119_/C vssd1 vssd1 vccd1 vccd1 _3119_/X sky130_fd_sc_hd__or3_1
XFILLER_43_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2781__A1 _3415_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1884__B_N _1794_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2850__A _2960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2772__A1 _3411_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3470_ _3474_/CLK _3470_/D vssd1 vssd1 vccd1 vccd1 _3470_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2421_ _2421_/A _2421_/B _3264_/B vssd1 vssd1 vccd1 vccd1 _2470_/A sky130_fd_sc_hd__and3_1
X_2352_ _2352_/A _2352_/B _2352_/C _2352_/D vssd1 vssd1 vccd1 vccd1 _2352_/X sky130_fd_sc_hd__or4_1
XFILLER_96_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2283_ _2333_/A _2323_/B vssd1 vssd1 vccd1 vccd1 _2290_/A sky130_fd_sc_hd__and2_1
XFILLER_96_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3806_ _3806_/A vssd1 vssd1 vccd1 vccd1 _3806_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2760__A _2760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3004__A2 _2711_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1998_ _1998_/A _1998_/B vssd1 vssd1 vccd1 vccd1 _1998_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_20_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2619_ _2654_/A vssd1 vssd1 vccd1 vccd1 _2619_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xrlbp_macro_205 vssd1 vssd1 vccd1 vccd1 rlbp_macro_205/HI la_data_out[7] sky130_fd_sc_hd__conb_1
Xrlbp_macro_238 vssd1 vssd1 vccd1 vccd1 rlbp_macro_238/HI la_data_out[40] sky130_fd_sc_hd__conb_1
Xrlbp_macro_227 vssd1 vssd1 vccd1 vccd1 rlbp_macro_227/HI la_data_out[29] sky130_fd_sc_hd__conb_1
Xrlbp_macro_216 vssd1 vssd1 vccd1 vccd1 rlbp_macro_216/HI la_data_out[18] sky130_fd_sc_hd__conb_1
Xrlbp_macro_249 vssd1 vssd1 vccd1 vccd1 rlbp_macro_249/HI la_data_out[51] sky130_fd_sc_hd__conb_1
XFILLER_87_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2000__A _3323_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2670__A _2780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2194__A_N _1949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input60_A wbs_dat_i[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3006__A _3006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2970_ _2970_/A _2973_/B vssd1 vssd1 vccd1 vccd1 _2970_/X sky130_fd_sc_hd__or2_1
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1921_ _3426_/Q vssd1 vssd1 vccd1 vccd1 _1921_/Y sky130_fd_sc_hd__inv_2
X_1852_ _3426_/Q _2121_/B vssd1 vssd1 vccd1 vccd1 _1893_/B sky130_fd_sc_hd__xnor2_1
X_1783_ _3441_/Q _2046_/B vssd1 vssd1 vccd1 vccd1 _1813_/C sky130_fd_sc_hd__or2_1
X_3522_ _3528_/CLK _3522_/D vssd1 vssd1 vccd1 vccd1 _3522_/Q sky130_fd_sc_hd__dfxtp_2
X_3453_ _3464_/CLK _3453_/D vssd1 vssd1 vccd1 vccd1 _3453_/Q sky130_fd_sc_hd__dfxtp_1
X_2404_ _2405_/A vssd1 vssd1 vccd1 vccd1 _2404_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3384_ _3387_/CLK _3384_/D vssd1 vssd1 vccd1 vccd1 _3384_/Q sky130_fd_sc_hd__dfxtp_1
X_2335_ _2335_/A _2335_/B vssd1 vssd1 vccd1 vccd1 _2336_/B sky130_fd_sc_hd__xor2_1
XFILLER_97_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2266_ _2258_/Y _2259_/X _2262_/X _2263_/Y _2265_/Y vssd1 vssd1 vccd1 vccd1 _2269_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_69_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2197_ _2264_/A _2241_/B vssd1 vssd1 vccd1 vccd1 _2198_/C sky130_fd_sc_hd__and2_1
XFILLER_65_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2474__B _2943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2736__A1 _3400_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_520 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2727__A1 _3397_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3152__B2 _3440_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2120_ _2120_/A _2120_/B vssd1 vssd1 vccd1 vccd1 _2169_/A sky130_fd_sc_hd__nor2_1
X_2051_ _3348_/Q vssd1 vssd1 vccd1 vccd1 _2051_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2294__B _2294_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2953_ _2953_/A _2960_/B vssd1 vssd1 vccd1 vccd1 _2953_/X sky130_fd_sc_hd__or2_1
X_1904_ _1907_/A _1907_/B _1881_/X vssd1 vssd1 vccd1 vccd1 _1906_/A sky130_fd_sc_hd__a21oi_1
X_2884_ _2957_/A _2886_/B vssd1 vssd1 vccd1 vccd1 _2884_/X sky130_fd_sc_hd__or2_1
X_1835_ _1833_/Y _1693_/A _1759_/A vssd1 vssd1 vccd1 vccd1 _1835_/X sky130_fd_sc_hd__o21a_1
XFILLER_30_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1766_ _3446_/Q _2106_/B vssd1 vssd1 vccd1 vccd1 _1808_/B sky130_fd_sc_hd__xnor2_1
X_3505_ _3507_/CLK _3505_/D vssd1 vssd1 vccd1 vccd1 _3505_/Q sky130_fd_sc_hd__dfxtp_1
X_1697_ _2026_/B vssd1 vssd1 vccd1 vccd1 _1698_/A sky130_fd_sc_hd__buf_2
XANTENNA__3143__A1 _3319_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3436_ _3436_/CLK _3436_/D vssd1 vssd1 vccd1 vccd1 _3436_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3367_ _3404_/CLK _3367_/D vssd1 vssd1 vccd1 vccd1 _3367_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2318_ _2318_/A _2318_/B vssd1 vssd1 vccd1 vccd1 _2352_/A sky130_fd_sc_hd__xnor2_1
X_3298_ _3356_/CLK _3298_/D vssd1 vssd1 vccd1 vccd1 _3298_/Q sky130_fd_sc_hd__dfxtp_1
X_2249_ _2249_/A _2251_/B vssd1 vssd1 vccd1 vccd1 _2250_/B sky130_fd_sc_hd__xnor2_1
XFILLER_26_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2379__B input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3134__A1 _3427_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput99 _3550_/Q vssd1 vssd1 vccd1 vccd1 Sw1 sky130_fd_sc_hd__buf_2
Xoutput77 _3786_/X vssd1 vssd1 vccd1 vccd1 Pd1_a sky130_fd_sc_hd__buf_2
Xoutput88 _3797_/X vssd1 vssd1 vccd1 vccd1 Pd6_b sky130_fd_sc_hd__buf_2
XANTENNA__3134__B2 _3511_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2395__A _2395_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input23_A la_data_in[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1739__A _3548_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2581__C1 _2580_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1923__A2 _1922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3221_ _3512_/Q _3221_/B vssd1 vssd1 vccd1 vccd1 _3221_/X sky130_fd_sc_hd__or2_1
XANTENNA__3125__B2 _3510_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3152_ _3428_/Q _2786_/A _2837_/A _3440_/Q _3151_/X vssd1 vssd1 vccd1 vccd1 _3153_/D
+ sky130_fd_sc_hd__a221o_1
X_2103_ _2049_/A _2102_/X _2049_/B vssd1 vssd1 vccd1 vccd1 _3547_/D sky130_fd_sc_hd__o21ai_1
X_3083_ _3083_/A _3083_/B _3083_/C _3083_/D vssd1 vssd1 vccd1 vccd1 _3083_/X sky130_fd_sc_hd__or4_1
X_2034_ _3349_/Q _2281_/B vssd1 vssd1 vccd1 vccd1 _2068_/A sky130_fd_sc_hd__xnor2_1
XFILLER_23_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1649__A _3511_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2936_ _2973_/A _2936_/B vssd1 vssd1 vccd1 vccd1 _2936_/X sky130_fd_sc_hd__or2_1
X_2867_ _3439_/Q _2853_/A _2866_/X _2864_/X vssd1 vssd1 vccd1 vccd1 _3439_/D sky130_fd_sc_hd__o211a_1
X_1818_ _1816_/A _1816_/B _1791_/X vssd1 vssd1 vccd1 vccd1 _1820_/A sky130_fd_sc_hd__a21oi_1
X_2798_ _3418_/Q _2789_/X _2796_/X _2797_/X vssd1 vssd1 vccd1 vccd1 _3418_/D sky130_fd_sc_hd__o211a_1
X_1749_ _1749_/A vssd1 vssd1 vccd1 vccd1 _1749_/X sky130_fd_sc_hd__buf_1
XFILLER_89_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2199__B _2294_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3419_ _3476_/CLK _3419_/D vssd1 vssd1 vccd1 vccd1 _3419_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3116__A1 _3413_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2943__A _2943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_423 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2158__A2 _1678_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3107__A1 _3400_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3107__B2 _3508_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2128__A_N _3360_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2721_ _3394_/Q _2713_/X _2720_/X _2718_/X vssd1 vssd1 vccd1 vccd1 _3394_/D sky130_fd_sc_hd__o211a_1
X_2652_ _3372_/Q _2642_/X _2651_/X _2635_/X vssd1 vssd1 vccd1 vccd1 _3372_/D sky130_fd_sc_hd__o211a_1
XFILLER_8_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2583_ _3354_/Q _2570_/X _2582_/X _2580_/X vssd1 vssd1 vccd1 vccd1 _3354_/D sky130_fd_sc_hd__o211a_1
XANTENNA__1932__A _3319_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3204_ _3207_/A vssd1 vssd1 vccd1 vccd1 _3219_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3135_ _3379_/Q _2997_/X _2711_/A _3403_/Q vssd1 vssd1 vccd1 vccd1 _3135_/X sky130_fd_sc_hd__a22o_1
XFILLER_27_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3066_ _3349_/Q _3000_/X _2837_/A _3433_/Q vssd1 vssd1 vccd1 vccd1 _3066_/X sky130_fd_sc_hd__a22o_1
XFILLER_70_518 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2017_ _2008_/Y _2009_/X _2012_/X _2013_/Y _2016_/Y vssd1 vssd1 vccd1 vccd1 _2021_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_50_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2919_ _2955_/A _2923_/B vssd1 vssd1 vccd1 vccd1 _2919_/X sky130_fd_sc_hd__or2_1
XANTENNA__2003__A _3322_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2938__A _2975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_450 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_570 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2848__A _2957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2303__A2 _1657_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_8_net107_A clkbuf_leaf_9_net107/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2704_ _3390_/Q _2692_/X _2703_/X _2699_/X vssd1 vssd1 vccd1 vccd1 _3390_/D sky130_fd_sc_hd__o211a_1
X_2635_ _2654_/A vssd1 vssd1 vccd1 vccd1 _2635_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2566_ _2566_/A vssd1 vssd1 vccd1 vccd1 _2566_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_99_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2758__A _2758_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2497_ _2574_/A _2505_/B vssd1 vssd1 vccd1 vccd1 _2497_/X sky130_fd_sc_hd__or2_1
XFILLER_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3118_ _3437_/Q _3021_/X _2875_/B _3449_/Q _3117_/X vssd1 vssd1 vccd1 vccd1 _3119_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_43_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3049_ _3444_/Q _3017_/X _3018_/X _3492_/Q vssd1 vssd1 vccd1 vccd1 _3049_/X sky130_fd_sc_hd__a22o_1
XFILLER_36_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_286 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2420_ _2420_/A _2420_/B _2420_/C vssd1 vssd1 vccd1 vccd1 _3264_/B sky130_fd_sc_hd__and3_1
XFILLER_89_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2578__A _2578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2351_ _3463_/Q _2351_/B vssd1 vssd1 vccd1 vccd1 _2352_/D sky130_fd_sc_hd__xnor2_1
XFILLER_96_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2282_ _3470_/Q _2282_/B vssd1 vssd1 vccd1 vccd1 _2323_/B sky130_fd_sc_hd__xnor2_1
XFILLER_96_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3805_ _3805_/A vssd1 vssd1 vccd1 vccd1 _3805_/X sky130_fd_sc_hd__clkbuf_1
X_1997_ _3324_/Q _1997_/B vssd1 vssd1 vccd1 vccd1 _1998_/B sky130_fd_sc_hd__xnor2_1
XFILLER_20_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1657__A _2026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2618_ _2771_/A _2628_/B vssd1 vssd1 vccd1 vccd1 _2618_/X sky130_fd_sc_hd__or2_1
Xrlbp_macro_206 vssd1 vssd1 vccd1 vccd1 rlbp_macro_206/HI la_data_out[8] sky130_fd_sc_hd__conb_1
X_2549_ _2586_/A _2549_/B vssd1 vssd1 vccd1 vccd1 _2549_/X sky130_fd_sc_hd__or2_1
Xrlbp_macro_217 vssd1 vssd1 vccd1 vccd1 rlbp_macro_217/HI la_data_out[19] sky130_fd_sc_hd__conb_1
Xrlbp_macro_228 vssd1 vssd1 vccd1 vccd1 rlbp_macro_228/HI la_data_out[30] sky130_fd_sc_hd__conb_1
Xrlbp_macro_239 vssd1 vssd1 vccd1 vccd1 rlbp_macro_239/HI la_data_out[41] sky130_fd_sc_hd__conb_1
XFILLER_0_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_186 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_8_net107 clkbuf_leaf_9_net107/A vssd1 vssd1 vccd1 vccd1 _3528_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__2951__A _2951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3782__A _3782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input53_A wbs_dat_i[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3006__B _3006_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2978__C1 _2971_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1920_ _1920_/A _1920_/B _1920_/C _1920_/D vssd1 vssd1 vccd1 vccd1 _1930_/B sky130_fd_sc_hd__and4_1
XFILLER_15_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2861__A _2970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1851_ _1851_/A _1851_/B vssd1 vssd1 vccd1 vccd1 _1911_/A sky130_fd_sc_hd__nor2_1
XFILLER_30_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3521_ _3528_/CLK _3521_/D vssd1 vssd1 vccd1 vccd1 _3521_/Q sky130_fd_sc_hd__dfxtp_2
X_1782_ _3452_/Q _2042_/B vssd1 vssd1 vccd1 vccd1 _1840_/B sky130_fd_sc_hd__xnor2_2
X_3452_ _3452_/CLK _3452_/D vssd1 vssd1 vccd1 vccd1 _3452_/Q sky130_fd_sc_hd__dfxtp_1
X_3383_ _3387_/CLK _3383_/D vssd1 vssd1 vccd1 vccd1 _3383_/Q sky130_fd_sc_hd__dfxtp_1
X_2403_ _2405_/B _2405_/C _2402_/Y _2397_/X vssd1 vssd1 vccd1 vccd1 _3303_/D sky130_fd_sc_hd__o211a_1
XFILLER_69_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2334_ _3457_/Q _2334_/B vssd1 vssd1 vccd1 vccd1 _2334_/Y sky130_fd_sc_hd__xnor2_1
X_2265_ _3389_/Q _2265_/B vssd1 vssd1 vccd1 vccd1 _2265_/Y sky130_fd_sc_hd__xnor2_1
X_2196_ _3402_/Q _3306_/Q vssd1 vssd1 vccd1 vccd1 _2241_/B sky130_fd_sc_hd__xnor2_1
XFILLER_37_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2771__A _2771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2433__A1 _3310_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3146__C1 _3145_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_495 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_307 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2681__A _2756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2050_ _2050_/A vssd1 vssd1 vccd1 vccd1 _3546_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2663__A1 _3376_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2415__A1 _2042_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_370 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2952_ _3465_/Q _2948_/X _2951_/X _2939_/X vssd1 vssd1 vccd1 vccd1 _3465_/D sky130_fd_sc_hd__o211a_1
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1903_ _3406_/Q _1900_/Y _1901_/X _1902_/Y vssd1 vssd1 vccd1 vccd1 _1903_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_30_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2883_ _3443_/Q _2874_/X _2881_/X _2882_/X vssd1 vssd1 vccd1 vccd1 _3443_/D sky130_fd_sc_hd__o211a_1
X_1834_ _1922_/A vssd1 vssd1 vccd1 vccd1 _1834_/X sky130_fd_sc_hd__buf_4
X_1765_ _3302_/Q vssd1 vssd1 vccd1 vccd1 _2106_/B sky130_fd_sc_hd__clkbuf_4
X_3504_ _3512_/CLK _3504_/D vssd1 vssd1 vccd1 vccd1 _3504_/Q sky130_fd_sc_hd__dfxtp_1
X_1696_ _3504_/Q vssd1 vssd1 vccd1 vccd1 _3202_/A sky130_fd_sc_hd__inv_2
X_3435_ _3435_/CLK _3435_/D vssd1 vssd1 vccd1 vccd1 _3435_/Q sky130_fd_sc_hd__dfxtp_1
X_3366_ _3407_/CLK _3366_/D vssd1 vssd1 vccd1 vccd1 _3366_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3297_ _3356_/CLK _3297_/D vssd1 vssd1 vccd1 vccd1 _3297_/Q sky130_fd_sc_hd__dfxtp_1
X_2317_ _3464_/Q _2317_/B vssd1 vssd1 vccd1 vccd1 _2318_/B sky130_fd_sc_hd__xnor2_1
X_2248_ _3383_/Q _2248_/B vssd1 vssd1 vccd1 vccd1 _2254_/B sky130_fd_sc_hd__xnor2_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2103__B1 _2049_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2179_ _3366_/Q vssd1 vssd1 vccd1 vccd1 _2179_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_395 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput67 _3808_/A vssd1 vssd1 vccd1 vccd1 CLR sky130_fd_sc_hd__buf_2
Xoutput78 _3787_/X vssd1 vssd1 vccd1 vccd1 Pd1_b sky130_fd_sc_hd__buf_2
Xoutput89 _3798_/X vssd1 vssd1 vccd1 vccd1 Pd7_a sky130_fd_sc_hd__buf_2
XFILLER_0_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2893__A1 _3447_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2395__B _2395_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input16_A la_data_in[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3220_ _2584_/A _3202_/B _3219_/Y _3213_/X vssd1 vssd1 vccd1 vccd1 _3511_/D sky130_fd_sc_hd__o211a_1
XFILLER_100_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2586__A _2586_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3151_ _3344_/Q _2996_/X _2872_/A _3452_/Q vssd1 vssd1 vccd1 vccd1 _3151_/X sky130_fd_sc_hd__a22o_1
XFILLER_94_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2102_ _2083_/X _2102_/B _2102_/C _2102_/D vssd1 vssd1 vccd1 vccd1 _2102_/X sky130_fd_sc_hd__and4b_1
XFILLER_39_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_15_net107_A clkbuf_2_3__f_net107/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3082_ _3398_/Q _3041_/X _3042_/X _3506_/Q vssd1 vssd1 vccd1 vccd1 _3083_/D sky130_fd_sc_hd__a22o_1
XANTENNA__2636__A1 _3368_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2033_ _2073_/A _2074_/B _2033_/C _2033_/D vssd1 vssd1 vccd1 vccd1 _2048_/A sky130_fd_sc_hd__and4_1
XFILLER_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_148 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2935_ _3461_/Q _2925_/X _2934_/X _2928_/X vssd1 vssd1 vccd1 vccd1 _3461_/D sky130_fd_sc_hd__o211a_1
X_2866_ _2975_/A _2868_/B vssd1 vssd1 vccd1 vccd1 _2866_/X sky130_fd_sc_hd__or2_1
XFILLER_30_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1817_ _3431_/Q _1817_/B vssd1 vssd1 vccd1 vccd1 _1817_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_30_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1665__A _3299_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2797_ _2815_/A vssd1 vssd1 vccd1 vccd1 _2797_/X sky130_fd_sc_hd__clkbuf_2
X_1748_ _1748_/A0 _3534_/Q _1748_/S vssd1 vssd1 vccd1 vccd1 _1749_/A sky130_fd_sc_hd__mux2_2
XFILLER_89_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1679_ _3506_/Q vssd1 vssd1 vccd1 vccd1 _3208_/A sky130_fd_sc_hd__inv_2
X_3418_ _3476_/CLK _3418_/D vssd1 vssd1 vccd1 vccd1 _3418_/Q sky130_fd_sc_hd__dfxtp_1
X_3349_ _3516_/CLK _3349_/D vssd1 vssd1 vccd1 vccd1 _3349_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA_input8_A la_data_in[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_568 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2943__B _3006_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_303 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_88 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3790__A _3790_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3030__A _3199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3043__A1 _3347_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3043__B2 _3431_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2720_ _2758_/A _2726_/B vssd1 vssd1 vccd1 vccd1 _2720_/X sky130_fd_sc_hd__or2_1
XFILLER_12_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2651_ _2762_/A _2653_/B vssd1 vssd1 vccd1 vccd1 _2651_/X sky130_fd_sc_hd__or2_1
XFILLER_8_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_402 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2582_ _2582_/A _2582_/B vssd1 vssd1 vccd1 vccd1 _2582_/X sky130_fd_sc_hd__or2_1
XFILLER_99_479 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3203_ _2565_/A _3191_/X _3202_/Y _3200_/X vssd1 vssd1 vccd1 vccd1 _3504_/D sky130_fd_sc_hd__o211a_1
XANTENNA__1932__B _1932_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3134_ _3427_/Q _2787_/A _3042_/X _3511_/Q vssd1 vssd1 vccd1 vccd1 _3134_/X sky130_fd_sc_hd__a22o_1
XFILLER_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3065_ _3325_/Q _2476_/A _2750_/A _3409_/Q _3064_/X vssd1 vssd1 vccd1 vccd1 _3070_/A
+ sky130_fd_sc_hd__a221o_1
X_2016_ _2016_/A _2016_/B vssd1 vssd1 vccd1 vccd1 _2016_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_35_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3034__B2 _3523_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2918_ _3454_/Q _2910_/X _2917_/X _2915_/X vssd1 vssd1 vccd1 vccd1 _3454_/D sky130_fd_sc_hd__o211a_1
X_2849_ _3432_/Q _2839_/X _2848_/X _2832_/X vssd1 vssd1 vccd1 vccd1 _3432_/D sky130_fd_sc_hd__o211a_1
XFILLER_88_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_462 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3025__B2 _3522_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3785__A _3785_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2703_ _2778_/A _2703_/B vssd1 vssd1 vccd1 vccd1 _2703_/X sky130_fd_sc_hd__or2_1
X_2634_ _2782_/A _2634_/B vssd1 vssd1 vccd1 vccd1 _2634_/X sky130_fd_sc_hd__or2_1
X_2565_ _2565_/A _2568_/B vssd1 vssd1 vccd1 vccd1 _2565_/X sky130_fd_sc_hd__or2_1
XFILLER_99_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1943__A _3314_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_30_net107_A _3436_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2496_ _3326_/Q _2493_/X _2495_/X _2487_/X vssd1 vssd1 vccd1 vccd1 _3326_/D sky130_fd_sc_hd__o211a_1
XFILLER_87_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3117_ _3341_/Q _2996_/X _3037_/A _3461_/Q vssd1 vssd1 vccd1 vccd1 _3117_/X sky130_fd_sc_hd__a22o_1
XFILLER_82_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3255__A1 _3524_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3048_ _3479_/Q _2990_/X _3047_/X _3031_/X vssd1 vssd1 vccd1 vccd1 _3479_/D sky130_fd_sc_hd__o211a_1
XFILLER_23_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2230__A2 _1922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2949__A _3160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2221__A2 _1878_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2859__A _2968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2350_ _2350_/A _2350_/B vssd1 vssd1 vccd1 vccd1 _2351_/B sky130_fd_sc_hd__xnor2_1
XFILLER_69_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2281_ _3469_/Q _2281_/B vssd1 vssd1 vccd1 vccd1 _2333_/A sky130_fd_sc_hd__xnor2_2
XFILLER_77_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2594__A _3227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3237__A1 _3525_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_563 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3804_ _3804_/A vssd1 vssd1 vccd1 vccd1 _3804_/X sky130_fd_sc_hd__clkbuf_1
X_1996_ _1999_/A _1999_/B _1969_/X vssd1 vssd1 vccd1 vccd1 _1998_/A sky130_fd_sc_hd__a21o_1
X_2617_ _3241_/A vssd1 vssd1 vccd1 vccd1 _2771_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__2769__A _2769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2548_ _3343_/Q _2533_/A _2546_/X _2547_/X vssd1 vssd1 vccd1 vccd1 _3343_/D sky130_fd_sc_hd__o211a_1
Xrlbp_macro_218 vssd1 vssd1 vccd1 vccd1 rlbp_macro_218/HI la_data_out[20] sky130_fd_sc_hd__conb_1
Xrlbp_macro_229 vssd1 vssd1 vccd1 vccd1 rlbp_macro_229/HI la_data_out[31] sky130_fd_sc_hd__conb_1
Xrlbp_macro_207 vssd1 vssd1 vccd1 vccd1 rlbp_macro_207/HI la_data_out[9] sky130_fd_sc_hd__conb_1
XFILLER_87_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2479_ _2493_/A vssd1 vssd1 vccd1 vccd1 _2479_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_18_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2436__C1 _2370_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2679__A _2679_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input46_A wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_496 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_135 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1850_ _3425_/Q _2119_/B vssd1 vssd1 vccd1 vccd1 _1851_/B sky130_fd_sc_hd__and2_1
XFILLER_30_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1781_ _3308_/Q vssd1 vssd1 vccd1 vccd1 _2042_/B sky130_fd_sc_hd__clkbuf_4
X_3520_ _3520_/CLK _3520_/D vssd1 vssd1 vccd1 vccd1 _3528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3451_ _3452_/CLK _3451_/D vssd1 vssd1 vccd1 vccd1 _3451_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2589__A _2983_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3382_ _3387_/CLK _3382_/D vssd1 vssd1 vccd1 vccd1 _3382_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2402_ _2405_/B _2405_/C vssd1 vssd1 vccd1 vccd1 _2402_/Y sky130_fd_sc_hd__nand2_1
X_2333_ _2333_/A _2333_/B vssd1 vssd1 vccd1 vccd1 _2334_/B sky130_fd_sc_hd__xor2_1
X_2264_ _2264_/A _2264_/B vssd1 vssd1 vccd1 vccd1 _2265_/B sky130_fd_sc_hd__xnor2_1
XFILLER_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1940__B _3304_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2195_ _3401_/Q _2407_/A vssd1 vssd1 vccd1 vccd1 _2264_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__3213__A _3251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1979_ _2011_/A _2015_/B _1976_/Y _1978_/X vssd1 vssd1 vccd1 vccd1 _1979_/X sky130_fd_sc_hd__a31o_1
XANTENNA__2499__A _2576_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3146__B1 _3195_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_408 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1850__B _2119_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_10_net107 clkbuf_opt_1_0_net107/X vssd1 vssd1 vccd1 vccd1 _3387_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__3793__A _3793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2202__A _3398_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2951_ _2951_/A _2960_/B vssd1 vssd1 vccd1 vccd1 _2951_/X sky130_fd_sc_hd__or2_1
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1902_ _1901_/B _1901_/C _3405_/Q vssd1 vssd1 vccd1 vccd1 _1902_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_15_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2882_ _2895_/A vssd1 vssd1 vccd1 vccd1 _2882_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1833_ _3450_/Q vssd1 vssd1 vccd1 vccd1 _1833_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1764_ _3445_/Q _2105_/B vssd1 vssd1 vccd1 vccd1 _1810_/A sky130_fd_sc_hd__xnor2_1
X_3503_ _3507_/CLK _3503_/D vssd1 vssd1 vccd1 vccd1 _3503_/Q sky130_fd_sc_hd__dfxtp_1
X_1695_ _3510_/Q _2412_/B vssd1 vssd1 vccd1 vccd1 _1695_/X sky130_fd_sc_hd__or2_1
X_3434_ _3435_/CLK _3434_/D vssd1 vssd1 vccd1 vccd1 _3434_/Q sky130_fd_sc_hd__dfxtp_1
X_3365_ _3407_/CLK _3365_/D vssd1 vssd1 vccd1 vccd1 _3365_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3296_ _1748_/A0 _3296_/D vssd1 vssd1 vccd1 vccd1 _3296_/Q sky130_fd_sc_hd__dfxtp_1
X_2316_ _2350_/A _2350_/B _2293_/A vssd1 vssd1 vccd1 vccd1 _2318_/A sky130_fd_sc_hd__a21o_1
X_2247_ _2247_/A _2247_/B vssd1 vssd1 vccd1 vccd1 _2248_/B sky130_fd_sc_hd__xor2_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2178_ _2178_/A _2178_/B _2178_/C _2178_/D vssd1 vssd1 vccd1 vccd1 _2187_/B sky130_fd_sc_hd__and4_1
XFILLER_65_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2782__A _2782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1845__B _2026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput68 _3253_/A2 vssd1 vssd1 vccd1 vccd1 CMP_out_c sky130_fd_sc_hd__buf_2
Xoutput79 _3788_/X vssd1 vssd1 vccd1 vccd1 Pd2_a sky130_fd_sc_hd__buf_2
XFILLER_88_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2957__A _2957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_216 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3788__A _3788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_378 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2581__A1 _3353_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3150_ _3500_/Q _3160_/B _3149_/X vssd1 vssd1 vccd1 vccd1 _3153_/C sky130_fd_sc_hd__a21o_1
XFILLER_94_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_536 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2101_ _2101_/A _2101_/B vssd1 vssd1 vccd1 vccd1 _2102_/D sky130_fd_sc_hd__xnor2_1
X_3081_ _3350_/Q _2554_/A _3021_/X _3434_/Q vssd1 vssd1 vccd1 vccd1 _3083_/C sky130_fd_sc_hd__a22o_1
XFILLER_94_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2032_ _2084_/A _2066_/B vssd1 vssd1 vccd1 vccd1 _2033_/D sky130_fd_sc_hd__and2_1
XFILLER_35_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2934_ _2970_/A _2936_/B vssd1 vssd1 vccd1 vccd1 _2934_/X sky130_fd_sc_hd__or2_1
X_2865_ _3438_/Q _2853_/X _2863_/X _2864_/X vssd1 vssd1 vccd1 vccd1 _3438_/D sky130_fd_sc_hd__o211a_1
XFILLER_30_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1816_ _1816_/A _1816_/B vssd1 vssd1 vccd1 vccd1 _1817_/B sky130_fd_sc_hd__xor2_1
XFILLER_7_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2796_ _2953_/A _2806_/B vssd1 vssd1 vccd1 vccd1 _2796_/X sky130_fd_sc_hd__or2_1
X_1747_ _1747_/A vssd1 vssd1 vccd1 vccd1 _3560_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1678_ _2190_/B vssd1 vssd1 vccd1 vccd1 _1678_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_89_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1681__A _1949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3417_ _3427_/CLK _3417_/D vssd1 vssd1 vccd1 vccd1 _3417_/Q sky130_fd_sc_hd__dfxtp_1
X_3348_ _3516_/CLK _3348_/D vssd1 vssd1 vccd1 vccd1 _3348_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3279_ _2372_/X _2374_/X _2376_/X vssd1 vssd1 vccd1 vccd1 _3279_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_85_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_315 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output115_A _3527_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2650_ _3371_/Q _2642_/X _2649_/X _2635_/X vssd1 vssd1 vccd1 vccd1 _3371_/D sky130_fd_sc_hd__o211a_1
XANTENNA__2024__A_N _1949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1766__A _3446_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2581_ _3353_/Q _2570_/X _2578_/X _2580_/X vssd1 vssd1 vccd1 vccd1 _3353_/D sky130_fd_sc_hd__o211a_1
XFILLER_99_414 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2597__A _2756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3202_ _3202_/A _3202_/B vssd1 vssd1 vccd1 vccd1 _3202_/Y sky130_fd_sc_hd__nand2_1
XFILLER_79_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3133_ _3486_/Q _3074_/X _3132_/X _3098_/X vssd1 vssd1 vccd1 vccd1 _3486_/D sky130_fd_sc_hd__o211a_1
X_3064_ _3445_/Q _2872_/A _3008_/A _3493_/Q vssd1 vssd1 vccd1 vccd1 _3064_/X sky130_fd_sc_hd__a22o_1
X_2015_ _3328_/Q _2015_/B vssd1 vssd1 vccd1 vccd1 _2016_/B sky130_fd_sc_hd__xnor2_1
XFILLER_63_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3034__A2 _2679_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2917_ _2953_/A _2923_/B vssd1 vssd1 vccd1 vccd1 _2917_/X sky130_fd_sc_hd__or2_1
XFILLER_12_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_48 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2848_ _2957_/A _2850_/B vssd1 vssd1 vccd1 vccd1 _2848_/X sky130_fd_sc_hd__or2_1
XANTENNA__2545__A1 _3342_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2779_ _3414_/Q _2767_/X _2778_/X _2776_/X vssd1 vssd1 vccd1 vccd1 _3414_/D sky130_fd_sc_hd__o211a_1
XFILLER_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2047__A_N _3549_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2970__A _2970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_380 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_428 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2702_ _3389_/Q _2692_/X _2701_/X _2699_/X vssd1 vssd1 vccd1 vccd1 _3389_/D sky130_fd_sc_hd__o211a_1
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2633_ _3188_/A vssd1 vssd1 vccd1 vccd1 _2782_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_99_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2564_ _3347_/Q _2556_/X _2563_/X _2547_/X vssd1 vssd1 vccd1 vccd1 _3347_/D sky130_fd_sc_hd__o211a_1
XFILLER_99_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2495_ _2572_/A _2505_/B vssd1 vssd1 vccd1 vccd1 _2495_/X sky130_fd_sc_hd__or2_1
XFILLER_101_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3116_ _3413_/Q _2751_/A _3115_/X vssd1 vssd1 vccd1 vccd1 _3119_/B sky130_fd_sc_hd__a21o_1
XFILLER_55_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3047_ _3311_/Q _2988_/X _3012_/A _3046_/X vssd1 vssd1 vccd1 vccd1 _3047_/X sky130_fd_sc_hd__a211o_1
XANTENNA__2790__A _3227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2766__A1 _3409_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3796__A input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_64 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2757__A1 _3405_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2205__A _3400_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3182__A1 _3497_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2280_ _2280_/A _2329_/A _2330_/B _2280_/D vssd1 vssd1 vccd1 vccd1 _2297_/A sky130_fd_sc_hd__and4_1
XFILLER_36_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2875__A _2875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_2_0__f_net107 clkbuf_0_net107/X vssd1 vssd1 vccd1 vccd1 _3494_/CLK sky130_fd_sc_hd__clkbuf_16
X_3803_ _3803_/A vssd1 vssd1 vccd1 vccd1 _3803_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_575 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1995_ _3321_/Q _1995_/B _1995_/C vssd1 vssd1 vccd1 vccd1 _1995_/X sky130_fd_sc_hd__or3_1
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2616_ _3362_/Q _2612_/X _2615_/X _2601_/X vssd1 vssd1 vccd1 vccd1 _3362_/D sky130_fd_sc_hd__o211a_1
XANTENNA__1971__A2 _1878_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2547_ _2566_/A vssd1 vssd1 vccd1 vccd1 _2547_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xrlbp_macro_219 vssd1 vssd1 vccd1 vccd1 rlbp_macro_219/HI la_data_out[21] sky130_fd_sc_hd__conb_1
Xrlbp_macro_208 vssd1 vssd1 vccd1 vccd1 rlbp_macro_208/HI la_data_out[10] sky130_fd_sc_hd__conb_1
XFILLER_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2920__A1 _3455_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2478_ _3223_/A _2480_/B vssd1 vssd1 vccd1 vccd1 _2493_/A sky130_fd_sc_hd__and2_1
XFILLER_87_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2025__A _3347_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2679__B _2679_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input39_A wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_33_net107 _3494_/CLK vssd1 vssd1 vccd1 vccd1 _3445_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_75_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_30 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1758__B _2119_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1780_ _1780_/A _1780_/B vssd1 vssd1 vccd1 vccd1 _1837_/A sky130_fd_sc_hd__nor2_1
XFILLER_30_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3450_ _3450_/CLK _3450_/D vssd1 vssd1 vccd1 vccd1 _3450_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2589__B _2709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3381_ _3396_/CLK _3381_/D vssd1 vssd1 vccd1 vccd1 _3381_/Q sky130_fd_sc_hd__dfxtp_1
X_2401_ _2399_/A _2399_/B _2400_/Y _2397_/X vssd1 vssd1 vccd1 vccd1 _3302_/D sky130_fd_sc_hd__o211a_1
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2902__A1 _3451_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2332_ _3454_/Q _2329_/Y _2330_/X _2331_/Y vssd1 vssd1 vccd1 vccd1 _2332_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2263_ _2262_/A _2262_/B _2262_/C vssd1 vssd1 vccd1 vccd1 _2263_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_84_228 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2194_ _1949_/A _3393_/Q vssd1 vssd1 vccd1 vccd1 _2251_/B sky130_fd_sc_hd__nand2b_2
XFILLER_65_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1949__A _1949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2108__A_N _2309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1978_ _1938_/A _1977_/X _1941_/B vssd1 vssd1 vccd1 vccd1 _1978_/X sky130_fd_sc_hd__a21o_1
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3137__A1 _3355_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_431 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_604 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2950_ _2977_/B vssd1 vssd1 vccd1 vccd1 _2960_/B sky130_fd_sc_hd__clkbuf_1
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1901_ _3405_/Q _1901_/B _1901_/C vssd1 vssd1 vccd1 vccd1 _1901_/X sky130_fd_sc_hd__and3_1
X_2881_ _2955_/A _2886_/B vssd1 vssd1 vccd1 vccd1 _2881_/X sky130_fd_sc_hd__or2_1
X_1832_ _1832_/A _1832_/B _1832_/C _1832_/D vssd1 vssd1 vccd1 vccd1 _1842_/B sky130_fd_sc_hd__and4_1
X_1763_ _3301_/Q vssd1 vssd1 vccd1 vccd1 _2105_/B sky130_fd_sc_hd__buf_4
X_3502_ _3512_/CLK _3502_/D vssd1 vssd1 vccd1 vccd1 _3502_/Q sky130_fd_sc_hd__dfxtp_1
X_1694_ _3510_/Q _2412_/B vssd1 vssd1 vccd1 vccd1 _1694_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__2112__B _2206_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3433_ _3440_/CLK _3433_/D vssd1 vssd1 vccd1 vccd1 _3433_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__3128__A1 _3474_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3128__B2 _3498_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3364_ _3407_/CLK _3364_/D vssd1 vssd1 vccd1 vccd1 _3364_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1951__B _3299_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3295_ _3295_/D _2356_/X vssd1 vssd1 vccd1 vccd1 _3295_/Q sky130_fd_sc_hd__dlxtn_2
X_2315_ _2299_/Y _1693_/A _2280_/A _2339_/B _2314_/X vssd1 vssd1 vccd1 vccd1 _2350_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_85_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2246_ _2246_/A _2246_/B vssd1 vssd1 vccd1 vccd1 _2254_/A sky130_fd_sc_hd__xnor2_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2103__A2 _2102_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2177_ _3375_/Q _2177_/B vssd1 vssd1 vccd1 vccd1 _2178_/D sky130_fd_sc_hd__or2_1
XFILLER_38_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput69 _3778_/X vssd1 vssd1 vccd1 vccd1 OTA_out_c sky130_fd_sc_hd__buf_2
XFILLER_88_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2973__A _2973_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_272 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3055__B1 _2643_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_320 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1771__B _2309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_548 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2100_ _3344_/Q _2100_/B vssd1 vssd1 vccd1 vccd1 _2101_/B sky130_fd_sc_hd__xnor2_1
X_3080_ _3326_/Q _2476_/A _2750_/A _3410_/Q _3079_/X vssd1 vssd1 vccd1 vccd1 _3083_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_94_367 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2031_ _3354_/Q _2121_/B vssd1 vssd1 vccd1 vccd1 _2066_/B sky130_fd_sc_hd__xnor2_1
XFILLER_35_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_434 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3046__B1 _3035_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2933_ _3460_/Q _2925_/X _2932_/X _2928_/X vssd1 vssd1 vccd1 vccd1 _3460_/D sky130_fd_sc_hd__o211a_1
XFILLER_50_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2864_ _2895_/A vssd1 vssd1 vccd1 vccd1 _2864_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_clkbuf_leaf_24_net107_A _3436_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1815_ _3430_/Q _1812_/Y _1813_/X _1814_/Y vssd1 vssd1 vccd1 vccd1 _1815_/Y sky130_fd_sc_hd__a211oi_1
X_2795_ _3230_/A vssd1 vssd1 vccd1 vccd1 _2953_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__2123__A _3358_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1746_ _3563_/Q _3564_/Q vssd1 vssd1 vccd1 vccd1 _1747_/A sky130_fd_sc_hd__and2b_1
XFILLER_7_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1940__A_N _3316_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1677_ _3299_/Q vssd1 vssd1 vccd1 vccd1 _2190_/B sky130_fd_sc_hd__clkbuf_4
X_3416_ _3427_/CLK _3416_/D vssd1 vssd1 vccd1 vccd1 _3416_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3347_ _3516_/CLK _3347_/D vssd1 vssd1 vccd1 vccd1 _3347_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3278_ _2372_/X _2374_/X _2376_/X vssd1 vssd1 vccd1 vccd1 _3278_/Y sky130_fd_sc_hd__a21oi_2
X_2229_ _3401_/Q _2313_/B vssd1 vssd1 vccd1 vccd1 _2229_/Y sky130_fd_sc_hd__nor2_1
XFILLER_66_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2793__A _2951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1856__B _2106_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2968__A _2968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2315__A2 _1693_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3799__A input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input21_A la_data_in[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3028__B1 _3016_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1766__B _2106_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2580_ _2654_/A vssd1 vssd1 vccd1 vccd1 _2580_/X sky130_fd_sc_hd__buf_2
XFILLER_99_426 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3201_ _2563_/A _3191_/X _3198_/Y _3200_/X vssd1 vssd1 vccd1 vccd1 _3503_/D sky130_fd_sc_hd__o211a_1
XFILLER_79_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3132_ _3155_/A _3132_/B vssd1 vssd1 vccd1 vccd1 _3132_/X sky130_fd_sc_hd__or2_1
XFILLER_94_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3063_ _3421_/Q _2791_/B _2949_/B _3469_/Q _3062_/X vssd1 vssd1 vccd1 vccd1 _3063_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_94_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2014_ _2011_/A _2011_/B _1938_/A vssd1 vssd1 vccd1 vccd1 _2016_/A sky130_fd_sc_hd__a21o_1
XFILLER_35_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2118__A _3365_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2490__A1 _3324_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2916_ _3453_/Q _2910_/X _2913_/X _2915_/X vssd1 vssd1 vccd1 vccd1 _3453_/D sky130_fd_sc_hd__o211a_1
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2847_ _3431_/Q _2839_/X _2846_/X _2832_/X vssd1 vssd1 vccd1 vccd1 _3431_/D sky130_fd_sc_hd__o211a_1
X_2778_ _2778_/A _2778_/B vssd1 vssd1 vccd1 vccd1 _2778_/X sky130_fd_sc_hd__or2_1
X_1729_ _1729_/A vssd1 vssd1 vccd1 vccd1 _3808_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__2788__A _2788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2028__A _3353_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1867__A _1932_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2698__A _2773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1777__A _3451_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2701_ _2775_/A _2703_/B vssd1 vssd1 vccd1 vccd1 _2701_/X sky130_fd_sc_hd__or2_1
X_2632_ _3367_/Q _2612_/A _2631_/X _2619_/X vssd1 vssd1 vccd1 vccd1 _3367_/D sky130_fd_sc_hd__o211a_1
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2563_ _2563_/A _2568_/B vssd1 vssd1 vccd1 vccd1 _2563_/X sky130_fd_sc_hd__or2_1
X_2494_ _2509_/B vssd1 vssd1 vccd1 vccd1 _2505_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_95_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3115_ _3425_/Q _2985_/B _3056_/A _3509_/Q vssd1 vssd1 vccd1 vccd1 _3115_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3232__A _3232_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3046_ _3419_/Q _2791_/B _3035_/X _3045_/X vssd1 vssd1 vccd1 vccd1 _3046_/X sky130_fd_sc_hd__a211o_1
XFILLER_82_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1726__B1 _1667_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_407 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2205__B _2285_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3167__C1 _3156_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2445__A1 _3313_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3802_ _3802_/A vssd1 vssd1 vccd1 vccd1 _3802_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_60_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_587 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_395 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1994_ _1995_/B _1995_/C _3321_/Q vssd1 vssd1 vccd1 vccd1 _1994_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_20_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2115__B _2115_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2615_ _2769_/A _2628_/B vssd1 vssd1 vccd1 vccd1 _2615_/X sky130_fd_sc_hd__or2_1
XANTENNA__1954__B _2118_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3227__A _3227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2546_ _2584_/A _2549_/B vssd1 vssd1 vccd1 vccd1 _2546_/X sky130_fd_sc_hd__or2_1
Xrlbp_macro_209 vssd1 vssd1 vccd1 vccd1 rlbp_macro_209/HI la_data_out[11] sky130_fd_sc_hd__conb_1
X_2477_ _2477_/A vssd1 vssd1 vccd1 vccd1 _2480_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_68_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_156 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3029_ _3121_/A _3029_/B vssd1 vssd1 vccd1 vccd1 _3029_/X sky130_fd_sc_hd__or2_1
XFILLER_24_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2025__B _2025_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_99 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_42 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2216__A _3396_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1774__B _1774_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2400_ _2405_/C vssd1 vssd1 vccd1 vccd1 _2400_/Y sky130_fd_sc_hd__inv_2
X_3380_ _3392_/CLK _3380_/D vssd1 vssd1 vccd1 vccd1 _3380_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2886__A _2960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2331_ _2330_/B _2330_/C _3453_/Q vssd1 vssd1 vccd1 vccd1 _2331_/Y sky130_fd_sc_hd__a21oi_1
X_2262_ _2262_/A _2262_/B _2262_/C vssd1 vssd1 vccd1 vccd1 _2262_/X sky130_fd_sc_hd__or3_1
XFILLER_2_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2193_ _3394_/Q _3298_/Q vssd1 vssd1 vccd1 vccd1 _2249_/A sky130_fd_sc_hd__xnor2_1
XFILLER_1_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3091__A1 _3447_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2126__A _3368_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1977_ _2285_/B _3316_/Q vssd1 vssd1 vccd1 vccd1 _1977_/X sky130_fd_sc_hd__or2b_1
XANTENNA_clkbuf_leaf_1_net107_A _3494_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3146__A2 _2557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2529_ _2565_/A _2531_/B vssd1 vssd1 vccd1 vccd1 _2529_/X sky130_fd_sc_hd__or2_1
XANTENNA__2796__A _2953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2409__A1 _2407_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1859__B _2309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3082__A1 _3398_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input51_A wbs_cyc_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2896__A1 _3448_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2648__A1 _3370_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1769__B _3448_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_6 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1900_ _1900_/A _1901_/B vssd1 vssd1 vccd1 vccd1 _1900_/Y sky130_fd_sc_hd__xnor2_1
X_2880_ _3442_/Q _2874_/X _2879_/X _2864_/X vssd1 vssd1 vccd1 vccd1 _3442_/D sky130_fd_sc_hd__o211a_1
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1831_ _1831_/A _1831_/B vssd1 vssd1 vccd1 vccd1 _1832_/D sky130_fd_sc_hd__xnor2_1
XFILLER_42_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1762_ _1762_/A _1812_/A _1813_/B _1762_/D vssd1 vssd1 vccd1 vccd1 _1785_/A sky130_fd_sc_hd__and4_1
X_1693_ _1693_/A vssd1 vssd1 vccd1 vccd1 _2412_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3501_ _3512_/CLK _3501_/D vssd1 vssd1 vccd1 vccd1 _3501_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3432_ _3440_/CLK _3432_/D vssd1 vssd1 vccd1 vccd1 _3432_/Q sky130_fd_sc_hd__dfxtp_1
X_3363_ _3414_/CLK _3363_/D vssd1 vssd1 vccd1 vccd1 _3363_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2887__A1 _3445_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3294_ _3464_/CLK _3294_/D _2377_/Y vssd1 vssd1 vccd1 vccd1 _3294_/Q sky130_fd_sc_hd__dfrtp_1
X_2314_ _2299_/Y _1922_/X _2313_/Y vssd1 vssd1 vccd1 vccd1 _2314_/X sky130_fd_sc_hd__o21a_1
X_2245_ _3384_/Q _2245_/B vssd1 vssd1 vccd1 vccd1 _2246_/B sky130_fd_sc_hd__xor2_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2176_ _3375_/Q _2177_/B vssd1 vssd1 vccd1 vccd1 _2178_/C sky130_fd_sc_hd__nand2_1
XFILLER_38_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3064__A1 _3445_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1695__A _3510_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3055__B2 _3372_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_387 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2869__A1 _3440_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2030_ _2030_/A _2030_/B vssd1 vssd1 vccd1 vccd1 _2084_/A sky130_fd_sc_hd__nor2_1
XFILLER_11_6 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_379 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_427 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2932_ _2968_/A _2936_/B vssd1 vssd1 vccd1 vccd1 _2932_/X sky130_fd_sc_hd__or2_1
X_2863_ _2973_/A _2863_/B vssd1 vssd1 vccd1 vccd1 _2863_/X sky130_fd_sc_hd__or2_1
X_1814_ _1813_/B _1813_/C _3429_/Q vssd1 vssd1 vccd1 vccd1 _1814_/Y sky130_fd_sc_hd__a21oi_1
X_2794_ _3417_/Q _2789_/X _2793_/X _2776_/X vssd1 vssd1 vccd1 vccd1 _3417_/D sky130_fd_sc_hd__o211a_1
X_1745_ _1745_/A vssd1 vssd1 vccd1 vccd1 _3555_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2123__B _2389_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_380 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1676_ _3505_/Q vssd1 vssd1 vccd1 vccd1 _3205_/A sky130_fd_sc_hd__inv_2
X_3415_ _3427_/CLK _3415_/D vssd1 vssd1 vccd1 vccd1 _3415_/Q sky130_fd_sc_hd__dfxtp_1
X_3346_ _3516_/CLK _3346_/D vssd1 vssd1 vccd1 vccd1 _3346_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_302 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3277_ _2372_/X _2374_/X _2376_/X vssd1 vssd1 vccd1 vccd1 _3277_/Y sky130_fd_sc_hd__a21oi_2
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2228_ _2212_/A _2212_/B _2235_/B _2227_/X vssd1 vssd1 vccd1 vccd1 _2264_/B sky130_fd_sc_hd__a31o_1
XFILLER_26_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2159_ _3372_/Q _2159_/B vssd1 vssd1 vccd1 vccd1 _2160_/B sky130_fd_sc_hd__xnor2_1
XFILLER_81_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1835__A2 _1693_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input14_A la_data_in[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3028__A1 _3310_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2208__B _2291_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1782__B _2042_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3200_ _3251_/A vssd1 vssd1 vccd1 vccd1 _3200_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3131_ _3318_/Q _2988_/A _3124_/X _3130_/X vssd1 vssd1 vccd1 vccd1 _3132_/B sky130_fd_sc_hd__a211o_1
XANTENNA__2894__A _2968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3062_ _3361_/Q _3036_/X _3037_/X _3457_/Q vssd1 vssd1 vccd1 vccd1 _3062_/X sky130_fd_sc_hd__a22o_1
X_2013_ _3327_/Q _2013_/B vssd1 vssd1 vccd1 vccd1 _2013_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__3019__A1 _3322_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2118__B _2118_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3019__B2 _3406_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2915_ _2971_/A vssd1 vssd1 vccd1 vccd1 _2915_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__1957__B _2121_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2846_ _2955_/A _2850_/B vssd1 vssd1 vccd1 vccd1 _2846_/X sky130_fd_sc_hd__or2_1
X_2777_ _3413_/Q _2767_/X _2775_/X _2776_/X vssd1 vssd1 vccd1 vccd1 _3413_/D sky130_fd_sc_hd__o211a_1
XANTENNA__1973__A _3314_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1728_ _1719_/X _1728_/B _1728_/C _1728_/D vssd1 vssd1 vccd1 vccd1 _1729_/A sky130_fd_sc_hd__and4b_1
X_1659_ _2285_/B vssd1 vssd1 vccd1 vccd1 _2037_/B sky130_fd_sc_hd__buf_2
XANTENNA_input6_A la_data_in[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3329_ _3332_/CLK _3329_/D vssd1 vssd1 vccd1 vccd1 _3329_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2309__A _2309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2028__B _2313_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2044__A _3355_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_16_net107 clkbuf_2_3__f_net107/X vssd1 vssd1 vccd1 vccd1 _3377_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_76_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2219__A _3395_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1777__B _2115_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2700_ _3388_/Q _2692_/X _2698_/X _2699_/X vssd1 vssd1 vccd1 vccd1 _3388_/D sky130_fd_sc_hd__o211a_1
XFILLER_13_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2631_ _2780_/A _2634_/B vssd1 vssd1 vccd1 vccd1 _2631_/X sky130_fd_sc_hd__or2_1
XFILLER_9_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2562_ _3346_/Q _2556_/X _2561_/X _2547_/X vssd1 vssd1 vccd1 vccd1 _3346_/D sky130_fd_sc_hd__o211a_1
XFILLER_57_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2493_ _2493_/A vssd1 vssd1 vccd1 vccd1 _2493_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_99_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3114_ _3365_/Q _3036_/A _3018_/X _3497_/Q _3113_/X vssd1 vssd1 vccd1 vccd1 _3119_/A
+ sky130_fd_sc_hd__a221o_1
X_3045_ _3467_/Q _2946_/A _3038_/X _3040_/X _3044_/X vssd1 vssd1 vccd1 vccd1 _3045_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_36_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2799__A _3232_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2829_ _3188_/A vssd1 vssd1 vccd1 vccd1 _2977_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_2_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_240 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2439__C1 _2370_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1878__A _2191_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1662__B1 _1657_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_463 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_3_net107 clkbuf_leaf_9_net107/A vssd1 vssd1 vccd1 vccd1 _3307_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_6_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1717__B2 _3489_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1717__A1 _3492_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2390__A1 _1667_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_2_3__f_net107_A clkbuf_0_net107/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3801_ _3801_/A vssd1 vssd1 vccd1 vccd1 _3801_/X sky130_fd_sc_hd__clkbuf_1
X_1993_ _2001_/B vssd1 vssd1 vccd1 vccd1 _1995_/B sky130_fd_sc_hd__inv_2
XFILLER_33_599 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2614_ _2634_/B vssd1 vssd1 vccd1 vccd1 _2628_/B sky130_fd_sc_hd__clkbuf_1
X_2545_ _3342_/Q _2533_/X _2544_/X _2536_/X vssd1 vssd1 vccd1 vccd1 _3342_/D sky130_fd_sc_hd__o211a_1
XFILLER_87_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2476_ _2476_/A vssd1 vssd1 vccd1 vccd1 _2477_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3243__A _3243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_496 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3028_ _3310_/Q _2993_/X _3016_/X _3027_/X vssd1 vssd1 vccd1 vccd1 _3029_/B sky130_fd_sc_hd__a211o_1
XFILLER_70_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1698__A _1698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_363 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3153__A _3153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_6 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2330_ _3453_/Q _2330_/B _2330_/C vssd1 vssd1 vccd1 vccd1 _2330_/X sky130_fd_sc_hd__and3_1
X_2261_ _3388_/Q _2261_/B vssd1 vssd1 vccd1 vccd1 _2262_/C sky130_fd_sc_hd__xnor2_1
XFILLER_69_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2192_ _2247_/A _2245_/B vssd1 vssd1 vccd1 vccd1 _2213_/A sky130_fd_sc_hd__nor2_1
XFILLER_77_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_18_net107_A clkbuf_2_3__f_net107/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2407__A _2407_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2126__B _2294_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1976_ _1972_/X _1973_/X _1975_/X vssd1 vssd1 vccd1 vccd1 _1976_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__3238__A _3238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2142__A _3362_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2528_ _3335_/Q _2518_/X _2527_/X _2523_/X vssd1 vssd1 vccd1 vccd1 _3335_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2459_ _3317_/Q _2446_/X _2458_/X _2444_/X vssd1 vssd1 vccd1 vccd1 _3317_/D sky130_fd_sc_hd__o211a_1
XFILLER_68_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2317__A _3464_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3082__A2 _3041_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input44_A wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1830_ _3436_/Q _1830_/B vssd1 vssd1 vccd1 vccd1 _1831_/B sky130_fd_sc_hd__xnor2_1
XFILLER_30_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1761_ _1827_/A _1805_/B vssd1 vssd1 vccd1 vccd1 _1762_/D sky130_fd_sc_hd__and2_1
X_3500_ _3507_/CLK _3500_/D vssd1 vssd1 vccd1 vccd1 _3500_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1692_ _1922_/A vssd1 vssd1 vccd1 vccd1 _1693_/A sky130_fd_sc_hd__buf_4
X_3431_ _3440_/CLK _3431_/D vssd1 vssd1 vccd1 vccd1 _3431_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__2897__A _2970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3362_ _3407_/CLK _3362_/D vssd1 vssd1 vccd1 vccd1 _3362_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2313_ _3473_/Q _2313_/B vssd1 vssd1 vccd1 vccd1 _2313_/Y sky130_fd_sc_hd__nor2_1
XFILLER_85_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3293_ _3436_/CLK _3293_/D _2370_/X vssd1 vssd1 vccd1 vccd1 _3293_/Q sky130_fd_sc_hd__dfrtp_1
X_2244_ _2219_/Y _1667_/X _2243_/X vssd1 vssd1 vccd1 vccd1 _2246_/A sky130_fd_sc_hd__a21o_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2175_ _2175_/A _2175_/B vssd1 vssd1 vccd1 vccd1 _2177_/B sky130_fd_sc_hd__xnor2_1
XFILLER_38_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_127 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2575__A1 _3351_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1959_ _1959_/A _1959_/B vssd1 vssd1 vccd1 vccd1 _1962_/B sky130_fd_sc_hd__nand2_1
XANTENNA__2600__A _2758_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_399 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_255 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2931_ _3459_/Q _2925_/X _2930_/X _2928_/X vssd1 vssd1 vccd1 vccd1 _3459_/D sky130_fd_sc_hd__o211a_1
XANTENNA__1796__A _2282_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2862_ _3437_/Q _2853_/X _2861_/X _2851_/X vssd1 vssd1 vccd1 vccd1 _3437_/D sky130_fd_sc_hd__o211a_1
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1813_ _3429_/Q _1813_/B _1813_/C vssd1 vssd1 vccd1 vccd1 _1813_/X sky130_fd_sc_hd__and3_1
X_2793_ _2951_/A _2806_/B vssd1 vssd1 vccd1 vccd1 _2793_/X sky130_fd_sc_hd__or2_1
X_1744_ _3559_/Q _2189_/B vssd1 vssd1 vccd1 vccd1 _1745_/A sky130_fd_sc_hd__and2_1
X_3414_ _3414_/CLK _3414_/D vssd1 vssd1 vccd1 vccd1 _3414_/Q sky130_fd_sc_hd__dfxtp_1
X_1675_ _3509_/Q _2313_/B _1667_/X _3198_/A _1674_/X vssd1 vssd1 vccd1 vccd1 _1686_/C
+ sky130_fd_sc_hd__a221o_1
X_3345_ _3516_/CLK _3345_/D vssd1 vssd1 vccd1 vccd1 _3345_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3276_ _2372_/X _2374_/X _2376_/X vssd1 vssd1 vccd1 vccd1 _3276_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA_clkbuf_leaf_33_net107_A _3494_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2227_ _2222_/Y _2037_/B _2212_/B _2224_/Y _2226_/X vssd1 vssd1 vccd1 vccd1 _2227_/X
+ sky130_fd_sc_hd__a221o_1
Xrepeater132 _3807_/A vssd1 vssd1 vccd1 vccd1 _3253_/A2 sky130_fd_sc_hd__buf_2
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3251__A _3251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2158_ _3359_/Q _1678_/Y _2157_/Y vssd1 vssd1 vccd1 vccd1 _2160_/A sky130_fd_sc_hd__o21ai_1
XFILLER_81_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2089_ _3339_/Q _2089_/B vssd1 vssd1 vccd1 vccd1 _2093_/C sky130_fd_sc_hd__nand2_1
XFILLER_81_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2548__A1 _3343_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2330__A _3453_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2505__A _2582_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2539__A1 _3339_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_39_net107 _3494_/CLK vssd1 vssd1 vccd1 vccd1 _3491_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_output75_A _3784_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3130_ _3414_/Q _2754_/B _3125_/X _3127_/X _3129_/X vssd1 vssd1 vccd1 vccd1 _3130_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_94_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrlbp_macro_190 vssd1 vssd1 vccd1 vccd1 rlbp_macro_190/HI io_out[33] sky130_fd_sc_hd__conb_1
XFILLER_67_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3061_ _3480_/Q _2990_/X _3060_/X _3031_/X vssd1 vssd1 vccd1 vccd1 _3480_/D sky130_fd_sc_hd__o211a_1
XFILLER_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2012_ _3327_/Q _2013_/B vssd1 vssd1 vccd1 vccd1 _2012_/X sky130_fd_sc_hd__or2_1
XFILLER_63_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2914_ _3199_/A vssd1 vssd1 vccd1 vccd1 _2971_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2845_ _3430_/Q _2839_/X _2844_/X _2832_/X vssd1 vssd1 vccd1 vccd1 _3430_/D sky130_fd_sc_hd__o211a_1
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2776_ _2815_/A vssd1 vssd1 vccd1 vccd1 _2776_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3246__A _3262_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1727_ _3494_/Q _1673_/Y _1724_/X _1725_/Y _1726_/X vssd1 vssd1 vccd1 vccd1 _1728_/D
+ sky130_fd_sc_hd__o221a_1
XANTENNA__2150__A _3378_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1658_ _3304_/Q vssd1 vssd1 vccd1 vccd1 _2285_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__2702__A1 _3389_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3328_ _3332_/CLK _3328_/D vssd1 vssd1 vccd1 vccd1 _3328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3259_ _3526_/Q _1707_/A _3251_/X _3258_/X vssd1 vssd1 vccd1 vccd1 _3526_/D sky130_fd_sc_hd__o211a_1
XFILLER_37_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2044__B _2115_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3194__A1 _2559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2060__A _3350_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_2_2__f_net107_A clkbuf_0_net107/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output113_A _3525_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2630_ _3186_/A vssd1 vssd1 vccd1 vccd1 _2780_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__3185__A1 _3498_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2561_ _2561_/A _2568_/B vssd1 vssd1 vccd1 vccd1 _2561_/X sky130_fd_sc_hd__or2_1
XFILLER_99_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2492_ _3325_/Q _2479_/X _2491_/X _2487_/X vssd1 vssd1 vccd1 vccd1 _3325_/D sky130_fd_sc_hd__o211a_1
XFILLER_4_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1755__A_N _2389_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3113_ _3389_/Q _3053_/X _2944_/A _3473_/Q vssd1 vssd1 vccd1 vccd1 _3113_/X sky130_fd_sc_hd__a22o_1
XFILLER_95_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3044_ _3395_/Q _3041_/X _3042_/X _3503_/Q _3043_/X vssd1 vssd1 vccd1 vccd1 _3044_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_82_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2999__B2 _3369_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_236 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2145__A _2145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1984__A _3331_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2828_ _3427_/Q _2808_/A _2827_/X _2815_/X vssd1 vssd1 vccd1 vccd1 _3427_/D sky130_fd_sc_hd__o211a_1
X_2759_ _3406_/Q _2753_/X _2758_/X _2743_/X vssd1 vssd1 vccd1 vccd1 _3406_/D sky130_fd_sc_hd__o211a_1
XFILLER_2_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_22_net107 _3436_/CLK vssd1 vssd1 vccd1 vccd1 _3476_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_98_291 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2039__B _2288_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3100__A1 _3448_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3100__B2 _3496_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1662__A1 _3511_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3167__A1 _3491_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1717__A2 _1657_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3800_ _3800_/A vssd1 vssd1 vccd1 vccd1 _3800_/X sky130_fd_sc_hd__clkbuf_1
X_1992_ _1992_/A _1992_/B vssd1 vssd1 vccd1 vccd1 _2006_/C sky130_fd_sc_hd__xnor2_1
X_2613_ _3238_/A vssd1 vssd1 vccd1 vccd1 _2769_/A sky130_fd_sc_hd__clkbuf_2
X_2544_ _2582_/A _2544_/B vssd1 vssd1 vccd1 vccd1 _2544_/X sky130_fd_sc_hd__or2_1
XFILLER_87_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2475_ _2981_/A vssd1 vssd1 vccd1 vccd1 _2476_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_95_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3027_ _3027_/A _3027_/B _3027_/C _3027_/D vssd1 vssd1 vccd1 vccd1 _3027_/X sky130_fd_sc_hd__or4_1
XFILLER_63_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_375 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2603__A _3232_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3149__B2 _3464_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3149__A1 _3368_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2260_ _2260_/A _2260_/B vssd1 vssd1 vccd1 vccd1 _2262_/B sky130_fd_sc_hd__nor2_1
XFILLER_2_460 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2191_ _3396_/Q _2191_/B vssd1 vssd1 vccd1 vccd1 _2245_/B sky130_fd_sc_hd__xor2_1
XFILLER_77_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1975_ _1974_/X _3314_/Q vssd1 vssd1 vccd1 vccd1 _1975_/X sky130_fd_sc_hd__and2b_1
XANTENNA__2587__C1 _2580_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2527_ _2563_/A _2531_/B vssd1 vssd1 vccd1 vccd1 _2527_/X sky130_fd_sc_hd__or2_1
XANTENNA__3254__A _3523_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2458_ _2578_/A _2461_/B vssd1 vssd1 vccd1 vccd1 _2458_/X sky130_fd_sc_hd__or2_1
XFILLER_96_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2389_ _2389_/A _2389_/B _2389_/C hold5/A vssd1 vssd1 vccd1 vccd1 _2395_/C sky130_fd_sc_hd__and4_1
XFILLER_29_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2052__B _2052_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3164__A _3230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input37_A la_data_in[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3058__B1 _3195_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1760_ _3450_/Q _1922_/A vssd1 vssd1 vccd1 vccd1 _1805_/B sky130_fd_sc_hd__xnor2_1
XFILLER_7_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1691_ _3306_/Q vssd1 vssd1 vccd1 vccd1 _1922_/A sky130_fd_sc_hd__clkbuf_2
X_3430_ _3440_/CLK _3430_/D vssd1 vssd1 vccd1 vccd1 _3430_/Q sky130_fd_sc_hd__dfxtp_2
X_3361_ _3377_/CLK _3361_/D vssd1 vssd1 vccd1 vccd1 _3361_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2312_ _2296_/A _2333_/B _2311_/X vssd1 vssd1 vccd1 vccd1 _2339_/B sky130_fd_sc_hd__a21o_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3292_ _3292_/D _2356_/X vssd1 vssd1 vccd1 vccd1 _3294_/D sky130_fd_sc_hd__dlxtn_1
XANTENNA__3802__A _3802_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2243_ _2247_/A _2247_/B vssd1 vssd1 vccd1 vccd1 _2243_/X sky130_fd_sc_hd__and2b_1
XFILLER_78_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2174_ _2174_/A _2174_/B vssd1 vssd1 vccd1 vccd1 _2178_/B sky130_fd_sc_hd__xnor2_1
XFILLER_38_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_139 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_278 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3249__A _3521_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2153__A _3374_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1958_ _2007_/A _1986_/B vssd1 vssd1 vccd1 vccd1 _1959_/B sky130_fd_sc_hd__and2_1
X_1889_ _1888_/X _1864_/B _1860_/B vssd1 vssd1 vccd1 vccd1 _1889_/X sky130_fd_sc_hd__a21o_1
XFILLER_88_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3559_ _3559_/CLK _3559_/D _3288_/Y vssd1 vssd1 vccd1 vccd1 _3559_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_88_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3288__B1 _3282_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2047__B _3548_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_492 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_599 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_540 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3543__RESET_B _3278_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2930_ _2966_/A _2936_/B vssd1 vssd1 vccd1 vccd1 _2930_/X sky130_fd_sc_hd__or2_1
XFILLER_15_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2861_ _2970_/A _2863_/B vssd1 vssd1 vccd1 vccd1 _2861_/X sky130_fd_sc_hd__or2_1
X_1812_ _1812_/A _1813_/B vssd1 vssd1 vccd1 vccd1 _1812_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_30_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2792_ _2830_/B vssd1 vssd1 vccd1 vccd1 _2806_/B sky130_fd_sc_hd__clkbuf_1
X_1743_ _3558_/Q vssd1 vssd1 vccd1 vccd1 _2189_/B sky130_fd_sc_hd__inv_2
XFILLER_7_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2701__A _2775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1674_ _3215_/A _2407_/A _1673_/Y _3506_/Q vssd1 vssd1 vccd1 vccd1 _1674_/X sky130_fd_sc_hd__a22o_1
X_3413_ _3414_/CLK _3413_/D vssd1 vssd1 vccd1 vccd1 _3413_/Q sky130_fd_sc_hd__dfxtp_1
X_3344_ _3356_/CLK _3344_/D vssd1 vssd1 vccd1 vccd1 _3344_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3275_ _3275_/A vssd1 vssd1 vccd1 vccd1 _3534_/D sky130_fd_sc_hd__clkbuf_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2226_ _2222_/Y _2037_/B _2262_/A vssd1 vssd1 vccd1 vccd1 _2226_/X sky130_fd_sc_hd__o21a_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2157_ _2161_/A _2161_/B vssd1 vssd1 vccd1 vccd1 _2157_/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_212 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2088_ _3339_/Q _2089_/B vssd1 vssd1 vccd1 vccd1 _2093_/B sky130_fd_sc_hd__or2_1
XFILLER_53_267 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_175 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2330__B _2330_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_2_1__f_net107_A clkbuf_0_net107/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output68_A _3253_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrlbp_macro_191 vssd1 vssd1 vccd1 vccd1 rlbp_macro_191/HI io_out[34] sky130_fd_sc_hd__conb_1
XFILLER_79_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3060_ _3312_/Q _2988_/X _3012_/A _3059_/X vssd1 vssd1 vccd1 vccd1 _3060_/X sky130_fd_sc_hd__a211o_1
Xrlbp_macro_180 vssd1 vssd1 vccd1 vccd1 rlbp_macro_180/HI io_out[9] sky130_fd_sc_hd__conb_1
XFILLER_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2011_ _2011_/A _2011_/B vssd1 vssd1 vccd1 vccd1 _2013_/B sky130_fd_sc_hd__xor2_1
XFILLER_94_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2913_ _2951_/A _2923_/B vssd1 vssd1 vccd1 vccd1 _2913_/X sky130_fd_sc_hd__or2_1
X_2844_ _2953_/A _2850_/B vssd1 vssd1 vccd1 vccd1 _2844_/X sky130_fd_sc_hd__or2_1
XFILLER_31_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2775_ _2775_/A _2778_/B vssd1 vssd1 vccd1 vccd1 _2775_/X sky130_fd_sc_hd__or2_1
XANTENNA__2431__A _3230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1726_ _3493_/Q _1648_/Y _1667_/X _1714_/Y vssd1 vssd1 vccd1 vccd1 _1726_/X sky130_fd_sc_hd__o22a_1
X_1657_ _2026_/B vssd1 vssd1 vccd1 vccd1 _1657_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_100_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3327_ _3332_/CLK _3327_/D vssd1 vssd1 vccd1 vccd1 _3327_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3262__A _3527_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3258_ _3525_/Q _3262_/B _3262_/C vssd1 vssd1 vccd1 vccd1 _3258_/X sky130_fd_sc_hd__or3_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3112__C1 _3111_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2209_ _3403_/Q _2292_/B vssd1 vssd1 vccd1 vccd1 _2210_/B sky130_fd_sc_hd__and2_1
XANTENNA__2466__A1 _3319_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3189_ _3500_/Q _3173_/A _3188_/X _3184_/X vssd1 vssd1 vccd1 vccd1 _3500_/D sky130_fd_sc_hd__o211a_1
XFILLER_39_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2606__A _3234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2979__C _2997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2341__A _3461_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2516__A _2516_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output106_A _2381_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_568 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2560_ _3345_/Q _2556_/X _2559_/X _2547_/X vssd1 vssd1 vccd1 vccd1 _3345_/D sky130_fd_sc_hd__o211a_1
X_2491_ _2568_/A _2491_/B vssd1 vssd1 vccd1 vccd1 _2491_/X sky130_fd_sc_hd__or2_1
XFILLER_101_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_123 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3112_ _3329_/Q _2480_/B _2557_/B _3353_/Q _3111_/X vssd1 vssd1 vccd1 vccd1 _3112_/X
+ sky130_fd_sc_hd__a221o_1
X_3043_ _3347_/Q _3000_/X _2837_/A _3431_/Q vssd1 vssd1 vccd1 vccd1 _3043_/X sky130_fd_sc_hd__a22o_1
XFILLER_82_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2999__A2 _2996_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2426__A _3227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2620__A1 _3363_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2827_ _2975_/A _2830_/B vssd1 vssd1 vccd1 vccd1 _2827_/X sky130_fd_sc_hd__or2_1
X_2758_ _2758_/A _2765_/B vssd1 vssd1 vccd1 vccd1 _2758_/X sky130_fd_sc_hd__or2_1
X_1709_ hold5/X vssd1 vssd1 vccd1 vccd1 _2385_/C sky130_fd_sc_hd__clkbuf_2
X_2689_ _3384_/Q _2678_/X _2688_/X _2686_/X vssd1 vssd1 vccd1 vccd1 _3384_/D sky130_fd_sc_hd__o211a_1
XFILLER_48_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2336__A _3455_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1662__A2 _2115_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2611__A1 _3361_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_104 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2223__B_N _2105_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1991_ _3326_/Q _1991_/B vssd1 vssd1 vccd1 vccd1 _1992_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__2602__A1 _3358_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_590 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2612_ _2612_/A vssd1 vssd1 vccd1 vccd1 _2612_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_70_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2543_ _3341_/Q _2533_/X _2542_/X _2536_/X vssd1 vssd1 vccd1 vccd1 _3341_/D sky130_fd_sc_hd__o211a_1
XANTENNA__3805__A _3805_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2474_ _2552_/A _2943_/A vssd1 vssd1 vccd1 vccd1 _2981_/A sky130_fd_sc_hd__nor2_1
XANTENNA__2669__A1 _3378_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3026_ _3334_/Q _2516_/A _2640_/A _3370_/Q _3025_/X vssd1 vssd1 vccd1 vccd1 _3027_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__2156__A _3373_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_118 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1995__A _3321_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1883__A2 _1878_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2066__A _3342_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2190_ _3395_/Q _2190_/B vssd1 vssd1 vccd1 vccd1 _2247_/A sky130_fd_sc_hd__xor2_1
XFILLER_2_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_490 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1974_ _3302_/Q vssd1 vssd1 vccd1 vccd1 _1974_/X sky130_fd_sc_hd__buf_2
X_2526_ _3334_/Q _2518_/X _2525_/X _2523_/X vssd1 vssd1 vccd1 vccd1 _3334_/D sky130_fd_sc_hd__o211a_1
X_2457_ _3181_/A vssd1 vssd1 vccd1 vccd1 _2578_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_29_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2388_ _2388_/A vssd1 vssd1 vccd1 vccd1 _3298_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3067__A1 _3397_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3009_ _3441_/Q _2875_/B _3160_/B _3489_/Q vssd1 vssd1 vccd1 vccd1 _3009_/X sky130_fd_sc_hd__a22o_1
XFILLER_36_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3058__A1 _3396_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1690_ _3502_/Q _2385_/A vssd1 vssd1 vccd1 vccd1 _1690_/X sky130_fd_sc_hd__or2_1
XFILLER_7_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output98_A _3560_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3360_ _3377_/CLK _3360_/D vssd1 vssd1 vccd1 vccd1 _3360_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2311_ _2347_/B _2343_/A _2308_/Y _2310_/X vssd1 vssd1 vccd1 vccd1 _2311_/X sky130_fd_sc_hd__a31o_1
XFILLER_97_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3291_ _3291_/D _2356_/X vssd1 vssd1 vccd1 vccd1 _3293_/D sky130_fd_sc_hd__dlxtn_1
X_2242_ _2242_/A _2242_/B vssd1 vssd1 vccd1 vccd1 _2255_/C sky130_fd_sc_hd__xnor2_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2173_ _3376_/Q _2173_/B vssd1 vssd1 vccd1 vccd1 _2174_/B sky130_fd_sc_hd__xnor2_1
XFILLER_38_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2418__B _2983_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3049__B2 _3492_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2434__A _3232_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_379 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1957_ _3318_/Q _2121_/B vssd1 vssd1 vccd1 vccd1 _1986_/B sky130_fd_sc_hd__xnor2_1
X_1888_ _2145_/A _3424_/Q vssd1 vssd1 vccd1 vccd1 _1888_/X sky130_fd_sc_hd__or2b_1
XANTENNA__2980__B1 _3006_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3558_ _3559_/CLK _3558_/D _3287_/Y vssd1 vssd1 vccd1 vccd1 _3558_/Q sky130_fd_sc_hd__dfrtp_1
X_2509_ _2586_/A _2509_/B vssd1 vssd1 vccd1 vccd1 _2509_/X sky130_fd_sc_hd__or2_1
XFILLER_88_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3489_ _3491_/CLK _3489_/D vssd1 vssd1 vccd1 vccd1 _3489_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3288__A1 hold2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_0__f_net107_A clkbuf_0_net107/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2609__A _3236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_107 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3175__A _3238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrlbp_macro_340 vssd1 vssd1 vccd1 vccd1 rlbp_macro_340/HI wbs_dat_o[26] sky130_fd_sc_hd__conb_1
XFILLER_47_210 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_9_net107 clkbuf_leaf_9_net107/A vssd1 vssd1 vccd1 vccd1 _3396_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_6 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2860_ _3436_/Q _2853_/X _2859_/X _2851_/X vssd1 vssd1 vccd1 vccd1 _3436_/D sky130_fd_sc_hd__o211a_1
XFILLER_30_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1811_ _3433_/Q _1811_/B vssd1 vssd1 vccd1 vccd1 _1822_/C sky130_fd_sc_hd__xnor2_1
XFILLER_30_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2791_ _2875_/A _2791_/B vssd1 vssd1 vccd1 vccd1 _2830_/B sky130_fd_sc_hd__nand2_1
XANTENNA__3203__A1 _2565_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1742_ _1742_/A vssd1 vssd1 vccd1 vccd1 _3550_/D sky130_fd_sc_hd__clkbuf_1
X_1673_ _2399_/A vssd1 vssd1 vccd1 vccd1 _1673_/Y sky130_fd_sc_hd__inv_2
X_3412_ _3414_/CLK _3412_/D vssd1 vssd1 vccd1 vccd1 _3412_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3343_ _3356_/CLK _3343_/D vssd1 vssd1 vccd1 vccd1 _3343_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3274_ _2378_/A _3296_/Q vssd1 vssd1 vccd1 vccd1 _3275_/A sky130_fd_sc_hd__and2b_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_187 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2225_ _3399_/Q _2288_/B vssd1 vssd1 vccd1 vccd1 _2262_/A sky130_fd_sc_hd__and2b_1
XANTENNA__2429__A _2559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2156_ _3373_/Q _2156_/B vssd1 vssd1 vccd1 vccd1 _2168_/C sky130_fd_sc_hd__xnor2_1
XFILLER_53_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2087_ _2087_/A _2087_/B vssd1 vssd1 vccd1 vccd1 _2089_/B sky130_fd_sc_hd__xnor2_1
XFILLER_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2164__A _3370_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2989_ _2427_/A _2988_/X _3264_/B vssd1 vssd1 vccd1 vccd1 _3074_/A sky130_fd_sc_hd__a21boi_1
XFILLER_21_187 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2330__C _2330_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2984__D _3024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2339__A _2339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2802__A _3234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrlbp_macro_192 vssd1 vssd1 vccd1 vccd1 rlbp_macro_192/HI io_out[35] sky130_fd_sc_hd__conb_1
XFILLER_67_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrlbp_macro_170 vssd1 vssd1 vccd1 vccd1 rlbp_macro_170/HI io_oeb[37] sky130_fd_sc_hd__conb_1
XFILLER_0_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrlbp_macro_181 vssd1 vssd1 vccd1 vccd1 rlbp_macro_181/HI io_out[10] sky130_fd_sc_hd__conb_1
X_2010_ _1945_/C _1988_/B _1976_/Y vssd1 vssd1 vccd1 vccd1 _2011_/B sky130_fd_sc_hd__a21o_1
XFILLER_82_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2111__A_N _1774_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2227__A2 _2037_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2912_ _2941_/B vssd1 vssd1 vccd1 vccd1 _2923_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_92_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2843_ _3429_/Q _2839_/X _2842_/X _2832_/X vssd1 vssd1 vccd1 vccd1 _3429_/D sky130_fd_sc_hd__o211a_1
XANTENNA__3808__A _3808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2712__A _2788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2774_ _3412_/Q _2767_/X _2773_/X _2763_/X vssd1 vssd1 vccd1 vccd1 _3412_/D sky130_fd_sc_hd__o211a_1
X_1725_ _3498_/Q _1922_/A vssd1 vssd1 vccd1 vccd1 _1725_/Y sky130_fd_sc_hd__nor2_1
X_1656_ _3300_/Q vssd1 vssd1 vccd1 vccd1 _2026_/B sky130_fd_sc_hd__clkbuf_4
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3326_ _3332_/CLK _3326_/D vssd1 vssd1 vccd1 vccd1 _3326_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3262__B _3262_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2159__A _3372_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3257_ _3525_/Q _1707_/A _3251_/X _3256_/X vssd1 vssd1 vccd1 vccd1 _3525_/D sky130_fd_sc_hd__o211a_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3112__B1 _2557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2208_ _3403_/Q _2291_/B vssd1 vssd1 vccd1 vccd1 _2210_/A sky130_fd_sc_hd__nor2_1
XFILLER_73_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3188_ _3188_/A _3188_/B vssd1 vssd1 vccd1 vccd1 _3188_/X sky130_fd_sc_hd__or2_1
XFILLER_39_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2139_ _2138_/X _2129_/A _2129_/B vssd1 vssd1 vccd1 vccd1 _2139_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_22_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2622__A _2773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2979__D _3053_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2284__A_N _2285_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input12_A la_data_in[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_412 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_456 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2393__A1 _2395_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2490_ _3324_/Q _2479_/X _2489_/X _2487_/X vssd1 vssd1 vccd1 vccd1 _3324_/D sky130_fd_sc_hd__o211a_1
XFILLER_4_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3111_ _3377_/Q _2640_/A _2715_/B _3401_/Q vssd1 vssd1 vccd1 vccd1 _3111_/X sky130_fd_sc_hd__a22o_1
XFILLER_67_135 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3042_ _3042_/A vssd1 vssd1 vccd1 vccd1 _3042_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2707__A _2782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2442__A _2442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2826_ _3186_/A vssd1 vssd1 vccd1 vccd1 _2975_/A sky130_fd_sc_hd__clkbuf_2
X_2757_ _3405_/Q _2753_/X _2756_/X _2743_/X vssd1 vssd1 vccd1 vccd1 _3405_/D sky130_fd_sc_hd__o211a_1
X_2688_ _2762_/A _2690_/B vssd1 vssd1 vccd1 vccd1 _2688_/X sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_4_net107_A clkbuf_leaf_9_net107/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1708_ input30/X hold4/X _1708_/S vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__mux2_2
XFILLER_2_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_603 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input4_A io_in[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3309_ _3322_/CLK _3309_/D vssd1 vssd1 vccd1 vccd1 _3309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2617__A _3241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3183__A _3183_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_455 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_116 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2527__A _2563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_160 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1990_ _1988_/A _1988_/B _1972_/X vssd1 vssd1 vccd1 vccd1 _1992_/A sky130_fd_sc_hd__a21bo_1
XFILLER_20_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2611_ _3361_/Q _2593_/X _2610_/X _2601_/X vssd1 vssd1 vccd1 vccd1 _3361_/D sky130_fd_sc_hd__o211a_1
X_2542_ _2578_/A _2544_/B vssd1 vssd1 vccd1 vccd1 _2542_/X sky130_fd_sc_hd__or2_1
X_2473_ _2511_/A _2551_/B vssd1 vssd1 vccd1 vccd1 _2943_/A sky130_fd_sc_hd__or2_2
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3025_ _3382_/Q _2676_/A _3033_/A _3522_/Q vssd1 vssd1 vccd1 vccd1 _3025_/X sky130_fd_sc_hd__a22o_1
XFILLER_55_127 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2437__A _3234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3094__A2 _3041_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3789_ _3789_/A vssd1 vssd1 vccd1 vccd1 _3789_/X sky130_fd_sc_hd__clkbuf_1
X_2809_ _3238_/A vssd1 vssd1 vccd1 vccd1 _2964_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_3_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_422 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_267 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_436 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_90 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1973_ _3314_/Q _2106_/B vssd1 vssd1 vccd1 vccd1 _1973_/X sky130_fd_sc_hd__or2b_1
XFILLER_33_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2720__A _2758_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2525_ _2561_/A _2531_/B vssd1 vssd1 vccd1 vccd1 _2525_/X sky130_fd_sc_hd__or2_1
X_2456_ _3316_/Q _2446_/X _2455_/X _2444_/X vssd1 vssd1 vccd1 vccd1 _3316_/D sky130_fd_sc_hd__o211a_1
XFILLER_56_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2387_ _2385_/X _2387_/B _2387_/C vssd1 vssd1 vccd1 vccd1 _2388_/A sky130_fd_sc_hd__and3b_1
XFILLER_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3067__A2 _3041_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_299 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3008_ _3008_/A vssd1 vssd1 vccd1 vccd1 _3160_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_101_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2630__A _3186_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2502__A1 _3328_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2805__A _3236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2569__A1 _3349_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1792__A2 _1698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2540__A _2576_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3290_ hold2/X _3281_/A _3282_/A vssd1 vssd1 vccd1 vccd1 _3290_/Y sky130_fd_sc_hd__a21oi_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2310_ _2309_/X _2289_/B _2286_/B vssd1 vssd1 vccd1 vccd1 _2310_/X sky130_fd_sc_hd__a21o_1
X_2241_ _3390_/Q _2241_/B vssd1 vssd1 vccd1 vccd1 _2242_/B sky130_fd_sc_hd__xnor2_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2172_ _2175_/A _2175_/B _2113_/B vssd1 vssd1 vccd1 vccd1 _2174_/A sky130_fd_sc_hd__a21oi_1
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2715__A _2875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1956_ _1956_/A _1956_/B vssd1 vssd1 vccd1 vccd1 _2007_/A sky130_fd_sc_hd__nor2_1
X_1887_ _1884_/X _1885_/X _1886_/X vssd1 vssd1 vccd1 vccd1 _1887_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__3436__CLK _3436_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3557_ _3557_/D _2366_/X vssd1 vssd1 vccd1 vccd1 _3559_/D sky130_fd_sc_hd__dlxtn_1
XFILLER_88_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2732__A1 _3398_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2508_ _3331_/Q _2493_/A _2507_/X _2501_/X vssd1 vssd1 vccd1 vccd1 _3331_/D sky130_fd_sc_hd__o211a_1
X_3488_ _3529_/CLK _3488_/D vssd1 vssd1 vccd1 vccd1 _3488_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3281__A _3281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3288__A2 _3281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2439_ _3312_/Q _2425_/X _2438_/X _2370_/X vssd1 vssd1 vccd1 vccd1 _3312_/D sky130_fd_sc_hd__o211a_1
XFILLER_56_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2047__D _2074_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2625__A _2775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2723__A1 _3395_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input42_A wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrlbp_macro_341 vssd1 vssd1 vccd1 vccd1 rlbp_macro_341/HI wbs_dat_o[27] sky130_fd_sc_hd__conb_1
Xrlbp_macro_330 vssd1 vssd1 vccd1 vccd1 rlbp_macro_330/HI wbs_dat_o[16] sky130_fd_sc_hd__conb_1
XFILLER_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2535__A _2572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1810_ _1810_/A _1810_/B vssd1 vssd1 vccd1 vccd1 _1811_/B sky130_fd_sc_hd__xnor2_1
X_2790_ _3227_/A vssd1 vssd1 vccd1 vccd1 _2951_/A sky130_fd_sc_hd__clkbuf_2
X_1741_ _3554_/Q _3553_/Q vssd1 vssd1 vccd1 vccd1 _1742_/A sky130_fd_sc_hd__and2b_1
XFILLER_7_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_380 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1672_ _2282_/B vssd1 vssd1 vccd1 vccd1 _2399_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3411_ _3414_/CLK _3411_/D vssd1 vssd1 vccd1 vccd1 _3411_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__3085__B _3085_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3342_ _3516_/CLK _3342_/D vssd1 vssd1 vccd1 vccd1 _3342_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3273_ _3273_/A vssd1 vssd1 vccd1 vccd1 _3533_/D sky130_fd_sc_hd__clkbuf_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_199 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2224_ _2223_/X _2203_/B _2201_/X vssd1 vssd1 vccd1 vccd1 _2224_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_38_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2155_ _2155_/A _2155_/B vssd1 vssd1 vccd1 vccd1 _2156_/B sky130_fd_sc_hd__xnor2_1
XFILLER_66_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2086_ _2041_/A _2068_/B _2062_/Y vssd1 vssd1 vccd1 vccd1 _2087_/B sky130_fd_sc_hd__a21o_1
XFILLER_22_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2988_ _2988_/A vssd1 vssd1 vccd1 vccd1 _2988_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3293__RESET_B _2370_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1939_ _3304_/Q _3316_/Q vssd1 vssd1 vccd1 vccd1 _1941_/A sky130_fd_sc_hd__and2b_1
XANTENNA_clkbuf_leaf_11_net107_A clkbuf_leaf_9_net107/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2181__A2 _1834_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3197__A1 _2561_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3186__A _3186_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrlbp_macro_160 vssd1 vssd1 vccd1 vccd1 rlbp_macro_160/HI io_oeb[27] sky130_fd_sc_hd__conb_1
Xrlbp_macro_193 vssd1 vssd1 vccd1 vccd1 rlbp_macro_193/HI io_out[36] sky130_fd_sc_hd__conb_1
Xrlbp_macro_171 vssd1 vssd1 vccd1 vccd1 rlbp_macro_171/HI io_out[0] sky130_fd_sc_hd__conb_1
XFILLER_0_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrlbp_macro_182 vssd1 vssd1 vccd1 vccd1 rlbp_macro_182/HI io_out[11] sky130_fd_sc_hd__conb_1
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2265__A _3389_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2911_ _3160_/A _2911_/B vssd1 vssd1 vccd1 vccd1 _2941_/B sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_11_net107 clkbuf_leaf_9_net107/A vssd1 vssd1 vccd1 vccd1 _3400_/CLK sky130_fd_sc_hd__clkbuf_16
X_2842_ _2951_/A _2850_/B vssd1 vssd1 vccd1 vccd1 _2842_/X sky130_fd_sc_hd__or2_1
X_2773_ _2773_/A _2778_/B vssd1 vssd1 vccd1 vccd1 _2773_/X sky130_fd_sc_hd__or2_1
X_1724_ _3498_/Q _2121_/B vssd1 vssd1 vccd1 vccd1 _1724_/X sky130_fd_sc_hd__and2_1
XANTENNA__2935__A1 _3461_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1655_ _1932_/B vssd1 vssd1 vccd1 vccd1 _2115_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_98_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3325_ _3332_/CLK _3325_/D vssd1 vssd1 vccd1 vccd1 _3325_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3256_ _3524_/Q _3256_/B _3256_/C vssd1 vssd1 vccd1 vccd1 _3256_/X sky130_fd_sc_hd__or3_1
XANTENNA__3262__C _3262_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_147 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2207_ _2261_/B _2260_/A vssd1 vssd1 vccd1 vccd1 _2212_/B sky130_fd_sc_hd__nor2_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3112__B2 _3353_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3187_ _3499_/Q _3173_/A _3186_/X _3184_/X vssd1 vssd1 vccd1 vccd1 _3499_/D sky130_fd_sc_hd__o211a_1
X_2138_ _3359_/Q _2389_/A vssd1 vssd1 vccd1 vccd1 _2138_/X sky130_fd_sc_hd__or2b_1
XFILLER_39_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2069_ _3337_/Q _2069_/B vssd1 vssd1 vccd1 vccd1 _2083_/B sky130_fd_sc_hd__xnor2_1
XFILLER_54_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2424__B_N _3225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2903__A _2977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_431 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3103__A1 _3364_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2085__A _3341_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_424 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2813__A _3241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_468 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3110_ _3484_/Q _3074_/X _3109_/X _3098_/X vssd1 vssd1 vccd1 vccd1 _3484_/D sky130_fd_sc_hd__o211a_1
XFILLER_68_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3041_ _3041_/A vssd1 vssd1 vccd1 vccd1 _3041_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_75_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_372 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_548 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2825_ _3426_/Q _2808_/X _2824_/X _2815_/X vssd1 vssd1 vccd1 vccd1 _3426_/D sky130_fd_sc_hd__o211a_1
X_2756_ _2756_/A _2765_/B vssd1 vssd1 vccd1 vccd1 _2756_/X sky130_fd_sc_hd__or2_1
X_2687_ _3383_/Q _2678_/X _2685_/X _2686_/X vssd1 vssd1 vccd1 vccd1 _3383_/D sky130_fd_sc_hd__o211a_1
X_1707_ _1707_/A vssd1 vssd1 vccd1 vccd1 _3807_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_98_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3308_ _3308_/CLK _3308_/D vssd1 vssd1 vccd1 vccd1 _3308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3239_ _3251_/A vssd1 vssd1 vccd1 vccd1 _3239_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_73_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2633__A _3188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_128 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_512 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output111_A _3523_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2610_ _2765_/A _2610_/B vssd1 vssd1 vccd1 vccd1 _2610_/X sky130_fd_sc_hd__or2_1
X_2541_ _3340_/Q _2533_/X _2540_/X _2536_/X vssd1 vssd1 vccd1 vccd1 _3340_/D sky130_fd_sc_hd__o211a_1
X_2472_ _2512_/A _2512_/B _2512_/C vssd1 vssd1 vccd1 vccd1 _2551_/B sky130_fd_sc_hd__or3b_1
XFILLER_48_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3024_ _3024_/A vssd1 vssd1 vccd1 vccd1 _3033_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_55_139 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3268__B input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3788_ _3788_/A vssd1 vssd1 vccd1 vccd1 _3788_/X sky130_fd_sc_hd__clkbuf_1
X_2808_ _2808_/A vssd1 vssd1 vccd1 vccd1 _2808_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2739_ _2778_/A _2739_/B vssd1 vssd1 vccd1 vccd1 _2739_/X sky130_fd_sc_hd__or2_1
XFILLER_59_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_434 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2628__A _2778_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2142__B_N _1796_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_279 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2538__A _2574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2273__A _3474_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1972_ _3313_/Q _2105_/B vssd1 vssd1 vccd1 vccd1 _1972_/X sky130_fd_sc_hd__or2b_1
X_2524_ _3333_/Q _2518_/X _2522_/X _2523_/X vssd1 vssd1 vccd1 vccd1 _3333_/D sky130_fd_sc_hd__o211a_1
X_2455_ _2576_/A _2461_/B vssd1 vssd1 vccd1 vccd1 _2455_/X sky130_fd_sc_hd__or2_1
XFILLER_68_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2386_ _2385_/B _2385_/C _2385_/A vssd1 vssd1 vccd1 vccd1 _2387_/B sky130_fd_sc_hd__a21o_1
XFILLER_29_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_36_net107_A _3494_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3007_ _3018_/A vssd1 vssd1 vccd1 vccd1 _3008_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2183__A _3380_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2911__A _3160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_470 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2974__C1 _2971_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2821__A _2970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2240_ _2264_/A _2264_/B _2229_/Y vssd1 vssd1 vccd1 vccd1 _2242_/A sky130_fd_sc_hd__a21o_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2268__A _3391_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2171_ _2114_/A _2155_/B _2144_/Y vssd1 vssd1 vccd1 vccd1 _2175_/B sky130_fd_sc_hd__a21o_1
XFILLER_76_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1955_ _3317_/Q _2119_/B vssd1 vssd1 vccd1 vccd1 _1956_/B sky130_fd_sc_hd__and2_1
X_1886_ _1796_/X _3422_/Q vssd1 vssd1 vccd1 vccd1 _1886_/X sky130_fd_sc_hd__and2b_1
XANTENNA__2980__A2 _3006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3556_ _3556_/D _2366_/X vssd1 vssd1 vccd1 vccd1 _3558_/D sky130_fd_sc_hd__dlxtn_1
XFILLER_88_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2507_ _2584_/A _2509_/B vssd1 vssd1 vccd1 vccd1 _2507_/X sky130_fd_sc_hd__or2_1
XFILLER_88_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3487_ _3529_/CLK _3487_/D vssd1 vssd1 vccd1 vccd1 _3487_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2438_ _2565_/A _2441_/B vssd1 vssd1 vccd1 vccd1 _2438_/X sky130_fd_sc_hd__or2_1
XFILLER_69_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2369_ _2442_/A vssd1 vssd1 vccd1 vccd1 _2742_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__2496__A1 _3326_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2906__A _2983_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2641__A _2788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrlbp_macro_342 vssd1 vssd1 vccd1 vccd1 rlbp_macro_342/HI wbs_dat_o[28] sky130_fd_sc_hd__conb_1
Xrlbp_macro_331 vssd1 vssd1 vccd1 vccd1 rlbp_macro_331/HI wbs_dat_o[17] sky130_fd_sc_hd__conb_1
Xrlbp_macro_320 vssd1 vssd1 vccd1 vccd1 rlbp_macro_320/HI la_data_out[122] sky130_fd_sc_hd__conb_1
XFILLER_94_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2088__A _3339_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input35_A la_data_in[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1740_ _2049_/A vssd1 vssd1 vccd1 vccd1 _3545_/D sky130_fd_sc_hd__clkinv_2
XFILLER_7_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1671_ _3302_/Q vssd1 vssd1 vccd1 vccd1 _2282_/B sky130_fd_sc_hd__clkbuf_4
X_3410_ _3414_/CLK _3410_/D vssd1 vssd1 vccd1 vccd1 _3410_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3341_ _3356_/CLK _3341_/D vssd1 vssd1 vccd1 vccd1 _3341_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3272_ _2378_/X input4/X vssd1 vssd1 vccd1 vccd1 _3273_/A sky130_fd_sc_hd__and2b_1
XANTENNA__3124__C1 _3123_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2223_ _3397_/Q _2105_/B vssd1 vssd1 vccd1 vccd1 _2223_/X sky130_fd_sc_hd__or2b_1
Xclkbuf_leaf_34_net107 _3494_/CLK vssd1 vssd1 vccd1 vccd1 _3544_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2154_ _2154_/A _2154_/B vssd1 vssd1 vccd1 vccd1 _2168_/B sky130_fd_sc_hd__xnor2_1
XFILLER_66_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2726__A _2765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2085_ _3341_/Q _2085_/B vssd1 vssd1 vccd1 vccd1 _2093_/A sky130_fd_sc_hd__xnor2_1
XFILLER_53_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2650__A1 _3371_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2987_ _2993_/A vssd1 vssd1 vccd1 vccd1 _2988_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__2461__A _2582_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1938_ _1938_/A _1938_/B vssd1 vssd1 vccd1 vccd1 _2011_/A sky130_fd_sc_hd__nor2_1
X_1869_ _3427_/Q _2292_/B vssd1 vssd1 vccd1 vccd1 _1870_/B sky130_fd_sc_hd__and2_1
X_3539_ _3539_/CLK _3539_/D _3277_/Y vssd1 vssd1 vccd1 vccd1 _3539_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_76_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2074__C _2074_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrlbp_macro_150 vssd1 vssd1 vccd1 vccd1 rlbp_macro_150/HI io_oeb[17] sky130_fd_sc_hd__conb_1
Xrlbp_macro_194 vssd1 vssd1 vccd1 vccd1 rlbp_macro_194/HI io_out[37] sky130_fd_sc_hd__conb_1
XFILLER_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrlbp_macro_161 vssd1 vssd1 vccd1 vccd1 rlbp_macro_161/HI io_oeb[28] sky130_fd_sc_hd__conb_1
XFILLER_0_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrlbp_macro_172 vssd1 vssd1 vccd1 vccd1 rlbp_macro_172/HI io_out[1] sky130_fd_sc_hd__conb_1
Xrlbp_macro_183 vssd1 vssd1 vccd1 vccd1 rlbp_macro_183/HI io_out[12] sky130_fd_sc_hd__conb_1
XFILLER_57_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2546__A _2584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2910_ _2925_/A vssd1 vssd1 vccd1 vccd1 _2910_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2841_ _2868_/B vssd1 vssd1 vccd1 vccd1 _2850_/B sky130_fd_sc_hd__clkbuf_1
X_2772_ _3411_/Q _2767_/X _2771_/X _2763_/X vssd1 vssd1 vccd1 vccd1 _3411_/D sky130_fd_sc_hd__o211a_1
X_1723_ _3306_/Q vssd1 vssd1 vccd1 vccd1 _2121_/B sky130_fd_sc_hd__clkbuf_4
X_1654_ _1654_/A vssd1 vssd1 vccd1 vccd1 _1932_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_98_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3324_ _3486_/CLK _3324_/D vssd1 vssd1 vccd1 vccd1 _3324_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3255_ _3524_/Q _3807_/A _3251_/X _3254_/X vssd1 vssd1 vccd1 vccd1 _3524_/D sky130_fd_sc_hd__o211a_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2206_ _3399_/Q _2206_/B vssd1 vssd1 vccd1 vccd1 _2260_/A sky130_fd_sc_hd__xor2_2
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3186_ _3186_/A _3188_/B vssd1 vssd1 vccd1 vccd1 _3186_/X sky130_fd_sc_hd__or2_1
XFILLER_93_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2137_ _2163_/A _2165_/B _2136_/X vssd1 vssd1 vccd1 vccd1 _2161_/B sky130_fd_sc_hd__a21o_1
XFILLER_54_546 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1674__A2 _2407_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2068_ _2068_/A _2068_/B vssd1 vssd1 vccd1 vccd1 _2069_/B sky130_fd_sc_hd__xnor2_1
XFILLER_26_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2623__A1 _3364_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2191__A _3396_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3103__A2 _2595_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_436 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_95 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3040_ _3323_/Q _2477_/A _2751_/A _3407_/Q _3039_/X vssd1 vssd1 vccd1 vccd1 _3040_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_48_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2605__A1 _3359_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_270 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2824_ _2973_/A _2824_/B vssd1 vssd1 vccd1 vccd1 _2824_/X sky130_fd_sc_hd__or2_1
X_2755_ _2782_/B vssd1 vssd1 vccd1 vccd1 _2765_/B sky130_fd_sc_hd__clkbuf_1
X_2686_ _2731_/A vssd1 vssd1 vccd1 vccd1 _2686_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1706_ _3262_/B _3262_/C vssd1 vssd1 vccd1 vccd1 _1707_/A sky130_fd_sc_hd__nor2_1
XFILLER_86_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3307_ _3307_/CLK _3307_/D vssd1 vssd1 vccd1 vccd1 _3307_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3238_ _3238_/A _3243_/B vssd1 vssd1 vccd1 vccd1 _3238_/X sky130_fd_sc_hd__or2_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2186__A _3379_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3169_ _3492_/Q _3159_/X _3168_/X _3156_/X vssd1 vssd1 vccd1 vccd1 _3492_/D sky130_fd_sc_hd__o211a_1
XFILLER_39_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2914__A _3199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2824__A _2973_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2540_ _2576_/A _2544_/B vssd1 vssd1 vccd1 vccd1 _2540_/X sky130_fd_sc_hd__or2_1
XFILLER_5_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2471_ _3160_/A vssd1 vssd1 vccd1 vccd1 _3223_/A sky130_fd_sc_hd__buf_2
XFILLER_79_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3079__A1 _3446_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3023_ _3394_/Q _2711_/A _3056_/A _3502_/Q vssd1 vssd1 vccd1 vccd1 _3027_/C sky130_fd_sc_hd__a22o_1
XFILLER_48_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3787_ _3787_/A vssd1 vssd1 vccd1 vccd1 _3787_/X sky130_fd_sc_hd__clkbuf_1
X_2807_ _3421_/Q _2789_/X _2806_/X _2797_/X vssd1 vssd1 vccd1 vccd1 _3421_/D sky130_fd_sc_hd__o211a_1
X_2738_ _3401_/Q _2728_/X _2737_/X _2731_/X vssd1 vssd1 vccd1 vccd1 _3401_/D sky130_fd_sc_hd__o211a_1
X_2669_ _3378_/Q _2656_/X _2666_/X _2668_/X vssd1 vssd1 vccd1 vccd1 _3378_/D sky130_fd_sc_hd__o211a_1
XFILLER_59_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1813__A _3429_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2909__A _3158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_107 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_490 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3242__A1 _3527_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input65_A wbs_stb_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1723__A _3306_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1936__A_N _3315_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_398 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_368 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3233__A1 _3523_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1971_ _1966_/Y _1878_/X _1959_/A _1999_/B _1970_/X vssd1 vssd1 vccd1 vccd1 _1988_/B
+ sky130_fd_sc_hd__a221o_2
XANTENNA__2273__B _3306_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2523_ _2566_/A vssd1 vssd1 vccd1 vccd1 _2523_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_291 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2454_ _3243_/A vssd1 vssd1 vccd1 vccd1 _2576_/A sky130_fd_sc_hd__clkbuf_2
X_2385_ _2385_/A _2385_/B _2385_/C vssd1 vssd1 vccd1 vccd1 _2385_/X sky130_fd_sc_hd__and3_1
XFILLER_68_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput1 CMP vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3006_ _3006_/A _3006_/B vssd1 vssd1 vccd1 vccd1 _3018_/A sky130_fd_sc_hd__nor2_1
XFILLER_64_493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2464__A _3186_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1808__A _3434_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2639__A _2997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_600 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_482 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2374__A _3281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1977__B_N _3316_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2549__A _2586_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_6 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2170_ _3377_/Q _2170_/B vssd1 vssd1 vccd1 vccd1 _2178_/A sky130_fd_sc_hd__xnor2_1
XFILLER_38_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3206__A1 _2568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1954_ _3317_/Q _2118_/B vssd1 vssd1 vccd1 vccd1 _1956_/A sky130_fd_sc_hd__nor2_1
X_1885_ _3422_/Q _1796_/X vssd1 vssd1 vccd1 vccd1 _1885_/X sky130_fd_sc_hd__or2b_1
X_3555_ _3555_/D _2366_/X vssd1 vssd1 vccd1 vccd1 _3555_/Q sky130_fd_sc_hd__dlxtn_1
X_3486_ _3486_/CLK _3486_/D vssd1 vssd1 vccd1 vccd1 _3486_/Q sky130_fd_sc_hd__dfxtp_1
X_2506_ _3330_/Q _2493_/X _2505_/X _2501_/X vssd1 vssd1 vccd1 vccd1 _3330_/D sky130_fd_sc_hd__o211a_1
X_2437_ _3234_/A vssd1 vssd1 vccd1 vccd1 _2565_/A sky130_fd_sc_hd__buf_2
XFILLER_69_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2368_ _2368_/A vssd1 vssd1 vccd1 vccd1 _2368_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_84_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2299_ _3474_/Q vssd1 vssd1 vccd1 vccd1 _2299_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2906__B _3006_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2641__B _2643_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrlbp_macro_332 vssd1 vssd1 vccd1 vccd1 rlbp_macro_332/HI wbs_dat_o[18] sky130_fd_sc_hd__conb_1
Xrlbp_macro_343 vssd1 vssd1 vccd1 vccd1 rlbp_macro_343/HI wbs_dat_o[29] sky130_fd_sc_hd__conb_1
Xrlbp_macro_310 vssd1 vssd1 vccd1 vccd1 rlbp_macro_310/HI la_data_out[112] sky130_fd_sc_hd__conb_1
Xrlbp_macro_321 vssd1 vssd1 vccd1 vccd1 rlbp_macro_321/HI la_data_out[123] sky130_fd_sc_hd__conb_1
XANTENNA__2369__A _2442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2287__A_N _2206_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input28_A la_data_in[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1670_ _3305_/Q vssd1 vssd1 vccd1 vccd1 _2407_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_7_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output96_A _3535_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3340_ _3520_/CLK _3340_/D vssd1 vssd1 vccd1 vccd1 _3340_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3271_ _3271_/A vssd1 vssd1 vccd1 vccd1 _3532_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3124__B1 _2557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2222_ _3400_/Q vssd1 vssd1 vccd1 vccd1 _2222_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2153_ _3374_/Q _2153_/B vssd1 vssd1 vccd1 vccd1 _2154_/B sky130_fd_sc_hd__xnor2_1
XFILLER_66_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2084_ _2084_/A _2084_/B vssd1 vssd1 vccd1 vccd1 _2085_/B sky130_fd_sc_hd__xor2_1
XANTENNA__2742__A _2742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2986_ _2986_/A _2986_/B vssd1 vssd1 vccd1 vccd1 _2993_/A sky130_fd_sc_hd__nor2_1
XANTENNA__3060__C1 _3059_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1937_ _2288_/B _3315_/Q vssd1 vssd1 vccd1 vccd1 _1938_/B sky130_fd_sc_hd__and2b_1
X_1868_ _3427_/Q _2291_/B vssd1 vssd1 vccd1 vccd1 _1870_/A sky130_fd_sc_hd__nor2_1
X_3538_ _3539_/CLK _3538_/D _3276_/Y vssd1 vssd1 vccd1 vccd1 _3538_/Q sky130_fd_sc_hd__dfrtp_1
X_1799_ _1795_/X _1797_/X _1798_/X vssd1 vssd1 vccd1 vccd1 _1799_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_1_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3469_ _3469_/CLK _3469_/D vssd1 vssd1 vccd1 vccd1 _3469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_20_net107_A clkbuf_2_3__f_net107/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2917__A _2953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrlbp_macro_140 vssd1 vssd1 vccd1 vccd1 rlbp_macro_140/HI io_oeb[7] sky130_fd_sc_hd__conb_1
Xrlbp_macro_151 vssd1 vssd1 vccd1 vccd1 rlbp_macro_151/HI io_oeb[18] sky130_fd_sc_hd__conb_1
XFILLER_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrlbp_macro_173 vssd1 vssd1 vccd1 vccd1 rlbp_macro_173/HI io_out[2] sky130_fd_sc_hd__conb_1
Xrlbp_macro_162 vssd1 vssd1 vccd1 vccd1 rlbp_macro_162/HI io_oeb[29] sky130_fd_sc_hd__conb_1
Xrlbp_macro_184 vssd1 vssd1 vccd1 vccd1 rlbp_macro_184/HI io_out[13] sky130_fd_sc_hd__conb_1
XFILLER_48_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrlbp_macro_195 vssd1 vssd1 vccd1 vccd1 rlbp_macro_195/HI irq[0] sky130_fd_sc_hd__conb_1
XANTENNA__2827__A _2975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2840_ _2875_/A _2840_/B vssd1 vssd1 vccd1 vccd1 _2868_/B sky130_fd_sc_hd__nand2_1
X_2771_ _2771_/A _2778_/B vssd1 vssd1 vccd1 vccd1 _2771_/X sky130_fd_sc_hd__or2_1
XANTENNA__2281__B _2281_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1722_ _3490_/Q _2385_/A vssd1 vssd1 vccd1 vccd1 _1728_/C sky130_fd_sc_hd__xnor2_1
XFILLER_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1653_ _3307_/Q vssd1 vssd1 vccd1 vccd1 _1654_/A sky130_fd_sc_hd__inv_2
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3323_ _3486_/CLK _3323_/D vssd1 vssd1 vccd1 vccd1 _3323_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3254_ _3523_/Q _3256_/B _3256_/C vssd1 vssd1 vccd1 vccd1 _3254_/X sky130_fd_sc_hd__or3_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2205_ _3400_/Q _2285_/B vssd1 vssd1 vccd1 vccd1 _2261_/B sky130_fd_sc_hd__xor2_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2737__A _2775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3185_ _3498_/Q _3173_/X _3183_/X _3184_/X vssd1 vssd1 vccd1 vccd1 _3498_/D sky130_fd_sc_hd__o211a_1
X_2136_ _3358_/Q _2389_/B vssd1 vssd1 vccd1 vccd1 _2136_/X sky130_fd_sc_hd__and2b_1
XFILLER_66_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2067_ _2067_/A _2067_/B vssd1 vssd1 vccd1 vccd1 _2083_/A sky130_fd_sc_hd__xnor2_1
XFILLER_54_558 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2191__B _2191_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2969_ _3472_/Q _2962_/X _2968_/X _2958_/X vssd1 vssd1 vccd1 vccd1 _3472_/D sky130_fd_sc_hd__o211a_1
XFILLER_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2647__A _2758_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2550__A1 _3344_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2557__A _2679_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_396 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2292__A _3475_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2823_ _3183_/A vssd1 vssd1 vccd1 vccd1 _2973_/A sky130_fd_sc_hd__clkbuf_2
X_2754_ _2875_/A _2754_/B vssd1 vssd1 vccd1 vccd1 _2782_/B sky130_fd_sc_hd__nand2_1
X_1705_ _1689_/Y _1690_/X _1694_/Y _1695_/X _1704_/X vssd1 vssd1 vccd1 vccd1 _3262_/C
+ sky130_fd_sc_hd__a221o_2
X_2685_ _2760_/A _2690_/B vssd1 vssd1 vccd1 vccd1 _2685_/X sky130_fd_sc_hd__or2_1
XFILLER_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3306_ _3409_/CLK _3306_/D vssd1 vssd1 vccd1 vccd1 _3306_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3237_ _3525_/Q _3224_/X _3236_/X _3228_/X vssd1 vssd1 vccd1 vccd1 _3517_/D sky130_fd_sc_hd__o211a_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2467__A _3188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3168_ _3234_/A _3170_/B vssd1 vssd1 vccd1 vccd1 _3168_/X sky130_fd_sc_hd__or2_1
X_2119_ _3365_/Q _2119_/B vssd1 vssd1 vccd1 vccd1 _2120_/B sky130_fd_sc_hd__and2_1
XFILLER_54_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3099_ _3483_/Q _3074_/X _3097_/X _3098_/X vssd1 vssd1 vccd1 vccd1 _3483_/D sky130_fd_sc_hd__o211a_1
XFILLER_14_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_580 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2930__A _2966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_436 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input10_A la_data_in[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2840__A _2875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2220__B1 _2389_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2470_ _2470_/A vssd1 vssd1 vccd1 vccd1 _3160_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_68_436 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3022_ _3346_/Q _3000_/X _3021_/X _3430_/Q vssd1 vssd1 vccd1 vccd1 _3027_/B sky130_fd_sc_hd__a22o_1
XFILLER_91_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3786_ input5/X vssd1 vssd1 vccd1 vccd1 _3786_/X sky130_fd_sc_hd__clkbuf_1
X_2806_ _2960_/A _2806_/B vssd1 vssd1 vccd1 vccd1 _2806_/X sky130_fd_sc_hd__or2_1
X_2737_ _2775_/A _2739_/B vssd1 vssd1 vccd1 vccd1 _2737_/X sky130_fd_sc_hd__or2_1
X_2668_ _2731_/A vssd1 vssd1 vccd1 vccd1 _2668_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_99_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2599_ _3230_/A vssd1 vssd1 vccd1 vccd1 _2758_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_101_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input2_A io_in[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_288 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2660__A _2771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_31 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input58_A wbs_dat_i[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2835__A _3006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1970_ _1966_/Y _1698_/A _1969_/X vssd1 vssd1 vccd1 vccd1 _1970_/X sky130_fd_sc_hd__o21a_1
XFILLER_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2522_ _2559_/A _2531_/B vssd1 vssd1 vccd1 vccd1 _2522_/X sky130_fd_sc_hd__or2_1
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2453_ _3315_/Q _2446_/X _2452_/X _2444_/X vssd1 vssd1 vccd1 vccd1 _3315_/D sky130_fd_sc_hd__o211a_1
XFILLER_96_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2384_ _2385_/B _2385_/C _2383_/Y vssd1 vssd1 vccd1 vccd1 _3297_/D sky130_fd_sc_hd__a21oi_1
XFILLER_29_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_17_net107 clkbuf_2_3__f_net107/X vssd1 vssd1 vccd1 vccd1 _3559_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_68_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput2 io_in[15] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_2
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3005_ _3005_/A _3005_/B _3005_/C _3005_/D vssd1 vssd1 vccd1 vccd1 _3005_/X sky130_fd_sc_hd__or4_1
XANTENNA__2745__A _2782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2480__A _3225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_100 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2974__A1 _3474_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3151__A1 _3344_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2565__A _2565_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1953_ _1999_/A _1997_/B vssd1 vssd1 vccd1 vccd1 _1959_/A sky130_fd_sc_hd__and2_1
XFILLER_33_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1884_ _3421_/Q _1794_/X vssd1 vssd1 vccd1 vccd1 _1884_/X sky130_fd_sc_hd__or2b_1
Xclkbuf_leaf_4_net107 clkbuf_leaf_9_net107/A vssd1 vssd1 vccd1 vccd1 _3356_/CLK sky130_fd_sc_hd__clkbuf_16
X_3554_ _3564_/CLK _3554_/D _3286_/Y vssd1 vssd1 vccd1 vccd1 _3554_/Q sky130_fd_sc_hd__dfrtp_1
X_3485_ _3486_/CLK _3485_/D vssd1 vssd1 vccd1 vccd1 _3485_/Q sky130_fd_sc_hd__dfxtp_1
X_2505_ _2582_/A _2505_/B vssd1 vssd1 vccd1 vccd1 _2505_/X sky130_fd_sc_hd__or2_1
XANTENNA__1644__A _1774_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2436_ _3311_/Q _2425_/X _2435_/X _2370_/X vssd1 vssd1 vccd1 vccd1 _3311_/D sky130_fd_sc_hd__o211a_1
XANTENNA__3142__A1 _3499_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2367_ _3564_/Q _3563_/Q vssd1 vssd1 vccd1 vccd1 _2368_/A sky130_fd_sc_hd__and2_1
XFILLER_56_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2298_ _3560_/D _2271_/X _2353_/A _3563_/Q vssd1 vssd1 vccd1 vccd1 _3561_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_29_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2194__B _3393_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1819__A _3432_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2956__A1 _3467_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrlbp_macro_300 vssd1 vssd1 vccd1 vccd1 rlbp_macro_300/HI la_data_out[102] sky130_fd_sc_hd__conb_1
XFILLER_79_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrlbp_macro_333 vssd1 vssd1 vccd1 vccd1 rlbp_macro_333/HI wbs_dat_o[19] sky130_fd_sc_hd__conb_1
Xrlbp_macro_311 vssd1 vssd1 vccd1 vccd1 rlbp_macro_311/HI la_data_out[113] sky130_fd_sc_hd__conb_1
Xrlbp_macro_322 vssd1 vssd1 vccd1 vccd1 rlbp_macro_322/HI la_data_out[124] sky130_fd_sc_hd__conb_1
Xrlbp_macro_344 vssd1 vssd1 vccd1 vccd1 rlbp_macro_344/HI wbs_dat_o[30] sky130_fd_sc_hd__conb_1
XFILLER_94_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3270_ _2378_/X _3533_/Q vssd1 vssd1 vccd1 vccd1 _3271_/A sky130_fd_sc_hd__and2b_1
XFILLER_3_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2221_ _2216_/Y _1878_/X _2213_/A _2247_/B _2220_/X vssd1 vssd1 vccd1 vccd1 _2235_/B
+ sky130_fd_sc_hd__a221o_2
XANTENNA__3124__B2 _3354_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2152_ _2155_/A _2155_/B _2141_/X vssd1 vssd1 vccd1 vccd1 _2154_/A sky130_fd_sc_hd__a21bo_1
XFILLER_16_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2083_ _2083_/A _2083_/B _2083_/C _2083_/D vssd1 vssd1 vccd1 vccd1 _2083_/X sky130_fd_sc_hd__or4_1
XFILLER_93_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_228 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_442 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2985_ _2985_/A _2985_/B _2985_/C _2985_/D vssd1 vssd1 vccd1 vccd1 _2986_/B sky130_fd_sc_hd__or4_1
X_1936_ _3315_/Q _2288_/B vssd1 vssd1 vccd1 vccd1 _1938_/A sky130_fd_sc_hd__and2b_1
X_1867_ _1932_/B vssd1 vssd1 vccd1 vccd1 _2291_/B sky130_fd_sc_hd__clkbuf_4
Xinput60 wbs_dat_i[6] vssd1 vssd1 vccd1 vccd1 _3241_/A sky130_fd_sc_hd__clkbuf_4
X_1798_ _2399_/A _3446_/Q vssd1 vssd1 vccd1 vccd1 _1798_/X sky130_fd_sc_hd__and2b_1
X_3537_ _3537_/D _2358_/X vssd1 vssd1 vccd1 vccd1 _3539_/D sky130_fd_sc_hd__dlxtn_1
XFILLER_1_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_7_net107_A clkbuf_leaf_9_net107/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3468_ _3469_/CLK _3468_/D vssd1 vssd1 vccd1 vccd1 _3468_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3399_ _3400_/CLK _3399_/D vssd1 vssd1 vccd1 vccd1 _3399_/Q sky130_fd_sc_hd__dfxtp_2
X_2419_ input45/X input44/X _2419_/C _2419_/D vssd1 vssd1 vccd1 vccd1 _2420_/C sky130_fd_sc_hd__and4bb_1
XANTENNA__3115__B2 _3509_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input40_A wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrlbp_macro_141 vssd1 vssd1 vccd1 vccd1 rlbp_macro_141/HI io_oeb[8] sky130_fd_sc_hd__conb_1
XFILLER_0_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3106__A1 _3352_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrlbp_macro_174 vssd1 vssd1 vccd1 vccd1 rlbp_macro_174/HI io_out[3] sky130_fd_sc_hd__conb_1
Xrlbp_macro_163 vssd1 vssd1 vccd1 vccd1 rlbp_macro_163/HI io_oeb[30] sky130_fd_sc_hd__conb_1
Xrlbp_macro_152 vssd1 vssd1 vccd1 vccd1 rlbp_macro_152/HI io_oeb[19] sky130_fd_sc_hd__conb_1
Xrlbp_macro_185 vssd1 vssd1 vccd1 vccd1 rlbp_macro_185/HI io_out[14] sky130_fd_sc_hd__conb_1
XANTENNA__3106__B2 _3436_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrlbp_macro_196 vssd1 vssd1 vccd1 vccd1 rlbp_macro_196/HI irq[1] sky130_fd_sc_hd__conb_1
XFILLER_75_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3290__B1 _3282_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2770_ _3410_/Q _2767_/X _2769_/X _2763_/X vssd1 vssd1 vccd1 vccd1 _3410_/D sky130_fd_sc_hd__o211a_1
XFILLER_78_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1721_ _3499_/Q _1932_/B _1645_/Y _3495_/Q _1720_/Y vssd1 vssd1 vccd1 vccd1 _1728_/B
+ sky130_fd_sc_hd__o221a_1
X_1652_ _3507_/Q _1645_/Y _1648_/Y _3505_/Q _1651_/X vssd1 vssd1 vccd1 vccd1 _1686_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_98_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3322_ _3322_/CLK _3322_/D vssd1 vssd1 vccd1 vccd1 _3322_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3253_ _3523_/Q _3253_/A2 _3251_/X _3252_/X vssd1 vssd1 vccd1 vccd1 _3523_/D sky130_fd_sc_hd__o211a_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2204_ _2235_/A _2238_/B vssd1 vssd1 vccd1 vccd1 _2212_/A sky130_fd_sc_hd__and2_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3184_ _3184_/A vssd1 vssd1 vccd1 vccd1 _3184_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_39_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2135_ _2135_/A vssd1 vssd1 vccd1 vccd1 _3551_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1771__A_N _3448_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2066_ _3342_/Q _2066_/B vssd1 vssd1 vccd1 vccd1 _2067_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__2127__A_N _2191_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2968_ _2968_/A _2973_/B vssd1 vssd1 vccd1 vccd1 _2968_/X sky130_fd_sc_hd__or2_1
X_1919_ _1919_/A _1919_/B vssd1 vssd1 vccd1 vccd1 _1920_/D sky130_fd_sc_hd__xnor2_1
X_2899_ _2973_/A _2899_/B vssd1 vssd1 vccd1 vccd1 _2899_/X sky130_fd_sc_hd__or2_1
XFILLER_1_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2145__B_N _3364_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2838__A _3158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2557__B _2557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2302__A2 _2330_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3263__B1 _3264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2292__B _2292_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2822_ _3425_/Q _2808_/X _2821_/X _2815_/X vssd1 vssd1 vccd1 vccd1 _3425_/D sky130_fd_sc_hd__o211a_1
X_2753_ _2767_/A vssd1 vssd1 vccd1 vccd1 _2753_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1704_ _3202_/A _2395_/B _2385_/B _3193_/A _1703_/X vssd1 vssd1 vccd1 vccd1 _1704_/X
+ sky130_fd_sc_hd__a221o_1
X_2684_ _3382_/Q _2678_/X _2683_/X _2668_/X vssd1 vssd1 vccd1 vccd1 _3382_/D sky130_fd_sc_hd__o211a_1
XFILLER_98_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3305_ _3409_/CLK _3305_/D vssd1 vssd1 vccd1 vccd1 _3305_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2748__A _2983_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3236_ _3236_/A _3236_/B vssd1 vssd1 vccd1 vccd1 _3236_/X sky130_fd_sc_hd__or2_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3167_ _3491_/Q _3159_/X _3166_/X _3156_/X vssd1 vssd1 vccd1 vccd1 _3491_/D sky130_fd_sc_hd__o211a_1
XFILLER_81_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2118_ _3365_/Q _2118_/B vssd1 vssd1 vccd1 vccd1 _2120_/A sky130_fd_sc_hd__nor2_1
X_3098_ _3184_/A vssd1 vssd1 vccd1 vccd1 _3098_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2049_ _2049_/A _2049_/B vssd1 vssd1 vccd1 vccd1 _2050_/A sky130_fd_sc_hd__and2_1
XFILLER_42_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_592 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2658__A _2769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2568__A _2568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3021_ _3021_/A vssd1 vssd1 vccd1 vccd1 _3021_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_76_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_186 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2805_ _3236_/A vssd1 vssd1 vccd1 vccd1 _2960_/A sky130_fd_sc_hd__clkbuf_2
X_3785_ _3785_/A vssd1 vssd1 vccd1 vccd1 _3785_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__1647__A _2281_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2736_ _3400_/Q _2728_/X _2735_/X _2731_/X vssd1 vssd1 vccd1 vccd1 _3400_/D sky130_fd_sc_hd__o211a_1
X_2667_ _2742_/A vssd1 vssd1 vccd1 vccd1 _2731_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_99_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2598_ _3357_/Q _2593_/X _2597_/X _2580_/X vssd1 vssd1 vccd1 vccd1 _3357_/D sky130_fd_sc_hd__o211a_1
XANTENNA__2478__A _3223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3219_ _3219_/A _3219_/B vssd1 vssd1 vccd1 vccd1 _3219_/Y sky130_fd_sc_hd__nand2_1
XFILLER_39_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2941__A _2977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2450__A1 _3314_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_43 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3163__C1 _3156_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2521_ _2549_/B vssd1 vssd1 vccd1 vccd1 _2531_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__3154__C1 _3153_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2452_ _2574_/A _2461_/B vssd1 vssd1 vccd1 vccd1 _2452_/X sky130_fd_sc_hd__or2_1
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2383_ _2385_/B _2385_/C _2397_/A vssd1 vssd1 vccd1 vccd1 _2383_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_96_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput3 io_in[16] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_2
X_3004_ _3393_/Q _2711_/A _3056_/A _3501_/Q vssd1 vssd1 vccd1 vccd1 _3005_/D sky130_fd_sc_hd__a22o_1
XFILLER_83_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2719_ _3393_/Q _2713_/X _2717_/X _2718_/X vssd1 vssd1 vccd1 vccd1 _3393_/D sky130_fd_sc_hd__o211a_1
XANTENNA_clkbuf_leaf_14_net107_A clkbuf_2_3__f_net107/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1840__A _3440_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2936__A _2973_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2671__A1 _3379_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_23_net107 _3436_/CLK vssd1 vssd1 vccd1 vccd1 _3474_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3151__A2 _2996_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2846__A _2955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2414__A1 _2042_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1952_ _3312_/Q _3300_/Q vssd1 vssd1 vccd1 vccd1 _1997_/B sky130_fd_sc_hd__xnor2_1
XFILLER_33_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1883_ _1876_/Y _1878_/X _1854_/A _1907_/B _1882_/X vssd1 vssd1 vccd1 vccd1 _1895_/B
+ sky130_fd_sc_hd__a221o_2
X_3553_ _3564_/CLK _3553_/D _3285_/Y vssd1 vssd1 vccd1 vccd1 _3553_/Q sky130_fd_sc_hd__dfrtp_1
X_3484_ _3529_/CLK _3484_/D vssd1 vssd1 vccd1 vccd1 _3484_/Q sky130_fd_sc_hd__dfxtp_1
X_2504_ _3329_/Q _2493_/X _2503_/X _2501_/X vssd1 vssd1 vccd1 vccd1 _3329_/D sky130_fd_sc_hd__o211a_1
XFILLER_69_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2435_ _2563_/A _2441_/B vssd1 vssd1 vccd1 vccd1 _2435_/X sky130_fd_sc_hd__or2_1
XANTENNA__3142__A2 _3160_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2366_ _2366_/A vssd1 vssd1 vccd1 vccd1 _2366_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2756__A _2756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1660__A _2037_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2297_ _2297_/A _2297_/B vssd1 vssd1 vccd1 vccd1 _2353_/A sky130_fd_sc_hd__nand2_1
XFILLER_84_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2491__A _2568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrlbp_macro_334 vssd1 vssd1 vccd1 vccd1 rlbp_macro_334/HI wbs_dat_o[20] sky130_fd_sc_hd__conb_1
Xrlbp_macro_301 vssd1 vssd1 vccd1 vccd1 rlbp_macro_301/HI la_data_out[103] sky130_fd_sc_hd__conb_1
Xrlbp_macro_312 vssd1 vssd1 vccd1 vccd1 rlbp_macro_312/HI la_data_out[114] sky130_fd_sc_hd__conb_1
Xrlbp_macro_323 vssd1 vssd1 vccd1 vccd1 rlbp_macro_323/HI la_data_out[125] sky130_fd_sc_hd__conb_1
Xrlbp_macro_345 vssd1 vssd1 vccd1 vccd1 rlbp_macro_345/HI wbs_dat_o[31] sky130_fd_sc_hd__conb_1
XFILLER_75_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2666__A _2778_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3109__C1 _3108_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2220_ _2216_/Y _2191_/B _2389_/A _2219_/Y vssd1 vssd1 vccd1 vccd1 _2220_/X sky130_fd_sc_hd__o211a_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2151_ _2151_/A _2151_/B vssd1 vssd1 vccd1 vccd1 _2168_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__2576__A _2576_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2082_ _3334_/Q _2073_/Y _2076_/Y _2079_/Y _2081_/Y vssd1 vssd1 vccd1 vccd1 _2083_/D
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_66_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2295__B _2295_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2984_ _3041_/A _3021_/A _3017_/A _3024_/A vssd1 vssd1 vccd1 vccd1 _2985_/D sky130_fd_sc_hd__or4_1
X_1935_ _3303_/Q vssd1 vssd1 vccd1 vccd1 _2288_/B sky130_fd_sc_hd__buf_2
XFILLER_21_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3200__A _3251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1866_ _3428_/Q _2042_/B vssd1 vssd1 vccd1 vccd1 _1926_/B sky130_fd_sc_hd__xnor2_2
Xinput61 wbs_dat_i[7] vssd1 vssd1 vccd1 vccd1 _3243_/A sky130_fd_sc_hd__clkbuf_4
Xinput50 wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 _2982_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__1655__A _1932_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1797_ _3446_/Q _1796_/X vssd1 vssd1 vccd1 vccd1 _1797_/X sky130_fd_sc_hd__or2b_1
X_3536_ _3536_/D _2358_/X vssd1 vssd1 vccd1 vccd1 _3538_/D sky130_fd_sc_hd__dlxtn_1
X_3467_ _3469_/CLK _3467_/D vssd1 vssd1 vccd1 vccd1 _3467_/Q sky130_fd_sc_hd__dfxtp_2
X_3398_ _3400_/CLK _3398_/D vssd1 vssd1 vccd1 vccd1 _3398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2418_ _2552_/A _2983_/A vssd1 vssd1 vccd1 vccd1 _2427_/A sky130_fd_sc_hd__or2_2
XFILLER_84_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2486__A _2563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2349_ _2340_/Y _2341_/X _2344_/Y _2345_/X _2348_/Y vssd1 vssd1 vccd1 vccd1 _2352_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_29_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2626__A1 _3365_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3051__A1 _3360_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3051__B2 _3456_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3780__A _3780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrlbp_macro_142 vssd1 vssd1 vccd1 vccd1 rlbp_macro_142/HI io_oeb[9] sky130_fd_sc_hd__conb_1
Xrlbp_macro_175 vssd1 vssd1 vccd1 vccd1 rlbp_macro_175/HI io_out[4] sky130_fd_sc_hd__conb_1
Xrlbp_macro_164 vssd1 vssd1 vccd1 vccd1 rlbp_macro_164/HI io_oeb[31] sky130_fd_sc_hd__conb_1
Xrlbp_macro_153 vssd1 vssd1 vccd1 vccd1 rlbp_macro_153/HI io_oeb[20] sky130_fd_sc_hd__conb_1
XFILLER_0_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrlbp_macro_197 vssd1 vssd1 vccd1 vccd1 rlbp_macro_197/HI irq[2] sky130_fd_sc_hd__conb_1
XFILLER_0_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input33_A la_data_in[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrlbp_macro_186 vssd1 vssd1 vccd1 vccd1 rlbp_macro_186/HI io_out[15] sky130_fd_sc_hd__conb_1
XFILLER_75_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_538 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3290__A1 hold2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1720_ _3495_/Q _1645_/Y _1648_/Y _3493_/Q vssd1 vssd1 vccd1 vccd1 _1720_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_7_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1651_ _3219_/A _3307_/Q _2405_/B _3210_/A vssd1 vssd1 vccd1 vccd1 _1651_/X sky130_fd_sc_hd__a22o_1
XFILLER_98_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3321_ _3322_/CLK _3321_/D vssd1 vssd1 vccd1 vccd1 _3321_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3252_ _3522_/Q _3256_/B _3256_/C vssd1 vssd1 vccd1 vccd1 _3252_/X sky130_fd_sc_hd__or3_1
XFILLER_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2203_ _2201_/X _2203_/B vssd1 vssd1 vccd1 vccd1 _2238_/B sky130_fd_sc_hd__and2b_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2856__A1 _3434_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3183_ _3183_/A _3183_/B vssd1 vssd1 vccd1 vccd1 _3183_/X sky130_fd_sc_hd__or2_1
XFILLER_78_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2134_ _2134_/A _2134_/B vssd1 vssd1 vccd1 vccd1 _2135_/A sky130_fd_sc_hd__and2_1
XFILLER_54_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2608__A1 _3360_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2065_ _2084_/A _2084_/B _2030_/A vssd1 vssd1 vccd1 vccd1 _2067_/A sky130_fd_sc_hd__a21o_1
XFILLER_54_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2967_ _3471_/Q _2962_/X _2966_/X _2958_/X vssd1 vssd1 vccd1 vccd1 _3471_/D sky130_fd_sc_hd__o211a_1
X_1918_ _3412_/Q _1918_/B vssd1 vssd1 vccd1 vccd1 _1919_/B sky130_fd_sc_hd__xnor2_1
X_2898_ _3449_/Q _2888_/X _2897_/X _2895_/X vssd1 vssd1 vccd1 vccd1 _3449_/D sky130_fd_sc_hd__o211a_1
Xclkbuf_2_3__f_net107 clkbuf_0_net107/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3__f_net107/X
+ sky130_fd_sc_hd__clkbuf_16
X_1849_ _3425_/Q _2118_/B vssd1 vssd1 vccd1 vccd1 _1851_/A sky130_fd_sc_hd__nor2_1
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3519_ _3520_/CLK _3519_/D vssd1 vssd1 vccd1 vccd1 _3527_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2847__A1 _3431_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_368 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2075__A2 _2074_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_435 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1939__A_N _3304_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3263__A1 _3528_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3015__A1 _3358_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3015__B2 _3454_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2821_ _2970_/A _2824_/B vssd1 vssd1 vccd1 vccd1 _2821_/X sky130_fd_sc_hd__or2_1
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2752_ _2788_/A _2754_/B vssd1 vssd1 vccd1 vccd1 _2767_/A sky130_fd_sc_hd__and2_1
X_1703_ _3512_/Q _2294_/B vssd1 vssd1 vccd1 vccd1 _1703_/X sky130_fd_sc_hd__xor2_1
X_2683_ _2758_/A _2690_/B vssd1 vssd1 vccd1 vccd1 _2683_/X sky130_fd_sc_hd__or2_1
XANTENNA__1713__A1_N _3497_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1933__A _3319_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3304_ _3445_/CLK _3304_/D vssd1 vssd1 vccd1 vccd1 _3304_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3235_ _3524_/Q _3224_/X _3234_/X _3228_/X vssd1 vssd1 vccd1 vccd1 _3516_/D sky130_fd_sc_hd__o211a_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_39_net107_A _3494_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3166_ _3232_/A _3170_/B vssd1 vssd1 vccd1 vccd1 _3166_/X sky130_fd_sc_hd__or2_1
XFILLER_39_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2117_ _2117_/A _2117_/B vssd1 vssd1 vccd1 vccd1 _2185_/A sky130_fd_sc_hd__nor2_1
XFILLER_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3097_ _3121_/A _3097_/B vssd1 vssd1 vccd1 vccd1 _3097_/X sky130_fd_sc_hd__or2_1
XFILLER_39_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2048_ _2048_/A _2048_/B _2100_/B _2048_/D vssd1 vssd1 vccd1 vccd1 _2049_/B sky130_fd_sc_hd__nand4_2
XFILLER_22_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_287 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_6 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2674__A _3006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2220__A2 _2191_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3020_ _3442_/Q _3017_/X _3018_/X _3490_/Q _3019_/X vssd1 vssd1 vccd1 vccd1 _3027_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_63_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2584__A _2584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_198 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2804_ _3420_/Q _2789_/X _2803_/X _2797_/X vssd1 vssd1 vccd1 vccd1 _3420_/D sky130_fd_sc_hd__o211a_1
X_3784_ _3784_/A vssd1 vssd1 vccd1 vccd1 _3784_/X sky130_fd_sc_hd__clkbuf_1
X_2735_ _2773_/A _2739_/B vssd1 vssd1 vccd1 vccd1 _2735_/X sky130_fd_sc_hd__or2_1
X_2666_ _2778_/A _2666_/B vssd1 vssd1 vccd1 vccd1 _2666_/X sky130_fd_sc_hd__or2_1
XFILLER_99_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2597_ _2756_/A _2610_/B vssd1 vssd1 vccd1 vccd1 _2597_/X sky130_fd_sc_hd__or2_1
XFILLER_99_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3218_ _2582_/A _3207_/X _3217_/X _3213_/X vssd1 vssd1 vccd1 vccd1 _3510_/D sky130_fd_sc_hd__o211a_1
XFILLER_54_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3149_ _3368_/Q _3036_/A _3037_/A _3464_/Q vssd1 vssd1 vccd1 vccd1 _3149_/X sky130_fd_sc_hd__a22o_1
XFILLER_39_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_368 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_18 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1838__A _3439_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_268 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_55 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_368 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3218__A1 _2582_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2520_ _2679_/A _2520_/B vssd1 vssd1 vccd1 vccd1 _2549_/B sky130_fd_sc_hd__nand2_1
XFILLER_60_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2579__A _2742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2451_ _3241_/A vssd1 vssd1 vccd1 vccd1 _2574_/A sky130_fd_sc_hd__clkbuf_2
X_2382_ _2387_/C vssd1 vssd1 vccd1 vccd1 _2397_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_96_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput4 io_in[17] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_2
X_3003_ _3042_/A vssd1 vssd1 vccd1 vccd1 _3056_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_51_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3209__A1 _2572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1658__A _3304_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2718_ _2731_/A vssd1 vssd1 vccd1 vccd1 _2718_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2649_ _2760_/A _2653_/B vssd1 vssd1 vccd1 vccd1 _2649_/X sky130_fd_sc_hd__or2_1
XANTENNA__2489__A _2565_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1840__B _1840_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3783__A _3783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input63_A wbs_dat_i[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_227 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1750__B _2025_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_488 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1951_ _3311_/Q _3299_/Q vssd1 vssd1 vccd1 vccd1 _1999_/A sky130_fd_sc_hd__xnor2_1
X_1882_ _1876_/Y _1698_/A _1881_/X vssd1 vssd1 vccd1 vccd1 _1882_/X sky130_fd_sc_hd__o21a_1
XFILLER_14_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3552_ _3552_/D _2364_/X vssd1 vssd1 vccd1 vccd1 _3554_/D sky130_fd_sc_hd__dlxtn_1
XFILLER_6_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2503_ _2578_/A _2505_/B vssd1 vssd1 vccd1 vccd1 _2503_/X sky130_fd_sc_hd__or2_1
X_3483_ _3529_/CLK _3483_/D vssd1 vssd1 vccd1 vccd1 _3483_/Q sky130_fd_sc_hd__dfxtp_1
X_2434_ _3232_/A vssd1 vssd1 vccd1 vccd1 _2563_/A sky130_fd_sc_hd__buf_2
X_2365_ _3559_/Q _3558_/Q vssd1 vssd1 vccd1 vccd1 _2366_/A sky130_fd_sc_hd__and2_1
XFILLER_69_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2296_ _2296_/A _2350_/A _2317_/B _2330_/C vssd1 vssd1 vccd1 vccd1 _2297_/B sky130_fd_sc_hd__and4_1
XFILLER_84_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_260 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_455 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_308 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrlbp_macro_324 vssd1 vssd1 vccd1 vccd1 rlbp_macro_324/HI la_data_out[126] sky130_fd_sc_hd__conb_1
Xrlbp_macro_302 vssd1 vssd1 vccd1 vccd1 rlbp_macro_302/HI la_data_out[104] sky130_fd_sc_hd__conb_1
Xrlbp_macro_313 vssd1 vssd1 vccd1 vccd1 rlbp_macro_313/HI la_data_out[115] sky130_fd_sc_hd__conb_1
XANTENNA__2012__A _3327_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrlbp_macro_335 vssd1 vssd1 vccd1 vccd1 rlbp_macro_335/HI wbs_dat_o[21] sky130_fd_sc_hd__conb_1
XANTENNA__2947__A _3158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3778__A _3778_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2857__A _2966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2332__A1 _3454_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2150_ _3378_/Q _2150_/B vssd1 vssd1 vccd1 vccd1 _2151_/B sky130_fd_sc_hd__xnor2_1
XFILLER_38_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2081_ _3335_/Q _2081_/B vssd1 vssd1 vccd1 vccd1 _2081_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_66_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2592__A _3223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2983_ _2983_/A _2983_/B vssd1 vssd1 vccd1 vccd1 _3024_/A sky130_fd_sc_hd__nor2_2
XFILLER_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1934_ _1934_/A _1934_/B vssd1 vssd1 vccd1 vccd1 _1983_/A sky130_fd_sc_hd__nand2_1
X_1865_ _1865_/A _1918_/B _1914_/A vssd1 vssd1 vccd1 vccd1 _1873_/B sky130_fd_sc_hd__and3_1
Xinput40 wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 _2512_/A sky130_fd_sc_hd__clkbuf_1
X_1796_ _2282_/B vssd1 vssd1 vccd1 vccd1 _1796_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput51 wbs_cyc_i vssd1 vssd1 vccd1 vccd1 _2420_/B sky130_fd_sc_hd__clkbuf_1
Xinput62 wbs_dat_i[8] vssd1 vssd1 vccd1 vccd1 _3181_/A sky130_fd_sc_hd__buf_2
X_3535_ _3535_/D _2358_/X vssd1 vssd1 vccd1 vccd1 _3535_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3466_ _3469_/CLK _3466_/D vssd1 vssd1 vccd1 vccd1 _3466_/Q sky130_fd_sc_hd__dfxtp_1
X_2417_ _2512_/A _2512_/B _2512_/C _2511_/A vssd1 vssd1 vccd1 vccd1 _2983_/A sky130_fd_sc_hd__or4_4
X_3397_ _3400_/CLK _3397_/D vssd1 vssd1 vccd1 vccd1 _3397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2348_ _2348_/A _2348_/B vssd1 vssd1 vccd1 vccd1 _2348_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_29_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2279_ _2335_/A _2327_/B vssd1 vssd1 vccd1 vccd1 _2280_/D sky130_fd_sc_hd__and2_1
XFILLER_83_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_182 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2562__A1 _3346_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2677__A _2788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrlbp_macro_176 vssd1 vssd1 vccd1 vccd1 rlbp_macro_176/HI io_out[5] sky130_fd_sc_hd__conb_1
Xrlbp_macro_154 vssd1 vssd1 vccd1 vccd1 rlbp_macro_154/HI io_oeb[21] sky130_fd_sc_hd__conb_1
Xrlbp_macro_143 vssd1 vssd1 vccd1 vccd1 rlbp_macro_143/HI io_oeb[10] sky130_fd_sc_hd__conb_1
Xrlbp_macro_165 vssd1 vssd1 vccd1 vccd1 rlbp_macro_165/HI io_oeb[32] sky130_fd_sc_hd__conb_1
XFILLER_0_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrlbp_macro_198 vssd1 vssd1 vccd1 vccd1 rlbp_macro_198/HI la_data_out[0] sky130_fd_sc_hd__conb_1
Xrlbp_macro_187 vssd1 vssd1 vccd1 vccd1 rlbp_macro_187/HI io_out[16] sky130_fd_sc_hd__conb_1
XFILLER_87_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input26_A la_data_in[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3290__A2 _3281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1650_ _3507_/Q vssd1 vssd1 vccd1 vccd1 _3210_/A sky130_fd_sc_hd__inv_2
XFILLER_7_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2002__B1 _3322_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3320_ _3322_/CLK _3320_/D vssd1 vssd1 vccd1 vccd1 _3320_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3251_ _3251_/A vssd1 vssd1 vccd1 vccd1 _3251_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2202_ _3398_/Q _2282_/B vssd1 vssd1 vccd1 vccd1 _2203_/B sky130_fd_sc_hd__or2b_1
XFILLER_21_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3182_ _3497_/Q _3173_/X _3181_/X _3171_/X vssd1 vssd1 vccd1 vccd1 _3497_/D sky130_fd_sc_hd__o211a_1
X_2133_ _3550_/D _2133_/B _2185_/A _2133_/D vssd1 vssd1 vccd1 vccd1 _2134_/B sky130_fd_sc_hd__nand4_1
XFILLER_66_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2064_ _2048_/B _2068_/B _2058_/X _2063_/X vssd1 vssd1 vccd1 vccd1 _2084_/B sky130_fd_sc_hd__a211o_1
XFILLER_81_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2966_ _2966_/A _2973_/B vssd1 vssd1 vccd1 vccd1 _2966_/X sky130_fd_sc_hd__or2_1
XANTENNA__1666__A _2025_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1917_ _1914_/A _1914_/B _1864_/B vssd1 vssd1 vccd1 vccd1 _1919_/A sky130_fd_sc_hd__a21oi_1
X_2897_ _2970_/A _2899_/B vssd1 vssd1 vccd1 vccd1 _2897_/X sky130_fd_sc_hd__or2_1
X_1848_ _2389_/C _3417_/Q vssd1 vssd1 vccd1 vccd1 _1901_/B sky130_fd_sc_hd__nand2b_1
X_1779_ _3451_/Q _2292_/B vssd1 vssd1 vccd1 vccd1 _1780_/B sky130_fd_sc_hd__and2_1
XFILLER_89_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3518_ _3520_/CLK _3518_/D vssd1 vssd1 vccd1 vccd1 _3526_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2497__A _2574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3449_ _3452_/CLK _3449_/D vssd1 vssd1 vccd1 vccd1 _3449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2960__A _2960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3791__A _3791_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2200__A _3397_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2870__A _3002_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3015__A2 _2595_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2820_ _3181_/A vssd1 vssd1 vccd1 vccd1 _2970_/A sky130_fd_sc_hd__clkbuf_2
X_2751_ _2751_/A vssd1 vssd1 vccd1 vccd1 _2754_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_2682_ _3381_/Q _2678_/X _2681_/X _2668_/X vssd1 vssd1 vccd1 vccd1 _3381_/D sky130_fd_sc_hd__o211a_1
XANTENNA__2774__A1 _3412_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1702_ _3308_/Q vssd1 vssd1 vccd1 vccd1 _2294_/B sky130_fd_sc_hd__buf_4
XFILLER_98_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_255 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3303_ _3307_/CLK _3303_/D vssd1 vssd1 vccd1 vccd1 _3303_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1933__B _2115_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3234_ _3234_/A _3236_/B vssd1 vssd1 vccd1 vccd1 _3234_/X sky130_fd_sc_hd__or2_1
XFILLER_58_119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3165_ _3490_/Q _3159_/X _3164_/X _3156_/X vssd1 vssd1 vccd1 vccd1 _3490_/D sky130_fd_sc_hd__o211a_1
X_2116_ _3367_/Q _2292_/B vssd1 vssd1 vccd1 vccd1 _2117_/B sky130_fd_sc_hd__and2_1
XFILLER_54_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3096_ _3315_/Q _2993_/X _3088_/X _3095_/X vssd1 vssd1 vccd1 vccd1 _3097_/B sky130_fd_sc_hd__a211o_1
X_2047_ _3549_/Q _3548_/Q _2097_/A _2074_/C vssd1 vssd1 vccd1 vccd1 _2048_/D sky130_fd_sc_hd__and4b_1
XFILLER_81_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2780__A _2780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2214__B1 _2213_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_428 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2949_ _3160_/A _2949_/B vssd1 vssd1 vccd1 vccd1 _2977_/B sky130_fd_sc_hd__nand2_1
XFILLER_13_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2955__A _2955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2674__B _2709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3786__A input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2690__A _2765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2508__A1 _3331_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1731__A2 _2373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_450 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2803_ _2957_/A _2806_/B vssd1 vssd1 vccd1 vccd1 _2803_/X sky130_fd_sc_hd__or2_1
X_3783_ _3783_/A vssd1 vssd1 vccd1 vccd1 _3783_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2105__A _3361_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2734_ _3399_/Q _2728_/X _2733_/X _2731_/X vssd1 vssd1 vccd1 vccd1 _3399_/D sky130_fd_sc_hd__o211a_1
X_2665_ _3377_/Q _2656_/X _2664_/X _2654_/X vssd1 vssd1 vccd1 vccd1 _3377_/D sky130_fd_sc_hd__o211a_1
X_2596_ _2634_/B vssd1 vssd1 vccd1 vccd1 _2610_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__1970__A2 _1698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2775__A _2775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3217_ _3510_/Q _3221_/B vssd1 vssd1 vccd1 vccd1 _3217_/X sky130_fd_sc_hd__or2_1
X_3148_ _3404_/Q _2711_/A _2750_/A _3416_/Q vssd1 vssd1 vccd1 vccd1 _3153_/B sky130_fd_sc_hd__a22o_1
XFILLER_94_291 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3079_ _3446_/Q _2872_/A _3008_/A _3494_/Q vssd1 vssd1 vccd1 vccd1 _3079_/X sky130_fd_sc_hd__a22o_1
XFILLER_42_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2015__A _3328_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3163__A1 _3489_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2685__A _2760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_opt_1_0_net107 clkbuf_leaf_9_net107/A vssd1 vssd1 vccd1 vccd1 clkbuf_opt_1_0_net107/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_81_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1764__A _3445_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2450_ _3314_/Q _2446_/X _2449_/X _2444_/X vssd1 vssd1 vccd1 vccd1 _3314_/D sky130_fd_sc_hd__o211a_1
XFILLER_96_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2381_ _3808_/A _2381_/B vssd1 vssd1 vccd1 vccd1 _2387_/C sky130_fd_sc_hd__nor2_1
XANTENNA__1704__A2 _2395_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2595__A _2679_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput5 la_data_in[0] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__buf_2
X_3002_ _3002_/A _3006_/B vssd1 vssd1 vccd1 vccd1 _3042_/A sky130_fd_sc_hd__nor2_1
XFILLER_64_442 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2717_ _2756_/A _2726_/B vssd1 vssd1 vccd1 vccd1 _2717_/X sky130_fd_sc_hd__or2_1
XFILLER_10_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2648_ _3370_/Q _2642_/X _2647_/X _2635_/X vssd1 vssd1 vccd1 vccd1 _3370_/D sky130_fd_sc_hd__o211a_1
XFILLER_10_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3145__A1 _3332_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2579_ _2742_/A vssd1 vssd1 vccd1 vccd1 _2654_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_59_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_23_net107_A _3436_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_272 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3136__A1 _3331_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input56_A wbs_dat_i[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3136__B2 _3451_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1950_ _2001_/A _2001_/B vssd1 vssd1 vccd1 vccd1 _2003_/B sky130_fd_sc_hd__nand2_1
X_1881_ _3419_/Q _2190_/B vssd1 vssd1 vccd1 vccd1 _1881_/X sky130_fd_sc_hd__and2b_1
X_3551_ _3551_/D _2364_/X vssd1 vssd1 vccd1 vccd1 _3553_/D sky130_fd_sc_hd__dlxtn_1
XANTENNA__2583__C1 _2580_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2502_ _3328_/Q _2493_/X _2499_/X _2501_/X vssd1 vssd1 vccd1 vccd1 _3328_/D sky130_fd_sc_hd__o211a_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3482_ _3529_/CLK _3482_/D vssd1 vssd1 vccd1 vccd1 _3482_/Q sky130_fd_sc_hd__dfxtp_1
X_2433_ _3310_/Q _2425_/X _2432_/X _2370_/X vssd1 vssd1 vccd1 vccd1 _3310_/D sky130_fd_sc_hd__o211a_1
X_2364_ _2364_/A vssd1 vssd1 vccd1 vccd1 _2364_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1774__A_N _3447_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2295_ _3465_/Q _2295_/B vssd1 vssd1 vccd1 vccd1 _2330_/C sky130_fd_sc_hd__or2_1
XFILLER_25_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_486 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1669__A _3509_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrlbp_macro_325 vssd1 vssd1 vccd1 vccd1 rlbp_macro_325/HI la_data_out[127] sky130_fd_sc_hd__conb_1
Xrlbp_macro_303 vssd1 vssd1 vccd1 vccd1 rlbp_macro_303/HI la_data_out[105] sky130_fd_sc_hd__conb_1
Xrlbp_macro_314 vssd1 vssd1 vccd1 vccd1 rlbp_macro_314/HI la_data_out[116] sky130_fd_sc_hd__conb_1
XFILLER_99_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrlbp_macro_336 vssd1 vssd1 vccd1 vccd1 rlbp_macro_336/HI wbs_dat_o[22] sky130_fd_sc_hd__conb_1
XFILLER_101_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_320 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_180 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3794__A _3794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_368 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3109__A1 _3316_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2080_ _2080_/A _2080_/B vssd1 vssd1 vccd1 vccd1 _2081_/B sky130_fd_sc_hd__xor2_1
XFILLER_81_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2873__A _3158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2592__B _2595_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2982_ _2982_/A _2982_/B _2982_/C _2905_/B vssd1 vssd1 vccd1 vccd1 _2983_/B sky130_fd_sc_hd__or4b_1
X_1933_ _3319_/Q _2115_/B vssd1 vssd1 vccd1 vccd1 _1934_/B sky130_fd_sc_hd__nand2_1
X_1864_ _1864_/A _1864_/B vssd1 vssd1 vccd1 vccd1 _1914_/A sky130_fd_sc_hd__nor2_1
Xinput30 la_data_in[33] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__1936__B _2288_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput41 wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 _2419_/D sky130_fd_sc_hd__clkbuf_1
Xinput63 wbs_dat_i[9] vssd1 vssd1 vccd1 vccd1 _3183_/A sky130_fd_sc_hd__clkbuf_2
Xinput52 wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 _3227_/A sky130_fd_sc_hd__clkbuf_4
X_1795_ _3445_/Q _1794_/X vssd1 vssd1 vccd1 vccd1 _1795_/X sky130_fd_sc_hd__or2b_1
X_3534_ _1748_/A0 _3534_/D vssd1 vssd1 vccd1 vccd1 _3534_/Q sky130_fd_sc_hd__dfxtp_1
X_3465_ _3469_/CLK _3465_/D vssd1 vssd1 vccd1 vccd1 _3465_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2416_ _2982_/A _2982_/B _2982_/C _2905_/B vssd1 vssd1 vccd1 vccd1 _2552_/A sky130_fd_sc_hd__or4_2
X_3396_ _3396_/CLK _3396_/D vssd1 vssd1 vccd1 vccd1 _3396_/Q sky130_fd_sc_hd__dfxtp_2
X_2347_ _3460_/Q _2347_/B vssd1 vssd1 vccd1 vccd1 _2348_/B sky130_fd_sc_hd__xnor2_1
XFILLER_69_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2278_ _3468_/Q _3300_/Q vssd1 vssd1 vccd1 vccd1 _2327_/B sky130_fd_sc_hd__xnor2_1
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2023__A _3346_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrlbp_macro_133 vssd1 vssd1 vccd1 vccd1 rlbp_macro_133/HI io_oeb[0] sky130_fd_sc_hd__conb_1
XANTENNA__2677__B _2679_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrlbp_macro_166 vssd1 vssd1 vccd1 vccd1 rlbp_macro_166/HI io_oeb[33] sky130_fd_sc_hd__conb_1
Xrlbp_macro_144 vssd1 vssd1 vccd1 vccd1 rlbp_macro_144/HI io_oeb[11] sky130_fd_sc_hd__conb_1
Xrlbp_macro_155 vssd1 vssd1 vccd1 vccd1 rlbp_macro_155/HI io_oeb[22] sky130_fd_sc_hd__conb_1
XANTENNA__2314__A2 _1922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrlbp_macro_199 vssd1 vssd1 vccd1 vccd1 rlbp_macro_199/HI la_data_out[1] sky130_fd_sc_hd__conb_1
Xrlbp_macro_177 vssd1 vssd1 vccd1 vccd1 rlbp_macro_177/HI io_out[6] sky130_fd_sc_hd__conb_1
Xrlbp_macro_188 vssd1 vssd1 vccd1 vccd1 rlbp_macro_188/HI io_out[17] sky130_fd_sc_hd__conb_1
XFILLER_0_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3789__A _3789_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input19_A la_data_in[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1756__B _2313_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2868__A _2977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3250_ _3522_/Q _3253_/A2 _3239_/X _3249_/X vssd1 vssd1 vccd1 vccd1 _3522_/D sky130_fd_sc_hd__o211a_1
XFILLER_3_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2201_ _2282_/B _3398_/Q vssd1 vssd1 vccd1 vccd1 _2201_/X sky130_fd_sc_hd__and2b_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3181_ _3181_/A _3183_/B vssd1 vssd1 vccd1 vccd1 _3181_/X sky130_fd_sc_hd__or2_1
X_2132_ _2132_/A _2163_/A _2165_/B _2132_/D vssd1 vssd1 vccd1 vccd1 _2133_/D sky130_fd_sc_hd__and4_1
XFILLER_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2063_ _2091_/B _2087_/A _2062_/Y _2405_/A _2057_/Y vssd1 vssd1 vccd1 vccd1 _2063_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_19_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2965_ _3470_/Q _2962_/X _2964_/X _2958_/X vssd1 vssd1 vccd1 vccd1 _3470_/D sky130_fd_sc_hd__o211a_1
X_1916_ _3411_/Q _1916_/B vssd1 vssd1 vccd1 vccd1 _1920_/C sky130_fd_sc_hd__nand2_1
X_2896_ _3448_/Q _2888_/X _2894_/X _2895_/X vssd1 vssd1 vccd1 vccd1 _3448_/D sky130_fd_sc_hd__o211a_1
X_1847_ _3418_/Q _2052_/B vssd1 vssd1 vccd1 vccd1 _1900_/A sky130_fd_sc_hd__xnor2_1
X_3517_ _3528_/CLK _3517_/D vssd1 vssd1 vccd1 vccd1 _3525_/Q sky130_fd_sc_hd__dfxtp_1
X_1778_ _1932_/B vssd1 vssd1 vccd1 vccd1 _2292_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__2778__A _2778_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3448_ _3452_/CLK _3448_/D vssd1 vssd1 vccd1 vccd1 _3448_/Q sky130_fd_sc_hd__dfxtp_1
X_3379_ _3392_/CLK _3379_/D vssd1 vssd1 vccd1 vccd1 _3379_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3009__B1 _3160_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2688__A _2762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2200__B _2395_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_29_net107 _3436_/CLK vssd1 vssd1 vccd1 vccd1 _3440_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2750_ _2750_/A vssd1 vssd1 vccd1 vccd1 _2751_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2681_ _2756_/A _2690_/B vssd1 vssd1 vccd1 vccd1 _2681_/X sky130_fd_sc_hd__or2_1
X_1701_ _3501_/Q vssd1 vssd1 vccd1 vccd1 _3193_/A sky130_fd_sc_hd__inv_2
X_3302_ _3307_/CLK _3302_/D vssd1 vssd1 vccd1 vccd1 _3302_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_267 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3233_ _3523_/Q _3224_/X _3232_/X _3228_/X vssd1 vssd1 vccd1 vccd1 _3515_/D sky130_fd_sc_hd__o211a_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3164_ _3230_/A _3170_/B vssd1 vssd1 vccd1 vccd1 _3164_/X sky130_fd_sc_hd__or2_1
XFILLER_39_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_175 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2115_ _3367_/Q _2115_/B vssd1 vssd1 vccd1 vccd1 _2117_/A sky130_fd_sc_hd__nor2_1
XFILLER_54_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3095_ _3095_/A _3095_/B _3095_/C _3095_/D vssd1 vssd1 vccd1 vccd1 _3095_/X sky130_fd_sc_hd__or4_1
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2046_ _3345_/Q _2046_/B vssd1 vssd1 vccd1 vccd1 _2074_/C sky130_fd_sc_hd__or2_1
XFILLER_54_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1677__A _3299_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2948_ _2962_/A vssd1 vssd1 vccd1 vccd1 _2948_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2879_ _2953_/A _2886_/B vssd1 vssd1 vccd1 vccd1 _2879_/X sky130_fd_sc_hd__or2_1
XFILLER_2_606 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1858__A_N _2145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_551 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_0_net107_A _3494_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2453__A1 _3315_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_411 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2211__A _3393_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_410 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2881__A _2955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3782_ _3782_/A vssd1 vssd1 vccd1 vccd1 _3782_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2802_ _3234_/A vssd1 vssd1 vccd1 vccd1 _2957_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_32_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2733_ _2771_/A _2739_/B vssd1 vssd1 vccd1 vccd1 _2733_/X sky130_fd_sc_hd__or2_1
XANTENNA__2105__B _2105_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2664_ _2775_/A _2666_/B vssd1 vssd1 vccd1 vccd1 _2664_/X sky130_fd_sc_hd__or2_1
XFILLER_8_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2595_ _2679_/A _2595_/B vssd1 vssd1 vccd1 vccd1 _2634_/B sky130_fd_sc_hd__nand2_1
XANTENNA__3157__C1 _3156_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3217__A _3510_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_226 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3216_ _2578_/A _3207_/X _3215_/Y _3213_/X vssd1 vssd1 vccd1 vccd1 _3509_/D sky130_fd_sc_hd__o211a_1
X_3147_ _3380_/Q _2997_/X _2679_/B _3392_/Q vssd1 vssd1 vccd1 vccd1 _3153_/A sky130_fd_sc_hd__a22o_1
XFILLER_67_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3078_ _3338_/Q _2516_/A _2997_/X _3374_/Q _3077_/X vssd1 vssd1 vccd1 vccd1 _3083_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_42_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2029_ _3353_/Q _2119_/B vssd1 vssd1 vccd1 vccd1 _2030_/B sky130_fd_sc_hd__and2_1
XANTENNA__2791__A _2875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_12_net107 clkbuf_2_3__f_net107/X vssd1 vssd1 vccd1 vccd1 _3409_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_10_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2031__A _3354_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2966__A _2966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3797__A input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1764__B _2105_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2380_ _2380_/A vssd1 vssd1 vccd1 vccd1 _3296_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2595__B _2595_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2665__A1 _3377_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput6 la_data_in[10] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_2
X_3001_ _3345_/Q _3000_/X _2837_/A _3429_/Q vssd1 vssd1 vccd1 vccd1 _3005_/C sky130_fd_sc_hd__a22o_1
XFILLER_64_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3090__A1 _3339_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1939__B _3316_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3090__B2 _3375_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2716_ _2745_/B vssd1 vssd1 vccd1 vccd1 _2726_/B sky130_fd_sc_hd__clkbuf_1
X_2647_ _2758_/A _2653_/B vssd1 vssd1 vccd1 vccd1 _2647_/X sky130_fd_sc_hd__or2_1
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2578_ _2578_/A _2582_/B vssd1 vssd1 vccd1 vccd1 _2578_/X sky130_fd_sc_hd__or2_1
XFILLER_101_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_295 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1849__B _2118_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3081__A1 _3350_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2026__A _3348_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3081__B2 _3434_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2696__A _2771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input49_A wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1880_ _1900_/A _1901_/B _1879_/X vssd1 vssd1 vccd1 vccd1 _1907_/B sky130_fd_sc_hd__a21o_1
XFILLER_41_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2201__A_N _2282_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3550_ _3550_/D _2364_/X vssd1 vssd1 vccd1 vccd1 _3550_/Q sky130_fd_sc_hd__dlxtn_1
X_2501_ _2566_/A vssd1 vssd1 vccd1 vccd1 _2501_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3481_ _3529_/CLK _3481_/D vssd1 vssd1 vccd1 vccd1 _3481_/Q sky130_fd_sc_hd__dfxtp_1
X_2432_ _2561_/A _2441_/B vssd1 vssd1 vccd1 vccd1 _2432_/X sky130_fd_sc_hd__or2_1
XFILLER_96_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2363_ _3553_/Q _3554_/Q vssd1 vssd1 vccd1 vccd1 _2364_/A sky130_fd_sc_hd__and2_1
XFILLER_69_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2294_ _3476_/Q _2294_/B vssd1 vssd1 vccd1 vccd1 _2317_/B sky130_fd_sc_hd__xnor2_1
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3230__A _3230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrlbp_macro_315 vssd1 vssd1 vccd1 vccd1 rlbp_macro_315/HI la_data_out[117] sky130_fd_sc_hd__conb_1
Xrlbp_macro_304 vssd1 vssd1 vccd1 vccd1 rlbp_macro_304/HI la_data_out[106] sky130_fd_sc_hd__conb_1
Xrlbp_macro_326 vssd1 vssd1 vccd1 vccd1 rlbp_macro_326/HI wbs_dat_o[12] sky130_fd_sc_hd__conb_1
Xrlbp_macro_337 vssd1 vssd1 vccd1 vccd1 rlbp_macro_337/HI wbs_dat_o[23] sky130_fd_sc_hd__conb_1
XFILLER_101_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3054__B2 _3524_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2096__A2 _1834_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2981_ _2981_/A _2996_/A _2981_/C _2981_/D vssd1 vssd1 vccd1 vccd1 _2986_/A sky130_fd_sc_hd__or4_1
XANTENNA__3045__A1 _3467_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1932_ _3319_/Q _1932_/B vssd1 vssd1 vccd1 vccd1 _1934_/A sky130_fd_sc_hd__or2_1
XFILLER_14_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1863_ _3423_/Q _2206_/B vssd1 vssd1 vccd1 vccd1 _1864_/B sky130_fd_sc_hd__and2b_1
Xinput31 la_data_in[3] vssd1 vssd1 vccd1 vccd1 _3789_/A sky130_fd_sc_hd__clkbuf_2
Xinput20 la_data_in[23] vssd1 vssd1 vccd1 vccd1 _3785_/A sky130_fd_sc_hd__clkbuf_2
Xinput42 wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 _2419_/C sky130_fd_sc_hd__clkbuf_1
Xinput64 wbs_sel_i[0] vssd1 vssd1 vccd1 vccd1 _2421_/B sky130_fd_sc_hd__clkbuf_1
Xinput53 wbs_dat_i[10] vssd1 vssd1 vccd1 vccd1 _3186_/A sky130_fd_sc_hd__clkbuf_2
X_1794_ _2281_/B vssd1 vssd1 vccd1 vccd1 _1794_/X sky130_fd_sc_hd__clkbuf_2
X_3533_ _3533_/CLK _3533_/D vssd1 vssd1 vccd1 vccd1 _3533_/Q sky130_fd_sc_hd__dfxtp_1
X_3464_ _3464_/CLK _3464_/D vssd1 vssd1 vccd1 vccd1 _3464_/Q sky130_fd_sc_hd__dfxtp_2
X_2415_ _2042_/B _2412_/X _2414_/Y vssd1 vssd1 vccd1 vccd1 _3308_/D sky130_fd_sc_hd__o21a_1
XANTENNA__1952__B _3300_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3395_ _3396_/CLK _3395_/D vssd1 vssd1 vccd1 vccd1 _3395_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__3225__A _3225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2346_ _2343_/A _2343_/B _2289_/B vssd1 vssd1 vccd1 vccd1 _2348_/A sky130_fd_sc_hd__a21o_1
XFILLER_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2277_ _3467_/Q _3299_/Q vssd1 vssd1 vccd1 vccd1 _2335_/A sky130_fd_sc_hd__xnor2_2
XFILLER_29_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2023__B _2052_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrlbp_macro_167 vssd1 vssd1 vccd1 vccd1 rlbp_macro_167/HI io_oeb[34] sky130_fd_sc_hd__conb_1
Xrlbp_macro_156 vssd1 vssd1 vccd1 vccd1 rlbp_macro_156/HI io_oeb[23] sky130_fd_sc_hd__conb_1
Xrlbp_macro_134 vssd1 vssd1 vccd1 vccd1 rlbp_macro_134/HI io_oeb[1] sky130_fd_sc_hd__conb_1
Xrlbp_macro_145 vssd1 vssd1 vccd1 vccd1 rlbp_macro_145/HI io_oeb[12] sky130_fd_sc_hd__conb_1
XFILLER_0_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrlbp_macro_178 vssd1 vssd1 vccd1 vccd1 rlbp_macro_178/HI io_out[7] sky130_fd_sc_hd__conb_1
Xrlbp_macro_189 vssd1 vssd1 vccd1 vccd1 rlbp_macro_189/HI io_out[18] sky130_fd_sc_hd__conb_1
XFILLER_87_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2200_ _3397_/Q _2395_/A vssd1 vssd1 vccd1 vccd1 _2235_/A sky130_fd_sc_hd__xnor2_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3180_ _3496_/Q _3173_/X _3179_/X _3171_/X vssd1 vssd1 vccd1 vccd1 _3496_/D sky130_fd_sc_hd__o211a_1
X_2131_ _2125_/Y _2183_/B _2159_/B _2161_/A vssd1 vssd1 vccd1 vccd1 _2132_/D sky130_fd_sc_hd__and4bb_1
XANTENNA__2884__A _2957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_527 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2062_ _2059_/X _2060_/X _2061_/X vssd1 vssd1 vccd1 vccd1 _2062_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_19_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2108__B _3364_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2964_ _2964_/A _2973_/B vssd1 vssd1 vccd1 vccd1 _2964_/X sky130_fd_sc_hd__or2_1
X_1915_ _3411_/Q _1916_/B vssd1 vssd1 vccd1 vccd1 _1920_/B sky130_fd_sc_hd__or2_1
X_2895_ _2895_/A vssd1 vssd1 vccd1 vccd1 _2895_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2124__A _2389_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1846_ _1907_/A _1905_/B vssd1 vssd1 vccd1 vccd1 _1854_/A sky130_fd_sc_hd__and2_1
X_1777_ _3451_/Q _2115_/B vssd1 vssd1 vccd1 vccd1 _1780_/A sky130_fd_sc_hd__nor2_1
X_3516_ _3516_/CLK _3516_/D vssd1 vssd1 vccd1 vccd1 _3524_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2138__B_N _2389_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3447_ _3450_/CLK _3447_/D vssd1 vssd1 vccd1 vccd1 _3447_/Q sky130_fd_sc_hd__dfxtp_1
X_3378_ _3392_/CLK _3378_/D vssd1 vssd1 vccd1 vccd1 _3378_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2329_ _2329_/A _2330_/B vssd1 vssd1 vccd1 vccd1 _2329_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_57_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3257__A1 _3525_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_571 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3009__B2 _3489_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2034__A _3349_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input31_A la_data_in[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3248__A1 _3521_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2680_ _2707_/B vssd1 vssd1 vccd1 vccd1 _2690_/B sky130_fd_sc_hd__clkbuf_1
X_1700_ _2389_/C vssd1 vssd1 vccd1 vccd1 _2385_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2879__A _2953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3301_ _3307_/CLK _3301_/D vssd1 vssd1 vccd1 vccd1 _3301_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_279 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3232_ _3232_/A _3236_/B vssd1 vssd1 vccd1 vccd1 _3232_/X sky130_fd_sc_hd__or2_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3163_ _3489_/Q _3159_/X _3162_/X _3156_/X vssd1 vssd1 vccd1 vccd1 _3489_/D sky130_fd_sc_hd__o211a_1
XFILLER_39_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2114_ _2114_/A _2173_/B _2175_/A vssd1 vssd1 vccd1 vccd1 _2133_/B sky130_fd_sc_hd__and3_1
XFILLER_66_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3094_ _3399_/Q _3041_/X _3042_/X _3507_/Q vssd1 vssd1 vccd1 vccd1 _3095_/D sky130_fd_sc_hd__a22o_1
XANTENNA__2119__A _3365_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2045_ _2045_/A _2045_/B vssd1 vssd1 vccd1 vccd1 _2097_/A sky130_fd_sc_hd__nor2_1
XFILLER_54_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2998__B1 _3024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2947_ _3158_/A _2949_/B vssd1 vssd1 vccd1 vccd1 _2962_/A sky130_fd_sc_hd__and2_1
X_2878_ _3441_/Q _2874_/X _2877_/X _2864_/X vssd1 vssd1 vccd1 vccd1 _3441_/D sky130_fd_sc_hd__o211a_1
XANTENNA__1693__A _1693_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1829_ _1824_/A _1824_/B _1775_/B vssd1 vssd1 vccd1 vccd1 _1831_/A sky130_fd_sc_hd__a21oi_1
XFILLER_2_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_17_net107_A clkbuf_2_3__f_net107/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2301__B _2301_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_268 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_35_net107 _3494_/CLK vssd1 vssd1 vccd1 vccd1 _3486_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_38_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2029__A _3353_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_563 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1868__A _3427_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_511 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_566 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_423 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2211__B _2295_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_422 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_308 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1778__A _1932_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3781_ _3781_/A vssd1 vssd1 vccd1 vccd1 _3781_/X sky130_fd_sc_hd__clkbuf_1
X_2801_ _3419_/Q _2789_/X _2800_/X _2797_/X vssd1 vssd1 vccd1 vccd1 _3419_/D sky130_fd_sc_hd__o211a_1
X_2732_ _3398_/Q _2728_/X _2730_/X _2731_/X vssd1 vssd1 vccd1 vccd1 _3398_/D sky130_fd_sc_hd__o211a_1
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2663_ _3376_/Q _2656_/X _2662_/X _2654_/X vssd1 vssd1 vccd1 vccd1 _3376_/D sky130_fd_sc_hd__o211a_1
X_2594_ _3227_/A vssd1 vssd1 vccd1 vccd1 _2756_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__2121__B _2121_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_238 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1960__B _2294_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3215_ _3215_/A _3219_/B vssd1 vssd1 vccd1 vccd1 _3215_/Y sky130_fd_sc_hd__nand2_1
XFILLER_67_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3146_ _3356_/Q _2557_/B _3195_/B _3512_/Q _3145_/X vssd1 vssd1 vccd1 vccd1 _3146_/X
+ sky130_fd_sc_hd__a221o_1
X_3077_ _3386_/Q _2676_/A _3033_/A _3526_/Q vssd1 vssd1 vccd1 vccd1 _3077_/X sky130_fd_sc_hd__a22o_1
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2028_ _3353_/Q _2313_/B vssd1 vssd1 vccd1 vccd1 _2030_/A sky130_fd_sc_hd__nor2_1
XFILLER_82_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1688__A _2389_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2031__B _2121_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1975__A_N _1974_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_466 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2206__B _2206_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2222__A _3400_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3053__A _3053_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput7 la_data_in[11] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_2
X_3000_ _3000_/A vssd1 vssd1 vccd1 vccd1 _3000_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2892__A _2966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3090__A2 _2996_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1848__A_N _2389_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2116__B _2292_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2715_ _2875_/A _2715_/B vssd1 vssd1 vccd1 vccd1 _2745_/B sky130_fd_sc_hd__nand2_1
XANTENNA__1955__B _2119_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2646_ _3369_/Q _2642_/X _2645_/X _2635_/X vssd1 vssd1 vccd1 vccd1 _3369_/D sky130_fd_sc_hd__o211a_1
XANTENNA__3228__A _3251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2577_ _3352_/Q _2570_/X _2576_/X _2566_/X vssd1 vssd1 vccd1 vccd1 _3352_/D sky130_fd_sc_hd__o211a_1
XFILLER_101_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3129_ _3366_/Q _3036_/X _2679_/B _3390_/Q _3128_/X vssd1 vssd1 vccd1 vccd1 _3129_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2026__B _2026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_32_net107_A _3436_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2977__A _2977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2583__A1 _3354_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3480_ _3529_/CLK _3480_/D vssd1 vssd1 vccd1 vccd1 _3480_/Q sky130_fd_sc_hd__dfxtp_1
X_2500_ _2742_/A vssd1 vssd1 vccd1 vccd1 _2566_/A sky130_fd_sc_hd__clkbuf_2
X_2431_ _3230_/A vssd1 vssd1 vccd1 vccd1 _2561_/A sky130_fd_sc_hd__buf_2
X_2362_ _2362_/A vssd1 vssd1 vccd1 vccd1 _2362_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_69_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2293_ _2293_/A _2293_/B vssd1 vssd1 vccd1 vccd1 _2350_/A sky130_fd_sc_hd__nor2_1
XFILLER_96_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1739__B_N _3549_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_491 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2629_ _3366_/Q _2612_/X _2628_/X _2619_/X vssd1 vssd1 vccd1 vccd1 _3366_/D sky130_fd_sc_hd__o211a_1
Xoutput130 _3485_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[8] sky130_fd_sc_hd__buf_2
Xrlbp_macro_305 vssd1 vssd1 vccd1 vccd1 rlbp_macro_305/HI la_data_out[107] sky130_fd_sc_hd__conb_1
Xrlbp_macro_316 vssd1 vssd1 vccd1 vccd1 rlbp_macro_316/HI la_data_out[118] sky130_fd_sc_hd__conb_1
XANTENNA__2326__A1 _3467_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrlbp_macro_338 vssd1 vssd1 vccd1 vccd1 rlbp_macro_338/HI wbs_dat_o[24] sky130_fd_sc_hd__conb_1
Xrlbp_macro_327 vssd1 vssd1 vccd1 vccd1 rlbp_macro_327/HI wbs_dat_o[13] sky130_fd_sc_hd__conb_1
XFILLER_87_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_528 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2037__A _3352_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3054__A2 _3053_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input61_A wbs_dat_i[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2500__A _2742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_591 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2980_ _2551_/B _3006_/A _3006_/B vssd1 vssd1 vccd1 vccd1 _2981_/D sky130_fd_sc_hd__a21oi_1
XFILLER_61_288 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1931_ _1874_/A _1930_/X _1874_/B vssd1 vssd1 vccd1 vccd1 _3537_/D sky130_fd_sc_hd__o21ai_1
XFILLER_14_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1862_ _3303_/Q vssd1 vssd1 vccd1 vccd1 _2206_/B sky130_fd_sc_hd__buf_2
Xinput10 la_data_in[14] vssd1 vssd1 vccd1 vccd1 _3800_/A sky130_fd_sc_hd__clkbuf_2
Xinput21 la_data_in[24] vssd1 vssd1 vccd1 vccd1 _3778_/A sky130_fd_sc_hd__clkbuf_2
Xinput43 wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 _2512_/C sky130_fd_sc_hd__clkbuf_1
Xinput32 la_data_in[4] vssd1 vssd1 vccd1 vccd1 _3790_/A sky130_fd_sc_hd__clkbuf_2
Xinput54 wbs_dat_i[11] vssd1 vssd1 vccd1 vccd1 _3188_/A sky130_fd_sc_hd__buf_2
X_1793_ _1788_/Y _2395_/B _1762_/A _1816_/B _1792_/X vssd1 vssd1 vccd1 vccd1 _1810_/B
+ sky130_fd_sc_hd__a221o_2
Xinput65 wbs_stb_i vssd1 vssd1 vccd1 vccd1 _2420_/A sky130_fd_sc_hd__clkbuf_1
X_3532_ _3533_/CLK _3532_/D vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__dfxtp_1
XFILLER_89_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3463_ _3464_/CLK _3463_/D vssd1 vssd1 vccd1 vccd1 _3463_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_69_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2414_ _2042_/B _2412_/X _2397_/A vssd1 vssd1 vccd1 vccd1 _2414_/Y sky130_fd_sc_hd__a21boi_1
X_3394_ _3396_/CLK _3394_/D vssd1 vssd1 vccd1 vccd1 _3394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2345_ _3459_/Q _2345_/B vssd1 vssd1 vccd1 vccd1 _2345_/X sky130_fd_sc_hd__or2_1
XFILLER_69_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2276_ _1949_/A _3465_/Q vssd1 vssd1 vccd1 vccd1 _2330_/B sky130_fd_sc_hd__nand2b_2
XANTENNA__3241__A _3241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2320__A _3462_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrlbp_macro_146 vssd1 vssd1 vccd1 vccd1 rlbp_macro_146/HI io_oeb[13] sky130_fd_sc_hd__conb_1
Xrlbp_macro_135 vssd1 vssd1 vccd1 vccd1 rlbp_macro_135/HI io_oeb[2] sky130_fd_sc_hd__conb_1
Xrlbp_macro_157 vssd1 vssd1 vccd1 vccd1 rlbp_macro_157/HI io_oeb[24] sky130_fd_sc_hd__conb_1
Xrlbp_macro_168 vssd1 vssd1 vccd1 vccd1 rlbp_macro_168/HI io_oeb[35] sky130_fd_sc_hd__conb_1
Xrlbp_macro_179 vssd1 vssd1 vccd1 vccd1 rlbp_macro_179/HI io_out[8] sky130_fd_sc_hd__conb_1
XFILLER_57_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_340 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2130_ _3359_/Q _2389_/A vssd1 vssd1 vccd1 vccd1 _2161_/A sky130_fd_sc_hd__xnor2_2
XFILLER_78_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_539 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2061_ _1974_/X _3350_/Q vssd1 vssd1 vccd1 vccd1 _2061_/X sky130_fd_sc_hd__and2b_1
XFILLER_54_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_306 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2963_ _2977_/B vssd1 vssd1 vccd1 vccd1 _2973_/B sky130_fd_sc_hd__clkbuf_1
X_1914_ _1914_/A _1914_/B vssd1 vssd1 vccd1 vccd1 _1916_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__2777__A1 _3413_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2894_ _2968_/A _2899_/B vssd1 vssd1 vccd1 vccd1 _2894_/X sky130_fd_sc_hd__or2_1
X_1845_ _3420_/Q _2026_/B vssd1 vssd1 vccd1 vccd1 _1905_/B sky130_fd_sc_hd__xnor2_1
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1776_ _1776_/A _1830_/B _1824_/A vssd1 vssd1 vccd1 vccd1 _1785_/B sky130_fd_sc_hd__and3_1
X_3515_ _3520_/CLK _3515_/D vssd1 vssd1 vccd1 vccd1 _3523_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__3236__A _3236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3446_ _3450_/CLK _3446_/D vssd1 vssd1 vccd1 vccd1 _3446_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_97_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3377_ _3377_/CLK _3377_/D vssd1 vssd1 vccd1 vccd1 _3377_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2328_ _2328_/A _2328_/B vssd1 vssd1 vccd1 vccd1 _2338_/C sky130_fd_sc_hd__xnor2_1
XFILLER_84_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2259_ _3387_/Q _2259_/B vssd1 vssd1 vccd1 vccd1 _2259_/X sky130_fd_sc_hd__or2_1
XFILLER_38_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2034__B _2281_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2940__A1 _3463_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_66 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input24_A la_data_in[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3248__A2 _3253_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2209__B _2292_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2759__A1 _3406_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1982__A2 _1834_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1783__B _2046_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3300_ _3307_/CLK _3300_/D vssd1 vssd1 vccd1 vccd1 _3300_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_98_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3231_ _3522_/Q _3224_/X _3230_/X _3228_/X vssd1 vssd1 vccd1 vccd1 _3514_/D sky130_fd_sc_hd__o211a_1
XFILLER_3_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3162_ _3227_/A _3170_/B vssd1 vssd1 vccd1 vccd1 _3162_/X sky130_fd_sc_hd__or2_1
XFILLER_66_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2113_ _2113_/A _2113_/B vssd1 vssd1 vccd1 vccd1 _2175_/A sky130_fd_sc_hd__nor2_1
XFILLER_39_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3093_ _3351_/Q _3000_/X _3021_/X _3435_/Q vssd1 vssd1 vccd1 vccd1 _3095_/C sky130_fd_sc_hd__a22o_1
XFILLER_81_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2119__B _2119_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2044_ _3355_/Q _2115_/B vssd1 vssd1 vccd1 vccd1 _2045_/B sky130_fd_sc_hd__and2_1
XANTENNA__2998__B2 _3521_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_258 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2946_ _2946_/A vssd1 vssd1 vccd1 vccd1 _2949_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_2877_ _2951_/A _2886_/B vssd1 vssd1 vccd1 vccd1 _2877_/X sky130_fd_sc_hd__or2_1
X_1828_ _3437_/Q _1828_/B vssd1 vssd1 vccd1 vccd1 _1832_/C sky130_fd_sc_hd__xnor2_1
XFILLER_89_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2922__A1 _3456_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1759_ _1759_/A _1759_/B vssd1 vssd1 vccd1 vccd1 _1827_/A sky130_fd_sc_hd__nor2_1
XFILLER_58_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3429_ _3440_/CLK _3429_/D vssd1 vssd1 vccd1 vccd1 _3429_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2029__B _2119_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2989__A1 _2427_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1868__B _2291_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_575 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_578 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_435 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_434 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_531 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3780_ _3780_/A vssd1 vssd1 vccd1 vccd1 _3780_/X sky130_fd_sc_hd__clkbuf_1
X_2800_ _2955_/A _2806_/B vssd1 vssd1 vccd1 vccd1 _2800_/X sky130_fd_sc_hd__or2_1
XFILLER_32_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2731_ _2731_/A vssd1 vssd1 vccd1 vccd1 _2731_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1794__A _2281_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2662_ _2773_/A _2666_/B vssd1 vssd1 vccd1 vccd1 _2662_/X sky130_fd_sc_hd__or2_1
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2593_ _2612_/A vssd1 vssd1 vccd1 vccd1 _2593_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_101_539 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3214_ _2576_/A _3207_/X _3212_/X _3213_/X vssd1 vssd1 vccd1 vccd1 _3508_/D sky130_fd_sc_hd__o211a_1
XFILLER_39_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3145_ _3332_/Q _2477_/A _2946_/A _3476_/Q vssd1 vssd1 vccd1 vccd1 _3145_/X sky130_fd_sc_hd__a22o_1
XFILLER_39_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3076_ _3422_/Q _2787_/A _2949_/B _3470_/Q _3075_/X vssd1 vssd1 vccd1 vccd1 _3076_/X
+ sky130_fd_sc_hd__a221o_1
X_2027_ _2080_/A _2078_/B vssd1 vssd1 vccd1 vccd1 _2033_/C sky130_fd_sc_hd__and2_1
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2929_ _3458_/Q _2925_/X _2927_/X _2928_/X vssd1 vssd1 vccd1 vccd1 _3458_/D sky130_fd_sc_hd__o211a_1
XFILLER_40_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1795__B_N _1794_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_478 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3084__B1 _3076_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2503__A _2578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3139__A1 _3391_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3139__B2 _3475_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput8 la_data_in[12] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2714_ _2834_/A vssd1 vssd1 vccd1 vccd1 _2875_/A sky130_fd_sc_hd__buf_2
X_2645_ _2756_/A _2653_/B vssd1 vssd1 vccd1 vccd1 _2645_/X sky130_fd_sc_hd__or2_1
XFILLER_10_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2576_ _2576_/A _2582_/B vssd1 vssd1 vccd1 vccd1 _2576_/X sky130_fd_sc_hd__or2_1
XFILLER_59_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3128_ _3474_/Q _2945_/A _3018_/X _3498_/Q vssd1 vssd1 vccd1 vccd1 _3128_/X sky130_fd_sc_hd__a22o_1
XFILLER_27_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3059_ _3059_/A _3059_/B _3059_/C _3059_/D vssd1 vssd1 vccd1 vccd1 _3059_/X sky130_fd_sc_hd__or4_2
XFILLER_70_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2042__B _2042_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1881__B _2190_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_294 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2217__B _2301_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2430_ _3309_/Q _2425_/X _2429_/X _2370_/X vssd1 vssd1 vccd1 vccd1 _3309_/D sky130_fd_sc_hd__o211a_1
XANTENNA__1791__B _2190_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2361_ _3549_/Q _3548_/Q vssd1 vssd1 vccd1 vccd1 _2362_/A sky130_fd_sc_hd__and2_1
XFILLER_96_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2292_ _3475_/Q _2292_/B vssd1 vssd1 vccd1 vccd1 _2293_/B sky130_fd_sc_hd__and2_1
XFILLER_96_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2127__B _3360_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3239__A _3251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2628_ _2778_/A _2628_/B vssd1 vssd1 vccd1 vccd1 _2628_/X sky130_fd_sc_hd__or2_1
Xrlbp_macro_306 vssd1 vssd1 vccd1 vccd1 rlbp_macro_306/HI la_data_out[108] sky130_fd_sc_hd__conb_1
Xoutput120 _3477_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[0] sky130_fd_sc_hd__buf_2
Xoutput131 _3486_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[9] sky130_fd_sc_hd__buf_2
XANTENNA__2326__A2 _1678_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2559_ _2559_/A _2568_/B vssd1 vssd1 vccd1 vccd1 _2559_/X sky130_fd_sc_hd__or2_1
Xrlbp_macro_339 vssd1 vssd1 vccd1 vccd1 rlbp_macro_339/HI wbs_dat_o[25] sky130_fd_sc_hd__conb_1
Xrlbp_macro_317 vssd1 vssd1 vccd1 vccd1 rlbp_macro_317/HI la_data_out[119] sky130_fd_sc_hd__conb_1
Xrlbp_macro_328 vssd1 vssd1 vccd1 vccd1 rlbp_macro_328/HI wbs_dat_o[14] sky130_fd_sc_hd__conb_1
XFILLER_99_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2037__B _2037_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_150 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input54_A wbs_dat_i[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_599 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_507 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_212 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1930_ _1910_/X _1930_/B _1930_/C _1930_/D vssd1 vssd1 vccd1 vccd1 _1930_/X sky130_fd_sc_hd__and4b_1
X_1861_ _1774_/B _3423_/Q vssd1 vssd1 vccd1 vccd1 _1864_/A sky130_fd_sc_hd__and2b_1
XFILLER_14_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput22 la_data_in[25] vssd1 vssd1 vccd1 vccd1 _3804_/A sky130_fd_sc_hd__clkbuf_2
Xinput11 la_data_in[15] vssd1 vssd1 vccd1 vccd1 _3801_/A sky130_fd_sc_hd__buf_2
Xinput44 wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 input44/X sky130_fd_sc_hd__clkbuf_1
X_3531_ _3533_/CLK _3531_/D vssd1 vssd1 vccd1 vccd1 _3531_/Q sky130_fd_sc_hd__dfxtp_1
Xinput55 wbs_dat_i[1] vssd1 vssd1 vccd1 vccd1 _3230_/A sky130_fd_sc_hd__clkbuf_4
Xinput33 la_data_in[5] vssd1 vssd1 vccd1 vccd1 _3791_/A sky130_fd_sc_hd__clkbuf_2
X_1792_ _1788_/Y _1698_/A _1791_/X vssd1 vssd1 vccd1 vccd1 _1792_/X sky130_fd_sc_hd__o21a_1
XFILLER_6_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput66 wbs_we_i vssd1 vssd1 vccd1 vccd1 _2421_/A sky130_fd_sc_hd__clkbuf_1
X_3462_ _3462_/CLK _3462_/D vssd1 vssd1 vccd1 vccd1 _3462_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3393_ _3396_/CLK _3393_/D vssd1 vssd1 vccd1 vccd1 _3393_/Q sky130_fd_sc_hd__dfxtp_1
X_2413_ _2291_/B _2410_/Y _2412_/X _3808_/A _2381_/B vssd1 vssd1 vccd1 vccd1 _3307_/D
+ sky130_fd_sc_hd__a2111oi_1
X_2344_ _3459_/Q _2345_/B vssd1 vssd1 vccd1 vccd1 _2344_/Y sky130_fd_sc_hd__nand2_1
XFILLER_96_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2275_ _3466_/Q _2301_/B vssd1 vssd1 vccd1 vccd1 _2329_/A sky130_fd_sc_hd__xnor2_1
XFILLER_84_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2138__A _3359_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2492__A1 _3325_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1977__A _2285_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2143__A_N _1796_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrlbp_macro_158 vssd1 vssd1 vccd1 vccd1 rlbp_macro_158/HI io_oeb[25] sky130_fd_sc_hd__conb_1
Xrlbp_macro_147 vssd1 vssd1 vccd1 vccd1 rlbp_macro_147/HI io_oeb[14] sky130_fd_sc_hd__conb_1
Xrlbp_macro_136 vssd1 vssd1 vccd1 vccd1 rlbp_macro_136/HI io_oeb[3] sky130_fd_sc_hd__conb_1
XFILLER_0_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_18_net107 clkbuf_2_3__f_net107/X vssd1 vssd1 vccd1 vccd1 _3564_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrlbp_macro_169 vssd1 vssd1 vccd1 vccd1 rlbp_macro_169/HI io_oeb[36] sky130_fd_sc_hd__conb_1
XFILLER_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2483__A1 _3321_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_404 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1994__B1 _3321_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2060_ _3350_/Q _1974_/X vssd1 vssd1 vccd1 vccd1 _2060_/X sky130_fd_sc_hd__or2b_1
XFILLER_14_6 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1797__A _3446_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2962_ _2962_/A vssd1 vssd1 vccd1 vccd1 _2962_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1913_ _1865_/A _1895_/B _1887_/Y vssd1 vssd1 vccd1 vccd1 _1914_/B sky130_fd_sc_hd__a21o_1
X_2893_ _3447_/Q _2888_/X _2892_/X _2882_/X vssd1 vssd1 vccd1 vccd1 _3447_/D sky130_fd_sc_hd__o211a_1
X_1844_ _3419_/Q _2025_/B vssd1 vssd1 vccd1 vccd1 _1907_/A sky130_fd_sc_hd__xnor2_1
X_1775_ _1775_/A _1775_/B vssd1 vssd1 vccd1 vccd1 _1824_/A sky130_fd_sc_hd__nor2_1
X_3514_ _3516_/CLK _3514_/D vssd1 vssd1 vccd1 vccd1 _3522_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_89_407 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3445_ _3445_/CLK _3445_/D vssd1 vssd1 vccd1 vccd1 _3445_/Q sky130_fd_sc_hd__dfxtp_2
X_3376_ _3377_/CLK _3376_/D vssd1 vssd1 vccd1 vccd1 _3376_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3252__A _3522_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2327_ _3456_/Q _2327_/B vssd1 vssd1 vccd1 vccd1 _2328_/B sky130_fd_sc_hd__xnor2_1
X_2258_ _3387_/Q _2259_/B vssd1 vssd1 vccd1 vccd1 _2258_/Y sky130_fd_sc_hd__nand2_1
XFILLER_27_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2189_ _3559_/Q _2189_/B vssd1 vssd1 vccd1 vccd1 _2189_/Y sky130_fd_sc_hd__nor2_1
XFILLER_53_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_5_net107 clkbuf_leaf_9_net107/A vssd1 vssd1 vccd1 vccd1 _3512_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2039__A_N _3351_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3162__A _3227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input17_A la_data_in[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2456__A1 _3316_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_554 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2225__B _2288_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3169__C1 _3156_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3230_ _3230_/A _3236_/B vssd1 vssd1 vccd1 vccd1 _3230_/X sky130_fd_sc_hd__or2_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3161_ _3188_/B vssd1 vssd1 vccd1 vccd1 _3170_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_39_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2112_ _3363_/Q _2206_/B vssd1 vssd1 vccd1 vccd1 _2113_/B sky130_fd_sc_hd__and2b_1
XFILLER_12_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3092_ _3327_/Q _2476_/A _2750_/A _3411_/Q _3091_/X vssd1 vssd1 vccd1 vccd1 _3095_/B
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3800__A _3800_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2043_ _3355_/Q _2291_/B vssd1 vssd1 vccd1 vccd1 _2045_/A sky130_fd_sc_hd__nor2_1
XFILLER_47_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2945_ _2945_/A vssd1 vssd1 vccd1 vccd1 _2946_/A sky130_fd_sc_hd__clkbuf_2
X_2876_ _2903_/B vssd1 vssd1 vccd1 vccd1 _2886_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_30_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1827_ _1827_/A _1827_/B vssd1 vssd1 vccd1 vccd1 _1828_/B sky130_fd_sc_hd__xor2_1
X_1758_ _3449_/Q _2119_/B vssd1 vssd1 vccd1 vccd1 _1759_/B sky130_fd_sc_hd__and2_1
X_1689_ _3502_/Q _2385_/A vssd1 vssd1 vccd1 vccd1 _1689_/Y sky130_fd_sc_hd__nand2_1
XFILLER_89_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3428_ _3452_/CLK _3428_/D vssd1 vssd1 vccd1 vccd1 _3428_/Q sky130_fd_sc_hd__dfxtp_1
X_3359_ _3377_/CLK _3359_/D vssd1 vssd1 vccd1 vccd1 _3359_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_58_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input9_A la_data_in[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_148 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_26_net107_A _3436_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_543 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2730_ _2769_/A _2739_/B vssd1 vssd1 vccd1 vccd1 _2730_/X sky130_fd_sc_hd__or2_1
X_2661_ _3375_/Q _2656_/X _2660_/X _2654_/X vssd1 vssd1 vccd1 vccd1 _3375_/D sky130_fd_sc_hd__o211a_1
XFILLER_12_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2592_ _3223_/A _2595_/B vssd1 vssd1 vccd1 vccd1 _2612_/A sky130_fd_sc_hd__and2_1
XFILLER_5_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3213_ _3251_/A vssd1 vssd1 vccd1 vccd1 _3213_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_79_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3144_ _3487_/Q _3074_/A _3143_/X _3098_/X vssd1 vssd1 vccd1 vccd1 _3487_/D sky130_fd_sc_hd__o211a_1
XFILLER_39_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3075_ _3362_/Q _3036_/X _3037_/X _3458_/Q vssd1 vssd1 vccd1 vccd1 _3075_/X sky130_fd_sc_hd__a22o_1
X_2026_ _3348_/Q _2026_/B vssd1 vssd1 vccd1 vccd1 _2078_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__1969__B _2025_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3093__A1 _3351_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3093__B2 _3435_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2928_ _2971_/A vssd1 vssd1 vccd1 vccd1 _2928_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2859_ _2968_/A _2863_/B vssd1 vssd1 vccd1 vccd1 _2859_/X sky130_fd_sc_hd__or2_1
XANTENNA__3148__A2 _2711_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2659__A1 _3374_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1882__A2 _1698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1879__B _2052_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3084__A1 _3314_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_78 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3139__A2 _3053_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput9 la_data_in[13] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__1789__B _2389_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3075__A1 _3362_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2713_ _2728_/A vssd1 vssd1 vccd1 vccd1 _2713_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2644_ _2672_/B vssd1 vssd1 vccd1 vccd1 _2653_/B sky130_fd_sc_hd__clkbuf_1
X_2575_ _3351_/Q _2570_/X _2574_/X _2566_/X vssd1 vssd1 vccd1 vccd1 _3351_/D sky130_fd_sc_hd__o211a_1
XFILLER_87_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_424 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3127_ _3438_/Q _3021_/X _2875_/B _3450_/Q _3126_/X vssd1 vssd1 vccd1 vccd1 _3127_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3260__A _3526_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3066__B2 _3433_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3066__A1 _3349_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3058_ _3396_/Q _2715_/B _3195_/B _3504_/Q _3057_/X vssd1 vssd1 vccd1 vccd1 _3059_/D
+ sky130_fd_sc_hd__a221o_1
X_2009_ _3329_/Q _2009_/B vssd1 vssd1 vccd1 vccd1 _2009_/X sky130_fd_sc_hd__or2_1
XFILLER_35_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2604__A _2760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_26 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3170__A _3236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3057__A1 _3348_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3057__B2 _3432_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_6 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2360_ _2360_/A vssd1 vssd1 vccd1 vccd1 _2360_/X sky130_fd_sc_hd__clkbuf_1
X_2291_ _3475_/Q _2291_/B vssd1 vssd1 vccd1 vccd1 _2293_/A sky130_fd_sc_hd__nor2_1
XFILLER_96_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_287 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_490 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2424__A _2427_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2143__B _3362_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3220__A1 _2584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput110 _3522_/Q vssd1 vssd1 vccd1 vccd1 io_out[24] sky130_fd_sc_hd__buf_2
Xrlbp_macro_307 vssd1 vssd1 vccd1 vccd1 rlbp_macro_307/HI la_data_out[109] sky130_fd_sc_hd__conb_1
Xoutput121 _3487_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[10] sky130_fd_sc_hd__buf_2
X_2627_ _3183_/A vssd1 vssd1 vccd1 vccd1 _2778_/A sky130_fd_sc_hd__buf_2
X_2558_ _2586_/B vssd1 vssd1 vccd1 vccd1 _2568_/B sky130_fd_sc_hd__clkbuf_1
Xrlbp_macro_318 vssd1 vssd1 vccd1 vccd1 rlbp_macro_318/HI la_data_out[120] sky130_fd_sc_hd__conb_1
Xrlbp_macro_329 vssd1 vssd1 vccd1 vccd1 rlbp_macro_329/HI wbs_dat_o[15] sky130_fd_sc_hd__conb_1
XFILLER_99_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2489_ _2565_/A _2491_/B vssd1 vssd1 vccd1 vccd1 _2489_/X sky130_fd_sc_hd__or2_1
XFILLER_83_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_479 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3039__B2 _3491_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2334__A _3457_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3211__A1 _2574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input47_A wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_519 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2509__A _2586_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1860_ _1860_/A _1860_/B vssd1 vssd1 vccd1 vccd1 _1918_/B sky130_fd_sc_hd__nor2_1
Xinput12 la_data_in[16] vssd1 vssd1 vccd1 vccd1 _3802_/A sky130_fd_sc_hd__clkbuf_2
X_1791_ _3443_/Q _2190_/B vssd1 vssd1 vccd1 vccd1 _1791_/X sky130_fd_sc_hd__and2b_1
Xinput45 wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 input45/X sky130_fd_sc_hd__clkbuf_1
Xinput34 la_data_in[6] vssd1 vssd1 vccd1 vccd1 _3792_/A sky130_fd_sc_hd__clkbuf_2
Xinput23 la_data_in[27] vssd1 vssd1 vccd1 vccd1 _3779_/A sky130_fd_sc_hd__buf_2
X_3530_ _3533_/CLK _3530_/D vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__dfxtp_1
XFILLER_10_390 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput56 wbs_dat_i[2] vssd1 vssd1 vccd1 vccd1 _3232_/A sky130_fd_sc_hd__clkbuf_4
X_3461_ _3462_/CLK _3461_/D vssd1 vssd1 vccd1 vccd1 _3461_/Q sky130_fd_sc_hd__dfxtp_1
X_3392_ _3392_/CLK _3392_/D vssd1 vssd1 vccd1 vccd1 _3392_/Q sky130_fd_sc_hd__dfxtp_1
X_2412_ _3307_/Q _2412_/B _2412_/C vssd1 vssd1 vccd1 vccd1 _2412_/X sky130_fd_sc_hd__and3_1
XFILLER_42_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2343_ _2343_/A _2343_/B vssd1 vssd1 vccd1 vccd1 _2345_/B sky130_fd_sc_hd__xor2_1
XANTENNA__3803__A _3803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2274_ _2339_/A _2320_/B vssd1 vssd1 vccd1 vccd1 _2280_/A sky130_fd_sc_hd__and2_1
XFILLER_65_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2244__A2 _1667_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1989_ _3325_/Q _1989_/B vssd1 vssd1 vccd1 vccd1 _2006_/B sky130_fd_sc_hd__xnor2_1
XFILLER_4_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrlbp_macro_148 vssd1 vssd1 vccd1 vccd1 rlbp_macro_148/HI io_oeb[15] sky130_fd_sc_hd__conb_1
XFILLER_0_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrlbp_macro_137 vssd1 vssd1 vccd1 vccd1 rlbp_macro_137/HI io_oeb[4] sky130_fd_sc_hd__conb_1
XANTENNA__1800__B_N _3448_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrlbp_macro_159 vssd1 vssd1 vccd1 vccd1 rlbp_macro_159/HI io_oeb[26] sky130_fd_sc_hd__conb_1
XFILLER_28_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_3_net107_A clkbuf_leaf_9_net107/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2306__B_N _1974_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_375 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2226__A2 _2037_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2961_ _3469_/Q _2948_/X _2960_/X _2958_/X vssd1 vssd1 vccd1 vccd1 _3469_/D sky130_fd_sc_hd__o211a_1
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1912_ _3413_/Q _1912_/B vssd1 vssd1 vccd1 vccd1 _1920_/A sky130_fd_sc_hd__xnor2_1
X_2892_ _2966_/A _2899_/B vssd1 vssd1 vccd1 vccd1 _2892_/X sky130_fd_sc_hd__or2_1
X_1843_ _1786_/A _1842_/X _1786_/B vssd1 vssd1 vccd1 vccd1 _3292_/D sky130_fd_sc_hd__o21ai_1
XFILLER_30_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1774_ _3447_/Q _1774_/B vssd1 vssd1 vccd1 vccd1 _1775_/B sky130_fd_sc_hd__and2b_1
Xclkbuf_leaf_24_net107 _3436_/CLK vssd1 vssd1 vccd1 vccd1 _3462_/CLK sky130_fd_sc_hd__clkbuf_16
X_3513_ _3528_/CLK _3513_/D vssd1 vssd1 vccd1 vccd1 _3521_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_89_419 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3444_ _3445_/CLK _3444_/D vssd1 vssd1 vccd1 vccd1 _3444_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3375_ _3377_/CLK _3375_/D vssd1 vssd1 vccd1 vccd1 _3375_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1973__B_N _2106_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2326_ _3467_/Q _1678_/Y _2325_/Y vssd1 vssd1 vccd1 vccd1 _2328_/A sky130_fd_sc_hd__o21ai_1
X_2257_ _2260_/A _2260_/B vssd1 vssd1 vccd1 vccd1 _2259_/B sky130_fd_sc_hd__xor2_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2188_ _2134_/A _2187_/X _2134_/B vssd1 vssd1 vccd1 vccd1 _3552_/D sky130_fd_sc_hd__o21ai_1
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2059__A _3349_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1898__A _3410_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_500 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_566 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2522__A _2559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3160_ _3160_/A _3160_/B vssd1 vssd1 vccd1 vccd1 _3188_/B sky130_fd_sc_hd__nand2_1
XFILLER_39_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2111_ _1774_/B _3363_/Q vssd1 vssd1 vccd1 vccd1 _2113_/A sky130_fd_sc_hd__and2b_1
XANTENNA__3072__B _3072_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1 hold3/X vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__dlygate4sd3_1
X_3091_ _3447_/Q _2872_/A _3008_/A _3495_/Q vssd1 vssd1 vccd1 vccd1 _3091_/X sky130_fd_sc_hd__a22o_1
XFILLER_94_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2042_ _3356_/Q _2042_/B vssd1 vssd1 vccd1 vccd1 _2100_/B sky130_fd_sc_hd__xnor2_2
XFILLER_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2944_ _2944_/A vssd1 vssd1 vccd1 vccd1 _2945_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2875_ _2875_/A _2875_/B vssd1 vssd1 vccd1 vccd1 _2903_/B sky130_fd_sc_hd__nand2_1
X_1826_ _3435_/Q _1826_/B vssd1 vssd1 vccd1 vccd1 _1832_/B sky130_fd_sc_hd__nand2_1
XANTENNA__2432__A _2561_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1757_ _1757_/A vssd1 vssd1 vccd1 vccd1 _2119_/B sky130_fd_sc_hd__buf_2
X_1688_ _2389_/B vssd1 vssd1 vccd1 vccd1 _2385_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3427_ _3427_/CLK _3427_/D vssd1 vssd1 vccd1 vccd1 _3427_/Q sky130_fd_sc_hd__dfxtp_1
X_3358_ _3377_/CLK _3358_/D vssd1 vssd1 vccd1 vccd1 _3358_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2309_ _2309_/A _3472_/Q vssd1 vssd1 vccd1 vccd1 _2309_/X sky130_fd_sc_hd__or2b_1
XFILLER_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3289_ hold2/X _3281_/A _3282_/A vssd1 vssd1 vccd1 vccd1 _3289_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_57_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2607__A _2762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2061__B _3350_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output116_A _3528_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2517__A _3223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_352 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2660_ _2771_/A _2666_/B vssd1 vssd1 vccd1 vccd1 _2660_/X sky130_fd_sc_hd__or2_1
XFILLER_60_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2591_ _3036_/A vssd1 vssd1 vccd1 vccd1 _2595_/B sky130_fd_sc_hd__clkbuf_2
X_3212_ _3508_/Q _3221_/B vssd1 vssd1 vccd1 vccd1 _3212_/X sky130_fd_sc_hd__or2_1
XFILLER_79_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3143_ _3319_/Q _2988_/X _3012_/A _3142_/X vssd1 vssd1 vccd1 vccd1 _3143_/X sky130_fd_sc_hd__a211o_1
XFILLER_82_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_116 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3074_ _3074_/A vssd1 vssd1 vccd1 vccd1 _3074_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_27_319 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2025_ _3347_/Q _2025_/B vssd1 vssd1 vccd1 vccd1 _2080_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__2427__A _2427_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2927_ _2964_/A _2936_/B vssd1 vssd1 vccd1 vccd1 _2927_/X sky130_fd_sc_hd__or2_1
XANTENNA__2162__A _3371_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3258__A _3525_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2858_ _3435_/Q _2853_/X _2857_/X _2851_/X vssd1 vssd1 vccd1 vccd1 _3435_/D sky130_fd_sc_hd__o211a_1
X_1809_ _1809_/A _1809_/B vssd1 vssd1 vccd1 vccd1 _1822_/B sky130_fd_sc_hd__xnor2_1
X_2789_ _2808_/A vssd1 vssd1 vccd1 vccd1 _2789_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_403 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_36 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3168__A _3234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2800__A _2955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_488 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3075__A2 _3036_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2712_ _2788_/A _2715_/B vssd1 vssd1 vccd1 vccd1 _2728_/A sky130_fd_sc_hd__and2_1
XFILLER_9_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2643_ _2679_/A _2643_/B vssd1 vssd1 vccd1 vccd1 _2672_/B sky130_fd_sc_hd__nand2_1
XANTENNA__3806__A _3806_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2574_ _2574_/A _2582_/B vssd1 vssd1 vccd1 vccd1 _2574_/X sky130_fd_sc_hd__or2_1
XFILLER_87_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2510__A1 _3332_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3126_ _3342_/Q _2996_/X _3037_/A _3462_/Q vssd1 vssd1 vccd1 vccd1 _3126_/X sky130_fd_sc_hd__a22o_1
XFILLER_82_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3260__B _3262_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_436 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3057_ _3348_/Q _2554_/A _2840_/B _3432_/Q vssd1 vssd1 vccd1 vccd1 _3057_/X sky130_fd_sc_hd__a22o_1
XFILLER_23_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2008_ _3329_/Q _2009_/B vssd1 vssd1 vccd1 vccd1 _2008_/Y sky130_fd_sc_hd__nand2_1
XFILLER_35_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2577__A1 _3352_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_403 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2514__B _3006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_82 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2290_ _2290_/A _2347_/B _2343_/A vssd1 vssd1 vccd1 vccd1 _2296_/A sky130_fd_sc_hd__and3_1
XFILLER_77_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_263 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2705__A _2780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1861__A_N _1774_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput100 _3555_/Q vssd1 vssd1 vccd1 vccd1 Sw2 sky130_fd_sc_hd__buf_2
X_2626_ _3365_/Q _2612_/X _2625_/X _2619_/X vssd1 vssd1 vccd1 vccd1 _3365_/D sky130_fd_sc_hd__o211a_1
XANTENNA__2440__A _3236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput111 _3523_/Q vssd1 vssd1 vccd1 vccd1 io_out[25] sky130_fd_sc_hd__buf_2
Xoutput122 _3488_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[11] sky130_fd_sc_hd__buf_2
XANTENNA__2217__A_N _3394_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2557_ _2679_/A _2557_/B vssd1 vssd1 vccd1 vccd1 _2586_/B sky130_fd_sc_hd__nand2_1
Xrlbp_macro_308 vssd1 vssd1 vccd1 vccd1 rlbp_macro_308/HI la_data_out[110] sky130_fd_sc_hd__conb_1
Xrlbp_macro_319 vssd1 vssd1 vccd1 vccd1 rlbp_macro_319/HI la_data_out[121] sky130_fd_sc_hd__conb_1
XFILLER_87_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2488_ _3323_/Q _2479_/X _2486_/X _2487_/X vssd1 vssd1 vccd1 vccd1 _3323_/D sky130_fd_sc_hd__o211a_1
XFILLER_95_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3109_ _3316_/Q _2988_/X _3012_/A _3108_/X vssd1 vssd1 vccd1 vccd1 _3109_/X sky130_fd_sc_hd__a211o_1
XFILLER_15_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2615__A _2769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_483 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_30 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3181__A _3181_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2525__A _2561_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput13 la_data_in[17] vssd1 vssd1 vccd1 vccd1 _3803_/A sky130_fd_sc_hd__clkbuf_2
X_1790_ _1812_/A _1813_/B _1789_/X vssd1 vssd1 vccd1 vccd1 _1816_/B sky130_fd_sc_hd__a21o_1
XANTENNA__3059__C _3059_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput35 la_data_in[7] vssd1 vssd1 vccd1 vccd1 _3793_/A sky130_fd_sc_hd__buf_2
Xinput46 wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 _2511_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput24 la_data_in[28] vssd1 vssd1 vccd1 vccd1 _3805_/A sky130_fd_sc_hd__buf_2
XFILLER_6_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput57 wbs_dat_i[3] vssd1 vssd1 vccd1 vccd1 _3234_/A sky130_fd_sc_hd__clkbuf_4
X_3460_ _3462_/CLK _3460_/D vssd1 vssd1 vccd1 vccd1 _3460_/Q sky130_fd_sc_hd__dfxtp_1
X_3391_ _3392_/CLK _3391_/D vssd1 vssd1 vccd1 vccd1 _3391_/Q sky130_fd_sc_hd__dfxtp_1
X_2411_ _2412_/B _2412_/C _2410_/Y _2397_/X vssd1 vssd1 vccd1 vccd1 _3306_/D sky130_fd_sc_hd__o211a_1
XFILLER_69_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2342_ _2290_/A _2333_/B _2308_/Y vssd1 vssd1 vccd1 vccd1 _2343_/B sky130_fd_sc_hd__a21o_1
XFILLER_96_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2273_ _3474_/Q _3306_/Q vssd1 vssd1 vccd1 vccd1 _2320_/B sky130_fd_sc_hd__xnor2_1
XFILLER_84_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2435__A _2563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_280 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1988_ _1988_/A _1988_/B vssd1 vssd1 vccd1 vccd1 _1989_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__2170__A _3377_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2609_ _3236_/A vssd1 vssd1 vccd1 vccd1 _2765_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrlbp_macro_138 vssd1 vssd1 vccd1 vccd1 rlbp_macro_138/HI io_oeb[5] sky130_fd_sc_hd__conb_1
Xrlbp_macro_149 vssd1 vssd1 vccd1 vccd1 rlbp_macro_149/HI io_oeb[16] sky130_fd_sc_hd__conb_1
XANTENNA__2180__A2 _1922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_59 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2329__B _2330_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_523 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2960_ _2960_/A _2960_/B vssd1 vssd1 vccd1 vccd1 _2960_/X sky130_fd_sc_hd__or2_1
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1911_ _1911_/A _1911_/B vssd1 vssd1 vccd1 vccd1 _1912_/B sky130_fd_sc_hd__xor2_1
X_2891_ _3446_/Q _2888_/X _2890_/X _2882_/X vssd1 vssd1 vccd1 vccd1 _3446_/D sky130_fd_sc_hd__o211a_1
X_1842_ _1822_/X _1842_/B _1842_/C _1842_/D vssd1 vssd1 vccd1 vccd1 _1842_/X sky130_fd_sc_hd__and4b_1
XFILLER_8_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3187__A1 _3499_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1773_ _1774_/B _3447_/Q vssd1 vssd1 vccd1 vccd1 _1775_/A sky130_fd_sc_hd__and2b_1
X_3512_ _3512_/CLK _3512_/D vssd1 vssd1 vccd1 vccd1 _3512_/Q sky130_fd_sc_hd__dfxtp_1
X_3443_ _3445_/CLK _3443_/D vssd1 vssd1 vccd1 vccd1 _3443_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3374_ _3377_/CLK _3374_/D vssd1 vssd1 vccd1 vccd1 _3374_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2325_ _2335_/A _2335_/B vssd1 vssd1 vccd1 vccd1 _2325_/Y sky130_fd_sc_hd__nand2_1
XFILLER_97_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2256_ _2212_/A _2235_/B _2224_/Y vssd1 vssd1 vccd1 vccd1 _2260_/B sky130_fd_sc_hd__a21oi_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3111__A1 _3377_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2187_ _2168_/X _2187_/B _2187_/C _2187_/D vssd1 vssd1 vccd1 vccd1 _2187_/X sky130_fd_sc_hd__and4b_1
XFILLER_65_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_486 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_512 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_30_net107 _3436_/CLK vssd1 vssd1 vccd1 vccd1 _3450_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_44_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_402 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2803__A _2957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3169__A1 _3492_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2916__A1 _3453_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_486 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3090_ _3339_/Q _2996_/X _2997_/X _3375_/Q _3089_/X vssd1 vssd1 vccd1 vccd1 _3095_/A
+ sky130_fd_sc_hd__a221o_1
X_2110_ _2110_/A _2110_/B vssd1 vssd1 vccd1 vccd1 _2173_/B sky130_fd_sc_hd__nor2_1
XFILLER_58_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2041_ _2041_/A _2091_/B _2087_/A vssd1 vssd1 vccd1 vccd1 _2048_/B sky130_fd_sc_hd__and3_1
XFILLER_54_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_331 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_90 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2943_ _2943_/A _3006_/B vssd1 vssd1 vccd1 vccd1 _2944_/A sky130_fd_sc_hd__nor2_1
X_2874_ _2888_/A vssd1 vssd1 vccd1 vccd1 _2874_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1825_ _3435_/Q _1826_/B vssd1 vssd1 vccd1 vccd1 _1832_/A sky130_fd_sc_hd__or2_1
X_1756_ _3449_/Q _2313_/B vssd1 vssd1 vccd1 vccd1 _1759_/A sky130_fd_sc_hd__nor2_1
X_1687_ _3298_/Q vssd1 vssd1 vccd1 vccd1 _2389_/B sky130_fd_sc_hd__clkbuf_4
X_3426_ _3427_/CLK _3426_/D vssd1 vssd1 vccd1 vccd1 _3426_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3357_ _3404_/CLK _3357_/D vssd1 vssd1 vccd1 vccd1 _3357_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_412 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2308_ _2305_/X _2306_/X _2307_/X vssd1 vssd1 vccd1 vccd1 _2308_/Y sky130_fd_sc_hd__a21oi_1
X_3288_ hold2/X _3281_/A _3282_/A vssd1 vssd1 vccd1 vccd1 _3288_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2239_ _2239_/A _2239_/B vssd1 vssd1 vccd1 vccd1 _2255_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__3096__B1 _3088_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_35_net107_A _3494_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_68 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input22_A la_data_in[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output109_A _3521_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2598__C1 _2580_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_272 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2590_ _2979_/B vssd1 vssd1 vccd1 vccd1 _3036_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3211_ _2574_/A _3207_/X _3210_/Y _3200_/X vssd1 vssd1 vccd1 vccd1 _3507_/D sky130_fd_sc_hd__o211a_1
XFILLER_79_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3142_ _3499_/Q _3160_/B _3138_/X _3141_/X vssd1 vssd1 vccd1 vccd1 _3142_/X sky130_fd_sc_hd__a211o_1
XFILLER_82_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3073_ _3481_/Q _2990_/X _3072_/X _3031_/X vssd1 vssd1 vccd1 vccd1 _3481_/D sky130_fd_sc_hd__o211a_1
X_2024_ _1949_/A _3345_/Q vssd1 vssd1 vccd1 vccd1 _2074_/B sky130_fd_sc_hd__nand2b_1
XFILLER_54_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2443__A _3199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2926_ _2941_/B vssd1 vssd1 vccd1 vccd1 _2936_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__3258__B _3262_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2857_ _2966_/A _2863_/B vssd1 vssd1 vccd1 vccd1 _2857_/X sky130_fd_sc_hd__or2_1
X_1808_ _3434_/Q _1808_/B vssd1 vssd1 vccd1 vccd1 _1809_/B sky130_fd_sc_hd__xnor2_1
X_2788_ _2788_/A _2791_/B vssd1 vssd1 vccd1 vccd1 _2808_/A sky130_fd_sc_hd__and2_1
X_1739_ _3548_/Q _3549_/Q vssd1 vssd1 vccd1 vccd1 _2049_/A sky130_fd_sc_hd__or2b_1
XFILLER_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3409_ _3409_/CLK _3409_/D vssd1 vssd1 vccd1 vccd1 _3409_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_242 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_415 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2618__A _2771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_212 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2711_ _2711_/A vssd1 vssd1 vccd1 vccd1 _2715_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__2141__B_N _1794_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2642_ _2656_/A vssd1 vssd1 vccd1 vccd1 _2642_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2573_ _3350_/Q _2570_/X _2572_/X _2566_/X vssd1 vssd1 vccd1 vccd1 _3350_/D sky130_fd_sc_hd__o211a_1
XFILLER_99_378 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2438__A _2565_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3125_ _3426_/Q _2786_/A _3042_/X _3510_/Q vssd1 vssd1 vccd1 vccd1 _3125_/X sky130_fd_sc_hd__a22o_1
XFILLER_82_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3260__C _3262_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3056_ _3056_/A vssd1 vssd1 vccd1 vccd1 _3195_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_70_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2007_ _2007_/A _2007_/B vssd1 vssd1 vccd1 vccd1 _2009_/B sky130_fd_sc_hd__xor2_1
XFILLER_70_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2173__A _3376_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2909_ _3158_/A _2911_/B vssd1 vssd1 vccd1 vccd1 _2925_/A sky130_fd_sc_hd__and2_1
XANTENNA__2901__A _2975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_334 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3179__A _3243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2811__A _2964_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_94 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_540 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2413__D1 _2381_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput101 _3540_/Q vssd1 vssd1 vccd1 vccd1 Vd1 sky130_fd_sc_hd__buf_2
X_2625_ _2775_/A _2628_/B vssd1 vssd1 vccd1 vccd1 _2625_/X sky130_fd_sc_hd__or2_1
Xoutput112 _3524_/Q vssd1 vssd1 vccd1 vccd1 io_out[26] sky130_fd_sc_hd__buf_2
Xoutput123 _3478_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[1] sky130_fd_sc_hd__buf_2
XFILLER_99_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2556_ _2570_/A vssd1 vssd1 vccd1 vccd1 _2556_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xrlbp_macro_309 vssd1 vssd1 vccd1 vccd1 rlbp_macro_309/HI la_data_out[111] sky130_fd_sc_hd__conb_1
XFILLER_99_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2487_ _3264_/A vssd1 vssd1 vccd1 vccd1 _2487_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_101_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3108_ _3108_/A _3108_/B _3108_/C _3108_/D vssd1 vssd1 vccd1 vccd1 _3108_/X sky130_fd_sc_hd__or4_2
XFILLER_55_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1800__A _2145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3039_ _3443_/Q _3017_/X _3008_/A _3491_/Q vssd1 vssd1 vccd1 vccd1 _3039_/X sky130_fd_sc_hd__a22o_1
XFILLER_43_418 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2631__A _2780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_42 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2806__A _2960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1710__A _3496_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput14 la_data_in[18] vssd1 vssd1 vccd1 vccd1 _3780_/A sky130_fd_sc_hd__buf_2
Xinput36 la_data_in[8] vssd1 vssd1 vccd1 vccd1 _3794_/A sky130_fd_sc_hd__clkbuf_2
Xinput25 la_data_in[29] vssd1 vssd1 vccd1 vccd1 _3806_/A sky130_fd_sc_hd__clkbuf_2
Xinput58 wbs_dat_i[4] vssd1 vssd1 vccd1 vccd1 _3236_/A sky130_fd_sc_hd__clkbuf_4
Xinput47 wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 _2982_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_2410_ _2412_/B _2412_/C vssd1 vssd1 vccd1 vccd1 _2410_/Y sky130_fd_sc_hd__nand2_1
X_3390_ _3392_/CLK _3390_/D vssd1 vssd1 vccd1 vccd1 _3390_/Q sky130_fd_sc_hd__dfxtp_1
X_2341_ _3461_/Q _2341_/B vssd1 vssd1 vccd1 vccd1 _2341_/X sky130_fd_sc_hd__or2_1
XFILLER_69_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2272_ _3473_/Q _2407_/A vssd1 vssd1 vccd1 vccd1 _2339_/A sky130_fd_sc_hd__xnor2_2
XFILLER_96_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_292 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1987_ _1987_/A _1987_/B vssd1 vssd1 vccd1 vccd1 _2006_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__2451__A _3241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2608_ _3360_/Q _2593_/X _2607_/X _2601_/X vssd1 vssd1 vccd1 vccd1 _3360_/D sky130_fd_sc_hd__o211a_1
XFILLER_88_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2539_ _3339_/Q _2533_/X _2538_/X _2536_/X vssd1 vssd1 vccd1 vccd1 _3339_/D sky130_fd_sc_hd__o211a_1
Xrlbp_macro_139 vssd1 vssd1 vccd1 vccd1 rlbp_macro_139/HI io_oeb[6] sky130_fd_sc_hd__conb_1
XANTENNA__3282__A _3282_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_59 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2202__B_N _2282_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2361__A _3549_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input52_A wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2536__A _2566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1910_ _1910_/A _1910_/B _1910_/C _1910_/D vssd1 vssd1 vccd1 vccd1 _1910_/X sky130_fd_sc_hd__or4_1
X_2890_ _2964_/A _2899_/B vssd1 vssd1 vccd1 vccd1 _2890_/X sky130_fd_sc_hd__or2_1
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1841_ _1841_/A _1841_/B vssd1 vssd1 vccd1 vccd1 _1842_/D sky130_fd_sc_hd__xnor2_1
XFILLER_8_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1772_ _1772_/A _1772_/B vssd1 vssd1 vccd1 vccd1 _1830_/B sky130_fd_sc_hd__nor2_1
X_3511_ _3511_/CLK _3511_/D vssd1 vssd1 vccd1 vccd1 _3511_/Q sky130_fd_sc_hd__dfxtp_1
X_3442_ _3445_/CLK _3442_/D vssd1 vssd1 vccd1 vccd1 _3442_/Q sky130_fd_sc_hd__dfxtp_1
X_3373_ _3377_/CLK _3373_/D vssd1 vssd1 vccd1 vccd1 _3373_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_134 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2324_ _2324_/A _2324_/B vssd1 vssd1 vccd1 vccd1 _2338_/B sky130_fd_sc_hd__xnor2_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_307 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2255_ _2255_/A _2255_/B _2255_/C _2255_/D vssd1 vssd1 vccd1 vccd1 _2269_/B sky130_fd_sc_hd__or4_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2186_ _3379_/Q _2186_/B vssd1 vssd1 vccd1 vccd1 _2187_/D sky130_fd_sc_hd__xnor2_1
XFILLER_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_94_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2040_ _2040_/A _2040_/B vssd1 vssd1 vccd1 vccd1 _2087_/A sky130_fd_sc_hd__nor2_1
XFILLER_35_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2852__A1 _3433_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_568 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2942_ _3464_/Q _2925_/A _2941_/X _2939_/X vssd1 vssd1 vccd1 vccd1 _3464_/D sky130_fd_sc_hd__o211a_1
X_2873_ _3158_/A _2875_/B vssd1 vssd1 vccd1 vccd1 _2888_/A sky130_fd_sc_hd__and2_1
X_1824_ _1824_/A _1824_/B vssd1 vssd1 vccd1 vccd1 _1826_/B sky130_fd_sc_hd__xnor2_1
X_1755_ _2389_/C _3441_/Q vssd1 vssd1 vccd1 vccd1 _1813_/B sky130_fd_sc_hd__nand2b_1
X_1686_ _1686_/A _1686_/B _1686_/C _1686_/D vssd1 vssd1 vccd1 vccd1 _3262_/B sky130_fd_sc_hd__or4_4
X_3425_ _3427_/CLK _3425_/D vssd1 vssd1 vccd1 vccd1 _3425_/Q sky130_fd_sc_hd__dfxtp_1
X_3356_ _3356_/CLK _3356_/D vssd1 vssd1 vccd1 vccd1 _3356_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_424 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3287_ _3280_/X _3281_/X _3282_/X vssd1 vssd1 vccd1 vccd1 _3287_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_57_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2307_ _1974_/X _3470_/Q vssd1 vssd1 vccd1 vccd1 _2307_/X sky130_fd_sc_hd__and2b_1
X_2238_ _3386_/Q _2238_/B vssd1 vssd1 vccd1 vccd1 _2239_/B sky130_fd_sc_hd__xnor2_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3096__A1 _3315_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2176__A _3375_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2169_ _2169_/A _2169_/B vssd1 vssd1 vccd1 vccd1 _2170_/B sky130_fd_sc_hd__xor2_1
XFILLER_53_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2843__A1 _3429_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3020__B2 _3490_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2052__A_N _3346_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input15_A la_data_in[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3087__A1 _3363_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2814__A _2966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3011__A1 _3309_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3210_ _3210_/A _3219_/B vssd1 vssd1 vccd1 vccd1 _3210_/Y sky130_fd_sc_hd__nand2_1
X_3141_ _3439_/Q _2840_/B _2911_/B _3463_/Q _3140_/X vssd1 vssd1 vccd1 vccd1 _3141_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_94_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3078__B2 _3374_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3072_ _3121_/A _3072_/B vssd1 vssd1 vccd1 vccd1 _3072_/X sky130_fd_sc_hd__or2_1
X_2023_ _3346_/Q _2052_/B vssd1 vssd1 vccd1 vccd1 _2073_/A sky130_fd_sc_hd__xnor2_1
XFILLER_35_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2724__A _2762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3250__A1 _3522_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2925_ _2925_/A vssd1 vssd1 vccd1 vccd1 _2925_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3258__C _3262_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2856_ _3434_/Q _2853_/X _2855_/X _2851_/X vssd1 vssd1 vccd1 vccd1 _3434_/D sky130_fd_sc_hd__o211a_1
X_1807_ _1810_/A _1810_/B _1795_/X vssd1 vssd1 vccd1 vccd1 _1809_/A sky130_fd_sc_hd__a21bo_1
X_2787_ _2787_/A vssd1 vssd1 vccd1 vccd1 _2791_/B sky130_fd_sc_hd__clkbuf_2
X_1738_ _1946_/A _3544_/Q vssd1 vssd1 vccd1 vccd1 _3540_/D sky130_fd_sc_hd__nor2_1
X_1669_ _3509_/Q vssd1 vssd1 vccd1 vccd1 _3215_/A sky130_fd_sc_hd__inv_2
X_3408_ _3409_/CLK _3408_/D vssd1 vssd1 vccd1 vccd1 _3408_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_input7_A la_data_in[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3339_ _3520_/CLK _3339_/D vssd1 vssd1 vccd1 vccd1 _3339_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_427 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3069__B2 _3373_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_376 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2634__A _2782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3293__CLK _3436_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2809__A _3238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2544__A _2582_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_368 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2710_ _3041_/A vssd1 vssd1 vccd1 vccd1 _2711_/A sky130_fd_sc_hd__clkbuf_2
X_2641_ _2788_/A _2643_/B vssd1 vssd1 vccd1 vccd1 _2656_/A sky130_fd_sc_hd__and2_1
XFILLER_9_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2572_ _2572_/A _2582_/B vssd1 vssd1 vccd1 vccd1 _2572_/X sky130_fd_sc_hd__or2_1
XFILLER_99_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_318 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3124_ _3330_/Q _2480_/B _2557_/B _3354_/Q _3123_/X vssd1 vssd1 vccd1 vccd1 _3124_/X
+ sky130_fd_sc_hd__a221o_1
X_3055_ _3336_/Q _2520_/B _2643_/B _3372_/Q _3054_/X vssd1 vssd1 vccd1 vccd1 _3059_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2006_ _2006_/A _2006_/B _2006_/C _2006_/D vssd1 vssd1 vccd1 vccd1 _2021_/B sky130_fd_sc_hd__or4_1
XFILLER_63_482 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2454__A _3243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2908_ _3037_/A vssd1 vssd1 vccd1 vccd1 _2911_/B sky130_fd_sc_hd__clkbuf_2
X_2839_ _2853_/A vssd1 vssd1 vccd1 vccd1 _2839_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_519 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3214__A1 _2576_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_390 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3195__A _3225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2274__A _2339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2413__C1 _3808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2624_ _3181_/A vssd1 vssd1 vccd1 vccd1 _2775_/A sky130_fd_sc_hd__buf_2
Xoutput102 _3545_/Q vssd1 vssd1 vccd1 vccd1 Vd2 sky130_fd_sc_hd__buf_2
Xoutput113 _3525_/Q vssd1 vssd1 vccd1 vccd1 io_out[27] sky130_fd_sc_hd__buf_2
Xoutput124 _3479_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[2] sky130_fd_sc_hd__buf_2
X_2555_ _3223_/A _2557_/B vssd1 vssd1 vccd1 vccd1 _2570_/A sky130_fd_sc_hd__and2_1
XFILLER_99_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2486_ _2563_/A _2491_/B vssd1 vssd1 vccd1 vccd1 _2486_/X sky130_fd_sc_hd__or2_1
XANTENNA__2449__A _2572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_148 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3107_ _3400_/Q _2715_/B _3195_/B _3508_/Q _3106_/X vssd1 vssd1 vccd1 vccd1 _3108_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_70_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3038_ _3359_/Q _3036_/X _3037_/X _3455_/Q vssd1 vssd1 vccd1 vccd1 _3038_/X sky130_fd_sc_hd__a22o_1
XFILLER_70_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_2_2__f_net107 clkbuf_0_net107/X vssd1 vssd1 vccd1 vccd1 _3436_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_87_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_13_net107 clkbuf_2_3__f_net107/X vssd1 vssd1 vccd1 vccd1 _3407_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_61_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2094__A _3354_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1710__B _2037_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput37 la_data_in[9] vssd1 vssd1 vccd1 vccd1 _3795_/A sky130_fd_sc_hd__buf_2
Xinput26 la_data_in[2] vssd1 vssd1 vccd1 vccd1 _3788_/A sky130_fd_sc_hd__clkbuf_2
Xinput15 la_data_in[19] vssd1 vssd1 vccd1 vccd1 _3781_/A sky130_fd_sc_hd__buf_2
Xinput59 wbs_dat_i[5] vssd1 vssd1 vccd1 vccd1 _3238_/A sky130_fd_sc_hd__clkbuf_4
Xinput48 wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 _2982_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2136__A_N _3358_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2340_ _3461_/Q _2341_/B vssd1 vssd1 vccd1 vccd1 _2340_/Y sky130_fd_sc_hd__nand2_1
X_2271_ _3564_/Q _3563_/Q vssd1 vssd1 vccd1 vccd1 _2271_/X sky130_fd_sc_hd__and2b_1
XFILLER_2_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3123__B1 _3041_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1901__A _3405_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1685__B1 _1678_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1986_ _3330_/Q _1986_/B vssd1 vssd1 vccd1 vccd1 _1987_/B sky130_fd_sc_hd__xnor2_1
XFILLER_20_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2607_ _2762_/A _2610_/B vssd1 vssd1 vccd1 vccd1 _2607_/X sky130_fd_sc_hd__or2_1
X_2538_ _2574_/A _2544_/B vssd1 vssd1 vccd1 vccd1 _2538_/X sky130_fd_sc_hd__or2_1
XFILLER_87_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2469_ _3320_/Q _2446_/A _2468_/X _2462_/X vssd1 vssd1 vccd1 vccd1 _3320_/D sky130_fd_sc_hd__o211a_1
XFILLER_68_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1811__A _3433_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_29_net107_A _3436_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2361__B _3548_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2089__A _3339_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1903__A1 _3406_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input45_A wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_0_net107 _3494_/CLK vssd1 vssd1 vccd1 vccd1 _3511_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_78_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3105__B1 _2643_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2817__A _3243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1840_ _3440_/Q _1840_/B vssd1 vssd1 vccd1 vccd1 _1841_/B sky130_fd_sc_hd__xnor2_1
XFILLER_42_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1771_ _3448_/Q _2309_/A vssd1 vssd1 vccd1 vccd1 _1772_/B sky130_fd_sc_hd__and2b_1
X_3510_ _3511_/CLK _3510_/D vssd1 vssd1 vccd1 vccd1 _3510_/Q sky130_fd_sc_hd__dfxtp_1
X_3441_ _3450_/CLK _3441_/D vssd1 vssd1 vccd1 vccd1 _3441_/Q sky130_fd_sc_hd__dfxtp_1
X_3372_ _3377_/CLK _3372_/D vssd1 vssd1 vccd1 vccd1 _3372_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2323_ _3458_/Q _2323_/B vssd1 vssd1 vccd1 vccd1 _2324_/B sky130_fd_sc_hd__xnor2_1
XFILLER_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2254_ _2254_/A _2254_/B _2254_/C _2254_/D vssd1 vssd1 vccd1 vccd1 _2255_/D sky130_fd_sc_hd__or4_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_319 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2185_ _2185_/A _2185_/B vssd1 vssd1 vccd1 vccd1 _2186_/B sky130_fd_sc_hd__xor2_1
XFILLER_80_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2462__A _3264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1969_ _3311_/Q _2025_/B vssd1 vssd1 vccd1 vccd1 _1969_/X sky130_fd_sc_hd__and2b_1
XFILLER_88_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2637__A _3160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_396 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2372__A hold2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_455 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_403 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_94_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2547__A _2566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2941_ _2977_/A _2941_/B vssd1 vssd1 vccd1 vccd1 _2941_/X sky130_fd_sc_hd__or2_1
XANTENNA__3097__B _3097_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2872_ _2872_/A vssd1 vssd1 vccd1 vccd1 _2875_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_1823_ _1776_/A _1810_/B _1799_/Y vssd1 vssd1 vccd1 vccd1 _1824_/B sky130_fd_sc_hd__a21o_1
X_1754_ _3442_/Q _2052_/B vssd1 vssd1 vccd1 vccd1 _1812_/A sky130_fd_sc_hd__xnor2_1
X_3424_ _3474_/CLK _3424_/D vssd1 vssd1 vccd1 vccd1 _3424_/Q sky130_fd_sc_hd__dfxtp_1
X_1685_ _3205_/A _2395_/A _1678_/Y _3503_/Q _1684_/X vssd1 vssd1 vccd1 vccd1 _1686_/D
+ sky130_fd_sc_hd__a221o_1
X_3355_ _3356_/CLK _3355_/D vssd1 vssd1 vccd1 vccd1 _3355_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3286_ _3280_/X _3281_/X _3282_/X vssd1 vssd1 vccd1 vccd1 _3286_/Y sky130_fd_sc_hd__a21oi_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2306_ _3470_/Q _1974_/X vssd1 vssd1 vccd1 vccd1 _2306_/X sky130_fd_sc_hd__or2b_1
XFILLER_85_436 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2237_ _2235_/A _2235_/B _2223_/X vssd1 vssd1 vccd1 vccd1 _2239_/A sky130_fd_sc_hd__a21bo_1
XFILLER_73_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2457__A _3181_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2168_ _2168_/A _2168_/B _2168_/C _2168_/D vssd1 vssd1 vccd1 vccd1 _2168_/X sky130_fd_sc_hd__or4_1
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2099_ _2097_/A _2097_/B _2045_/A vssd1 vssd1 vccd1 vccd1 _2101_/A sky130_fd_sc_hd__a21oi_1
XFILLER_53_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3087__A2 _3036_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2598__A1 _3357_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2830__A _2977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2770__A1 _3410_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output76_A _3785_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3140_ _3343_/Q _2516_/A _2595_/B _3367_/Q _3139_/X vssd1 vssd1 vccd1 vccd1 _3140_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_39_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrlbp_macro_290 vssd1 vssd1 vccd1 vccd1 rlbp_macro_290/HI la_data_out[92] sky130_fd_sc_hd__conb_1
XFILLER_94_255 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3078__A2 _2516_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2277__A _3467_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3071_ _3313_/Q _2993_/X _3063_/X _3070_/X vssd1 vssd1 vccd1 vccd1 _3072_/B sky130_fd_sc_hd__a211o_1
XFILLER_82_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2022_ _1946_/A _3544_/Q _2021_/X _1963_/Y vssd1 vssd1 vccd1 vccd1 _3542_/D sky130_fd_sc_hd__a31o_1
XFILLER_47_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3250__A2 _3253_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2924_ _3457_/Q _2910_/X _2923_/X _2915_/X vssd1 vssd1 vccd1 vccd1 _3457_/D sky130_fd_sc_hd__o211a_1
XFILLER_31_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2855_ _2964_/A _2863_/B vssd1 vssd1 vccd1 vccd1 _2855_/X sky130_fd_sc_hd__or2_1
X_1806_ _1806_/A _1806_/B vssd1 vssd1 vccd1 vccd1 _1822_/A sky130_fd_sc_hd__xnor2_1
X_2786_ _2786_/A vssd1 vssd1 vccd1 vccd1 _2787_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__2761__A1 _3407_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1737_ _3543_/Q vssd1 vssd1 vccd1 vccd1 _1946_/A sky130_fd_sc_hd__inv_2
X_1668_ _3503_/Q vssd1 vssd1 vccd1 vccd1 _3198_/A sky130_fd_sc_hd__inv_2
X_3407_ _3407_/CLK _3407_/D vssd1 vssd1 vccd1 vccd1 _3407_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3338_ _3520_/CLK _3338_/D vssd1 vssd1 vccd1 vccd1 _3338_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3069__A2 _2516_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3269_ _3269_/A vssd1 vssd1 vccd1 vccd1 _3531_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output114_A _3526_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2640_ _2640_/A vssd1 vssd1 vccd1 vccd1 _2643_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__2991__A1 _2427_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2571_ _2586_/B vssd1 vssd1 vccd1 vccd1 _2582_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_4_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3123_ _3378_/Q _2640_/A _3041_/X _3402_/Q vssd1 vssd1 vccd1 vccd1 _3123_/X sky130_fd_sc_hd__a22o_1
XFILLER_95_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3054_ _3384_/Q _3053_/X _3225_/B _3524_/Q vssd1 vssd1 vccd1 vccd1 _3054_/X sky130_fd_sc_hd__a22o_1
XFILLER_27_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2735__A _2773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2005_ _1994_/Y _1995_/X _1998_/Y _2000_/Y _2004_/Y vssd1 vssd1 vccd1 vccd1 _2006_/D
+ sky130_fd_sc_hd__a2111o_1
XFILLER_90_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2907_ _2985_/C vssd1 vssd1 vccd1 vccd1 _3037_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2838_ _3158_/A _2840_/B vssd1 vssd1 vccd1 vccd1 _2853_/A sky130_fd_sc_hd__and2_1
X_2769_ _2769_/A _2778_/B vssd1 vssd1 vccd1 vccd1 _2769_/X sky130_fd_sc_hd__or2_1
XFILLER_86_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2645__A _2756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_6_net107_A clkbuf_leaf_9_net107/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2060__B_N _1974_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3195__B _3195_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2725__A1 _3396_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_36_net107 _3494_/CLK vssd1 vssd1 vccd1 vccd1 _3529_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__1724__A _3498_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2555__A _3223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_70 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2623_ _3364_/Q _2612_/X _2622_/X _2619_/X vssd1 vssd1 vccd1 vccd1 _3364_/D sky130_fd_sc_hd__o211a_1
Xoutput103 _3805_/X vssd1 vssd1 vccd1 vccd1 Vref_cmp_c sky130_fd_sc_hd__buf_2
XFILLER_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput114 _3526_/Q vssd1 vssd1 vccd1 vccd1 io_out[28] sky130_fd_sc_hd__buf_2
Xoutput125 _3480_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[3] sky130_fd_sc_hd__buf_2
X_2554_ _2554_/A vssd1 vssd1 vccd1 vccd1 _2557_/B sky130_fd_sc_hd__clkbuf_2
X_2485_ _3322_/Q _2479_/X _2484_/X _2462_/X vssd1 vssd1 vccd1 vccd1 _3322_/D sky130_fd_sc_hd__o211a_1
XFILLER_68_520 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3141__B2 _3463_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3141__A1 _3439_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3106_ _3352_/Q _2554_/A _2840_/B _3436_/Q vssd1 vssd1 vccd1 vccd1 _3106_/X sky130_fd_sc_hd__a22o_1
XANTENNA__2465__A _2584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3037_ _3037_/A vssd1 vssd1 vccd1 vccd1 _3037_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_43_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput16 la_data_in[1] vssd1 vssd1 vccd1 vccd1 _3787_/A sky130_fd_sc_hd__buf_2
Xinput27 la_data_in[30] vssd1 vssd1 vccd1 vccd1 _1708_/S sky130_fd_sc_hd__clkbuf_1
XFILLER_6_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput38 wb_rst_i vssd1 vssd1 vccd1 vccd1 _2378_/A sky130_fd_sc_hd__clkbuf_2
Xinput49 wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 _2905_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2270_ _2189_/Y _2213_/X _2269_/X _3555_/D vssd1 vssd1 vccd1 vccd1 _3557_/D sky130_fd_sc_hd__a22o_1
XFILLER_69_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3123__A1 _3378_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1985_ _2007_/A _2007_/B _1956_/A vssd1 vssd1 vccd1 vccd1 _1987_/A sky130_fd_sc_hd__a21o_1
XANTENNA__3539__RESET_B _3277_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2937__A1 _3462_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2606_ _3234_/A vssd1 vssd1 vccd1 vccd1 _2762_/A sky130_fd_sc_hd__clkbuf_2
X_2537_ _3338_/Q _2533_/X _2535_/X _2536_/X vssd1 vssd1 vccd1 vccd1 _3338_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2468_ _2586_/A _2468_/B vssd1 vssd1 vccd1 vccd1 _2468_/X sky130_fd_sc_hd__or2_1
XFILLER_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3114__A1 _3365_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3114__B2 _3497_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2399_ _2399_/A _2399_/B vssd1 vssd1 vccd1 vccd1 _2405_/C sky130_fd_sc_hd__and2_1
XFILLER_83_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2923__A _2960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3105__B2 _3376_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input38_A wb_rst_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2552__B _3002_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1770_ _3304_/Q vssd1 vssd1 vccd1 vccd1 _2309_/A sky130_fd_sc_hd__clkbuf_2
X_3440_ _3440_/CLK _3440_/D vssd1 vssd1 vccd1 vccd1 _3440_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3371_ _3377_/CLK _3371_/D vssd1 vssd1 vccd1 vccd1 _3371_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2322_ _2333_/A _2333_/B _2305_/X vssd1 vssd1 vccd1 vccd1 _2324_/A sky130_fd_sc_hd__a21bo_1
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2253_ _2253_/A _2253_/B vssd1 vssd1 vccd1 vccd1 _2254_/D sky130_fd_sc_hd__or2_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1912__A _3413_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2184_ _2184_/A _2184_/B vssd1 vssd1 vccd1 vccd1 _2187_/C sky130_fd_sc_hd__xnor2_1
XFILLER_65_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_38_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1968_ _2001_/A _2001_/B _1967_/X vssd1 vssd1 vccd1 vccd1 _1999_/B sky130_fd_sc_hd__a21o_1
X_1899_ _1899_/A _1899_/B vssd1 vssd1 vccd1 vccd1 _1910_/C sky130_fd_sc_hd__xnor2_1
XFILLER_88_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2653__A _2765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1821__A1 _3430_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2276__A_N _1949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_611 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_467 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_50 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1732__A _2442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_62_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_507 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2563__A _2563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2940_ _3463_/Q _2925_/A _2938_/X _2939_/X vssd1 vssd1 vccd1 vccd1 _3463_/D sky130_fd_sc_hd__o211a_1
X_2871_ _3017_/A vssd1 vssd1 vccd1 vccd1 _2872_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2282__B _2282_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1822_ _1822_/A _1822_/B _1822_/C _1822_/D vssd1 vssd1 vccd1 vccd1 _1822_/X sky130_fd_sc_hd__or4_1
XFILLER_30_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3494__CLK _3494_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1753_ _3298_/Q vssd1 vssd1 vccd1 vccd1 _2052_/B sky130_fd_sc_hd__clkbuf_4
X_1684_ _3208_/A _2399_/A _2046_/B _3501_/Q vssd1 vssd1 vccd1 vccd1 _1684_/X sky130_fd_sc_hd__a22o_1
X_3423_ _3474_/CLK _3423_/D vssd1 vssd1 vccd1 vccd1 _3423_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3354_ _3512_/CLK _3354_/D vssd1 vssd1 vccd1 vccd1 _3354_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3285_ _3280_/X _3281_/X _3282_/X vssd1 vssd1 vccd1 vccd1 _3285_/Y sky130_fd_sc_hd__a21oi_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2305_ _3469_/Q _1794_/X vssd1 vssd1 vccd1 vccd1 _2305_/X sky130_fd_sc_hd__or2b_1
X_2236_ _3385_/Q _2236_/B vssd1 vssd1 vccd1 vccd1 _2255_/A sky130_fd_sc_hd__xnor2_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2167_ _2167_/A _2167_/B _2167_/C _2167_/D vssd1 vssd1 vccd1 vccd1 _2168_/D sky130_fd_sc_hd__or4_1
XFILLER_53_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2098_ _3343_/Q _2098_/B vssd1 vssd1 vccd1 vccd1 _2102_/C sky130_fd_sc_hd__xnor2_1
XFILLER_80_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1817__A _3431_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_172 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_13_net107_A clkbuf_2_3__f_net107/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output69_A _3778_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrlbp_macro_291 vssd1 vssd1 vccd1 vccd1 rlbp_macro_291/HI la_data_out[93] sky130_fd_sc_hd__conb_1
Xrlbp_macro_280 vssd1 vssd1 vccd1 vccd1 rlbp_macro_280/HI la_data_out[82] sky130_fd_sc_hd__conb_1
XFILLER_39_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3070_ _3070_/A _3070_/B _3070_/C vssd1 vssd1 vccd1 vccd1 _3070_/X sky130_fd_sc_hd__or3_1
XFILLER_94_267 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2021_ _2021_/A _2021_/B _2021_/C _2021_/D vssd1 vssd1 vccd1 vccd1 _2021_/X sky130_fd_sc_hd__or4_1
XANTENNA__2277__B _3299_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_175 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2923_ _2960_/A _2923_/B vssd1 vssd1 vccd1 vccd1 _2923_/X sky130_fd_sc_hd__or2_1
X_2854_ _2868_/B vssd1 vssd1 vccd1 vccd1 _2863_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_31_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1805_ _3438_/Q _1805_/B vssd1 vssd1 vccd1 vccd1 _1806_/B sky130_fd_sc_hd__xnor2_1
X_2785_ _2985_/B vssd1 vssd1 vccd1 vccd1 _2786_/A sky130_fd_sc_hd__clkbuf_2
X_1736_ _1874_/A vssd1 vssd1 vccd1 vccd1 _3535_/D sky130_fd_sc_hd__clkinv_2
X_1667_ _2389_/A vssd1 vssd1 vccd1 vccd1 _1667_/X sky130_fd_sc_hd__clkbuf_2
X_3406_ _3407_/CLK _3406_/D vssd1 vssd1 vccd1 vccd1 _3406_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3337_ _3520_/CLK _3337_/D vssd1 vssd1 vccd1 vccd1 _3337_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2468__A _2586_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3268_ _2378_/X input3/X vssd1 vssd1 vccd1 vccd1 _3269_/A sky130_fd_sc_hd__and2b_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2219_ _3395_/Q vssd1 vssd1 vccd1 vccd1 _2219_/Y sky130_fd_sc_hd__inv_2
X_3199_ _3199_/A vssd1 vssd1 vccd1 vccd1 _3251_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_26_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2378__A _2378_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input20_A la_data_in[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3002__A _3002_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2976__C1 _2971_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2570_ _2570_/A vssd1 vssd1 vccd1 vccd1 _2570_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_99_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3122_ _3485_/Q _3074_/X _3121_/X _3098_/X vssd1 vssd1 vccd1 vccd1 _3485_/D sky130_fd_sc_hd__o211a_1
XFILLER_55_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3053_ _3053_/A vssd1 vssd1 vccd1 vccd1 _3053_/X sky130_fd_sc_hd__buf_2
XFILLER_67_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2004_ _2004_/A _2004_/B vssd1 vssd1 vccd1 vccd1 _2004_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2906_ _2983_/A _3006_/B vssd1 vssd1 vccd1 vccd1 _2985_/C sky130_fd_sc_hd__nor2_1
XFILLER_31_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2837_ _2837_/A vssd1 vssd1 vccd1 vccd1 _2840_/B sky130_fd_sc_hd__clkbuf_2
X_2768_ _2782_/B vssd1 vssd1 vccd1 vccd1 _2778_/B sky130_fd_sc_hd__clkbuf_1
X_2699_ _2731_/A vssd1 vssd1 vccd1 vccd1 _2699_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1719_ _1719_/A _1719_/B _1719_/C _1718_/Y vssd1 vssd1 vccd1 vccd1 _1719_/X sky130_fd_sc_hd__or4b_1
XFILLER_58_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2498__A1 _3327_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1830__A _3436_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_42 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1724__B _2121_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3150__A2 _3160_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2555__B _2557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2661__A1 _3375_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2413__A1 _2291_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2622_ _2773_/A _2628_/B vssd1 vssd1 vccd1 vccd1 _2622_/X sky130_fd_sc_hd__or2_1
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput104 _3806_/X vssd1 vssd1 vccd1 vccd1 Vref_sel_c sky130_fd_sc_hd__buf_2
Xoutput115 _3527_/Q vssd1 vssd1 vccd1 vccd1 io_out[29] sky130_fd_sc_hd__buf_2
X_2553_ _3000_/A vssd1 vssd1 vccd1 vccd1 _2554_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__1915__A _3411_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput126 _3481_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[4] sky130_fd_sc_hd__buf_2
X_2484_ _2561_/A _2491_/B vssd1 vssd1 vccd1 vccd1 _2484_/X sky130_fd_sc_hd__or2_1
XFILLER_101_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3105_ _3340_/Q _2520_/B _2643_/B _3376_/Q _3104_/X vssd1 vssd1 vccd1 vccd1 _3108_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_68_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3036_ _3036_/A vssd1 vssd1 vccd1 vccd1 _3036_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__2652__A1 _3372_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1825__A _3435_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2891__A1 _3446_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput17 la_data_in[20] vssd1 vssd1 vccd1 vccd1 _3782_/A sky130_fd_sc_hd__buf_2
Xinput28 la_data_in[31] vssd1 vssd1 vccd1 vccd1 _2373_/A sky130_fd_sc_hd__clkbuf_2
Xinput39 wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 _2512_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_6_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2566__A _2566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2331__B1 _3453_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1685__A2 _2395_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2285__B _2285_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1984_ _3331_/Q _1984_/B vssd1 vssd1 vccd1 vccd1 _2021_/A sky130_fd_sc_hd__xnor2_1
XFILLER_20_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2605_ _3359_/Q _2593_/X _2604_/X _2601_/X vssd1 vssd1 vccd1 vccd1 _3359_/D sky130_fd_sc_hd__o211a_1
X_2536_ _2566_/A vssd1 vssd1 vccd1 vccd1 _2536_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2467_ _3188_/A vssd1 vssd1 vccd1 vccd1 _2586_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_87_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2398_ _2395_/A _2394_/A _2396_/Y _2397_/X vssd1 vssd1 vccd1 vccd1 _3301_/D sky130_fd_sc_hd__o211a_1
XFILLER_95_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2195__B _2407_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3019_ _3322_/Q _2981_/A _2985_/A _3406_/Q vssd1 vssd1 vccd1 vccd1 _3019_/X sky130_fd_sc_hd__a22o_1
XFILLER_43_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3050__A1 _3324_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_38_net107_A _3494_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_104 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2616__A1 _3362_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_476 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3370_ _3377_/CLK _3370_/D vssd1 vssd1 vccd1 vccd1 _3370_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2321_ _2321_/A _2321_/B vssd1 vssd1 vccd1 vccd1 _2338_/A sky130_fd_sc_hd__xnor2_1
X_2252_ _2251_/B _2251_/C _3381_/Q vssd1 vssd1 vccd1 vccd1 _2253_/B sky130_fd_sc_hd__a21oi_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2183_ _3380_/Q _2183_/B vssd1 vssd1 vccd1 vccd1 _2184_/B sky130_fd_sc_hd__xor2_1
XFILLER_38_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_535 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1967_ _3310_/Q _2301_/B vssd1 vssd1 vccd1 vccd1 _1967_/X sky130_fd_sc_hd__and2b_1
X_1898_ _3410_/Q _1898_/B vssd1 vssd1 vccd1 vccd1 _1899_/B sky130_fd_sc_hd__xnor2_1
XFILLER_88_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2519_ _2834_/A vssd1 vssd1 vccd1 vccd1 _2679_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_88_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3499_ _3507_/CLK _3499_/D vssd1 vssd1 vccd1 vccd1 _3499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2934__A _2970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3023__A1 _3394_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input50_A wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2844__A _2953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_519 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2870_ _3002_/A _2870_/B vssd1 vssd1 vccd1 vccd1 _3017_/A sky130_fd_sc_hd__nor2_1
X_1821_ _3430_/Q _1812_/Y _1815_/Y _1817_/Y _1820_/Y vssd1 vssd1 vccd1 vccd1 _1822_/D
+ sky130_fd_sc_hd__o2111ai_1
X_1752_ _1816_/A _1819_/B vssd1 vssd1 vccd1 vccd1 _1762_/A sky130_fd_sc_hd__and2_1
X_1683_ _2295_/B vssd1 vssd1 vccd1 vccd1 _2046_/B sky130_fd_sc_hd__buf_2
XFILLER_7_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3422_ _3427_/CLK _3422_/D vssd1 vssd1 vccd1 vccd1 _3422_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3353_ _3512_/CLK _3353_/D vssd1 vssd1 vccd1 vccd1 _3353_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3284_ _3280_/X _3281_/X _3282_/X vssd1 vssd1 vccd1 vccd1 _3284_/Y sky130_fd_sc_hd__a21oi_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2304_ _2300_/Y _1878_/X _2280_/D _2335_/B _2303_/Y vssd1 vssd1 vccd1 vccd1 _2333_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_85_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2235_ _2235_/A _2235_/B vssd1 vssd1 vccd1 vccd1 _2236_/B sky130_fd_sc_hd__xnor2_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2828__A1 _3427_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2166_ _3369_/Q _2166_/B vssd1 vssd1 vccd1 vccd1 _2167_/D sky130_fd_sc_hd__xnor2_1
XFILLER_26_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2097_ _2097_/A _2097_/B vssd1 vssd1 vccd1 vccd1 _2098_/B sky130_fd_sc_hd__xor2_1
XANTENNA__2754__A _2875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3253__A1 _3523_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2056__A2 _1878_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2999_ _3333_/Q _2996_/X _2997_/X _3369_/Q _2998_/X vssd1 vssd1 vccd1 vccd1 _3005_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2664__A _2775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3244__A1 _3528_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_19_net107 clkbuf_2_3__f_net107/X vssd1 vssd1 vccd1 vccd1 _3539_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_67_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrlbp_macro_270 vssd1 vssd1 vccd1 vccd1 rlbp_macro_270/HI la_data_out[72] sky130_fd_sc_hd__conb_1
Xrlbp_macro_281 vssd1 vssd1 vccd1 vccd1 rlbp_macro_281/HI la_data_out[83] sky130_fd_sc_hd__conb_1
Xrlbp_macro_292 vssd1 vssd1 vccd1 vccd1 rlbp_macro_292/HI la_data_out[94] sky130_fd_sc_hd__conb_1
X_2020_ _2020_/A _2020_/B vssd1 vssd1 vccd1 vccd1 _2021_/D sky130_fd_sc_hd__xnor2_1
XFILLER_47_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_279 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2574__A _2574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3235__A1 _3524_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2922_ _3456_/Q _2910_/X _2921_/X _2915_/X vssd1 vssd1 vccd1 vccd1 _3456_/D sky130_fd_sc_hd__o211a_1
XFILLER_93_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1918__A _3412_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2853_ _2853_/A vssd1 vssd1 vccd1 vccd1 _2853_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1804_ _1827_/A _1827_/B _1759_/A vssd1 vssd1 vccd1 vccd1 _1806_/A sky130_fd_sc_hd__a21o_1
X_2784_ _2943_/A _2870_/B vssd1 vssd1 vccd1 vccd1 _2985_/B sky130_fd_sc_hd__nor2_1
X_1735_ _3538_/Q _3539_/Q vssd1 vssd1 vccd1 vccd1 _1874_/A sky130_fd_sc_hd__or2b_1
X_1666_ _2025_/B vssd1 vssd1 vccd1 vccd1 _2389_/A sky130_fd_sc_hd__clkbuf_4
X_3405_ _3407_/CLK _3405_/D vssd1 vssd1 vccd1 vccd1 _3405_/Q sky130_fd_sc_hd__dfxtp_1
X_3336_ _3520_/CLK _3336_/D vssd1 vssd1 vccd1 vccd1 _3336_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1721__A1 _3499_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3267_ _3267_/A vssd1 vssd1 vccd1 vccd1 _3530_/D sky130_fd_sc_hd__clkbuf_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2218_ _2249_/A _2251_/B _2217_/X vssd1 vssd1 vccd1 vccd1 _2247_/B sky130_fd_sc_hd__a21o_1
XFILLER_38_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3198_ _3198_/A _3202_/B vssd1 vssd1 vccd1 vccd1 _3198_/Y sky130_fd_sc_hd__nand2_1
XFILLER_81_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2149_ _2169_/A _2169_/B _2120_/A vssd1 vssd1 vccd1 vccd1 _2151_/A sky130_fd_sc_hd__a21o_1
XANTENNA__2484__A _2561_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_335 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input13_A la_data_in[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3002__B _3006_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_530 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_6_net107 clkbuf_leaf_9_net107/A vssd1 vssd1 vccd1 vccd1 _3516_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_13_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3121_ _3121_/A _3121_/B vssd1 vssd1 vccd1 vccd1 _3121_/X sky130_fd_sc_hd__or2_1
XANTENNA__2288__B _2288_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3052_ _3420_/Q _2787_/A _2946_/A _3468_/Q _3051_/X vssd1 vssd1 vccd1 vccd1 _3059_/B
+ sky130_fd_sc_hd__a221o_1
X_2003_ _3322_/Q _2003_/B _2003_/C vssd1 vssd1 vccd1 vccd1 _2004_/B sky130_fd_sc_hd__and3_1
XFILLER_63_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2905_ _2982_/C _2905_/B _2982_/A _2982_/B vssd1 vssd1 vccd1 vccd1 _3006_/B sky130_fd_sc_hd__or4bb_4
X_2836_ _3021_/A vssd1 vssd1 vccd1 vccd1 _2837_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__1648__A _2395_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2767_ _2767_/A vssd1 vssd1 vccd1 vccd1 _2767_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2698_ _2773_/A _2703_/B vssd1 vssd1 vccd1 vccd1 _2698_/X sky130_fd_sc_hd__or2_1
X_1718_ _3489_/Q _2295_/B _1717_/X vssd1 vssd1 vccd1 vccd1 _1718_/Y sky130_fd_sc_hd__a21boi_1
X_1649_ _3511_/Q vssd1 vssd1 vccd1 vccd1 _3219_/A sky130_fd_sc_hd__inv_2
XFILLER_86_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input5_A la_data_in[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3319_ _3322_/CLK _3319_/D vssd1 vssd1 vccd1 vccd1 _3319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2389__A _2389_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3135__B1 _2711_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2621_ _3243_/A vssd1 vssd1 vccd1 vccd1 _2773_/A sky130_fd_sc_hd__clkbuf_2
Xoutput116 _3528_/Q vssd1 vssd1 vccd1 vccd1 io_out[30] sky130_fd_sc_hd__buf_2
XFILLER_56_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput105 _2385_/C vssd1 vssd1 vccd1 vccd1 io_out[19] sky130_fd_sc_hd__buf_2
X_2552_ _2552_/A _3002_/A vssd1 vssd1 vccd1 vccd1 _3000_/A sky130_fd_sc_hd__nor2_1
XFILLER_99_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput127 _3482_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[5] sky130_fd_sc_hd__buf_2
XANTENNA__2299__A _3474_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2483_ _3321_/Q _2479_/X _2482_/X _2462_/X vssd1 vssd1 vccd1 vccd1 _3321_/D sky130_fd_sc_hd__o211a_1
XFILLER_68_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3104_ _3388_/Q _3053_/X _3225_/B _3528_/Q vssd1 vssd1 vccd1 vccd1 _3104_/X sky130_fd_sc_hd__a22o_1
X_3035_ _3335_/Q _2520_/B _2643_/B _3371_/Q _3034_/X vssd1 vssd1 vccd1 vccd1 _3035_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_55_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2762__A _2762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_308 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3799_ input9/X vssd1 vssd1 vccd1 vccd1 _3799_/X sky130_fd_sc_hd__clkbuf_1
X_2819_ _3424_/Q _2808_/X _2818_/X _2815_/X vssd1 vssd1 vccd1 vccd1 _3424_/D sky130_fd_sc_hd__o211a_1
XFILLER_3_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_102 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2672__A _2782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput18 la_data_in[21] vssd1 vssd1 vccd1 vccd1 _3783_/A sky130_fd_sc_hd__buf_2
Xinput29 la_data_in[32] vssd1 vssd1 vccd1 vccd1 _1748_/S sky130_fd_sc_hd__clkbuf_1
XFILLER_6_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2331__A1 _2330_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2582__A _2582_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2398__A1 _2395_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1983_ _1983_/A _1983_/B vssd1 vssd1 vccd1 vccd1 _1984_/B sky130_fd_sc_hd__xnor2_1
X_2604_ _2760_/A _2610_/B vssd1 vssd1 vccd1 vccd1 _2604_/X sky130_fd_sc_hd__or2_1
X_2535_ _2572_/A _2544_/B vssd1 vssd1 vccd1 vccd1 _2535_/X sky130_fd_sc_hd__or2_1
XFILLER_87_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2466_ _3319_/Q _2446_/A _2465_/X _2462_/X vssd1 vssd1 vccd1 vccd1 _3319_/D sky130_fd_sc_hd__o211a_1
XFILLER_87_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2397_ _2397_/A vssd1 vssd1 vccd1 vccd1 _2397_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_3_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1661__A _3508_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3018_ _3018_/A vssd1 vssd1 vccd1 vccd1 _3018_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2667__A _2742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_547 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_411 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_488 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2320_ _3462_/Q _2320_/B vssd1 vssd1 vccd1 vccd1 _2321_/B sky130_fd_sc_hd__xnor2_1
XFILLER_97_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2251_ _3381_/Q _2251_/B _2251_/C vssd1 vssd1 vccd1 vccd1 _2253_/A sky130_fd_sc_hd__and3_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2182_ _2185_/A _2185_/B _2117_/A vssd1 vssd1 vccd1 vccd1 _2184_/A sky130_fd_sc_hd__a21oi_1
XFILLER_38_547 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1966_ _3312_/Q vssd1 vssd1 vccd1 vccd1 _1966_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1897_ _1895_/A _1895_/B _1884_/X vssd1 vssd1 vccd1 vccd1 _1899_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__1656__A _3300_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2518_ _2533_/A vssd1 vssd1 vccd1 vccd1 _2518_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2543__A1 _3341_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2487__A _3264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3498_ _3507_/CLK _3498_/D vssd1 vssd1 vccd1 vccd1 _3498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2449_ _2572_/A _2461_/B vssd1 vssd1 vccd1 vccd1 _2449_/X sky130_fd_sc_hd__or2_1
XFILLER_84_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1885__B_N _1796_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3023__A2 _2711_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3781__A _3781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input43_A wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_6 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1820_ _1820_/A _1820_/B vssd1 vssd1 vccd1 vccd1 _1820_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1751_ _3444_/Q _2026_/B vssd1 vssd1 vccd1 vccd1 _1819_/B sky130_fd_sc_hd__xnor2_1
XFILLER_30_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1682_ _1682_/A vssd1 vssd1 vccd1 vccd1 _2295_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_99_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3421_ _3476_/CLK _3421_/D vssd1 vssd1 vccd1 vccd1 _3421_/Q sky130_fd_sc_hd__dfxtp_1
X_3352_ _3512_/CLK _3352_/D vssd1 vssd1 vccd1 vccd1 _3352_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_211 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2303_ _3468_/Q _1657_/Y _1678_/Y _3467_/Q vssd1 vssd1 vccd1 vccd1 _2303_/Y sky130_fd_sc_hd__a211oi_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3283_ _3280_/X _3281_/X _3282_/X vssd1 vssd1 vccd1 vccd1 _3283_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_57_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2234_ _2234_/A _2234_/B vssd1 vssd1 vccd1 vccd1 _2269_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__2100__A _3344_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2165_ _2125_/Y _2165_/B vssd1 vssd1 vccd1 vccd1 _2166_/B sky130_fd_sc_hd__and2b_1
XFILLER_38_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2096_ _2094_/Y _1834_/X _2033_/D _2084_/B _2095_/X vssd1 vssd1 vccd1 vccd1 _2097_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_26_539 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3253__A2 _3253_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2998_ _3381_/Q _2676_/A _3024_/A _3521_/Q vssd1 vssd1 vccd1 vccd1 _2998_/X sky130_fd_sc_hd__a22o_1
X_1949_ _1949_/A _3309_/Q vssd1 vssd1 vccd1 vccd1 _2001_/B sky130_fd_sc_hd__or2b_1
XFILLER_95_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_300 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_491 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_71 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_22_net107_A _3436_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3180__A1 _3496_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrlbp_macro_260 vssd1 vssd1 vccd1 vccd1 rlbp_macro_260/HI la_data_out[62] sky130_fd_sc_hd__conb_1
XFILLER_67_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrlbp_macro_282 vssd1 vssd1 vccd1 vccd1 rlbp_macro_282/HI la_data_out[84] sky130_fd_sc_hd__conb_1
Xrlbp_macro_271 vssd1 vssd1 vccd1 vccd1 rlbp_macro_271/HI la_data_out[73] sky130_fd_sc_hd__conb_1
Xrlbp_macro_293 vssd1 vssd1 vccd1 vccd1 rlbp_macro_293/HI la_data_out[95] sky130_fd_sc_hd__conb_1
XFILLER_82_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2855__A _2964_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2921_ _2957_/A _2923_/B vssd1 vssd1 vccd1 vccd1 _2921_/X sky130_fd_sc_hd__or2_1
XFILLER_31_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2994__A1 _3357_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2852_ _3433_/Q _2839_/X _2850_/X _2851_/X vssd1 vssd1 vccd1 vccd1 _3433_/D sky130_fd_sc_hd__o211a_1
XANTENNA__2994__B2 _3453_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2783_ _3416_/Q _2767_/A _2782_/X _2776_/X vssd1 vssd1 vccd1 vccd1 _3416_/D sky130_fd_sc_hd__o211a_1
X_1803_ _1785_/B _1810_/B _1802_/X vssd1 vssd1 vccd1 vccd1 _1827_/B sky130_fd_sc_hd__a21o_1
XFILLER_31_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1734_ _1786_/A vssd1 vssd1 vccd1 vccd1 _3295_/D sky130_fd_sc_hd__clkinv_2
XFILLER_7_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3404_ _3404_/CLK _3404_/D vssd1 vssd1 vccd1 vccd1 _3404_/Q sky130_fd_sc_hd__dfxtp_1
X_1665_ _3299_/Q vssd1 vssd1 vccd1 vccd1 _2025_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_98_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3335_ _3520_/CLK _3335_/D vssd1 vssd1 vccd1 vccd1 _3335_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3266_ _2378_/X _3531_/Q vssd1 vssd1 vccd1 vccd1 _3267_/A sky130_fd_sc_hd__and2b_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1721__A2 _1932_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2217_ _3394_/Q _2301_/B vssd1 vssd1 vccd1 vccd1 _2217_/X sky130_fd_sc_hd__and2b_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2765__A _2765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3197_ _2561_/A _3191_/X _3196_/X _3184_/X vssd1 vssd1 vccd1 vccd1 _3502_/D sky130_fd_sc_hd__o211a_1
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2148_ _2133_/B _2155_/B _2147_/X vssd1 vssd1 vccd1 vccd1 _2169_/B sky130_fd_sc_hd__a21o_1
XFILLER_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2079_ _2079_/A _2079_/B vssd1 vssd1 vccd1 vccd1 _2079_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_81_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_25_net107 _3436_/CLK vssd1 vssd1 vccd1 vccd1 _3469_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_30_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2675__A _3053_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_542 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2976__A1 _3475_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3120_ _3317_/Q _2988_/A _3112_/X _3119_/X vssd1 vssd1 vccd1 vccd1 _3121_/B sky130_fd_sc_hd__a211o_1
XFILLER_67_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3051_ _3360_/Q _3036_/A _3037_/X _3456_/Q vssd1 vssd1 vccd1 vccd1 _3051_/X sky130_fd_sc_hd__a22o_1
X_2002_ _2003_/B _2003_/C _3322_/Q vssd1 vssd1 vccd1 vccd1 _2004_/A sky130_fd_sc_hd__a21oi_1
XFILLER_35_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1929__A _3415_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2904_ _3452_/Q _2888_/A _2903_/X _2895_/X vssd1 vssd1 vccd1 vccd1 _3452_/D sky130_fd_sc_hd__o211a_1
X_2835_ _3006_/A _2870_/B vssd1 vssd1 vccd1 vccd1 _3021_/A sky130_fd_sc_hd__nor2_1
XANTENNA__2719__A1 _3393_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2766_ _3409_/Q _2753_/X _2765_/X _2763_/X vssd1 vssd1 vccd1 vccd1 _3409_/D sky130_fd_sc_hd__o211a_1
X_2697_ _3387_/Q _2692_/X _2696_/X _2686_/X vssd1 vssd1 vccd1 vccd1 _3387_/D sky130_fd_sc_hd__o211a_1
X_1717_ _3492_/Q _1657_/Y _1682_/A _3489_/Q _1716_/Y vssd1 vssd1 vccd1 vccd1 _1717_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_6_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1648_ _2395_/A vssd1 vssd1 vccd1 vccd1 _1648_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3318_ _3491_/CLK _3318_/D vssd1 vssd1 vccd1 vccd1 _3318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3249_ _3521_/Q _3256_/B _3256_/C vssd1 vssd1 vccd1 vccd1 _3249_/X sky130_fd_sc_hd__or3_1
XFILLER_58_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2495__A _2572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2389__B _2389_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3135__A1 _3379_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_420 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output112_A _3524_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_423 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2620_ _3363_/Q _2612_/X _2618_/X _2619_/X vssd1 vssd1 vccd1 vccd1 _3363_/D sky130_fd_sc_hd__o211a_1
Xoutput106 _2381_/B vssd1 vssd1 vccd1 vccd1 io_out[20] sky130_fd_sc_hd__buf_2
X_2551_ _2551_/A _2551_/B vssd1 vssd1 vccd1 vccd1 _3002_/A sky130_fd_sc_hd__or2_2
XFILLER_99_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput117 _3808_/X vssd1 vssd1 vccd1 vccd1 io_out[31] sky130_fd_sc_hd__buf_2
XANTENNA__1924__A2 _1834_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput128 _3483_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[6] sky130_fd_sc_hd__buf_2
XFILLER_5_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2482_ _2559_/A _2491_/B vssd1 vssd1 vccd1 vccd1 _2482_/X sky130_fd_sc_hd__or2_1
XFILLER_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_opt_1_0_net107_A clkbuf_leaf_9_net107/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3126__A1 _3342_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3126__B2 _3462_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3103_ _3364_/Q _2595_/B _2911_/B _3460_/Q _3102_/X vssd1 vssd1 vccd1 vccd1 _3108_/B
+ sky130_fd_sc_hd__a221o_1
X_3034_ _3383_/Q _2679_/B _3225_/B _3523_/Q vssd1 vssd1 vccd1 vccd1 _3034_/X sky130_fd_sc_hd__a22o_1
XFILLER_83_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1659__A _2285_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2124__B_N _3357_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3798_ input8/X vssd1 vssd1 vccd1 vccd1 _3798_/X sky130_fd_sc_hd__clkbuf_1
X_2818_ _2968_/A _2824_/B vssd1 vssd1 vccd1 vccd1 _2818_/X sky130_fd_sc_hd__or2_1
X_2749_ _2985_/A vssd1 vssd1 vccd1 vccd1 _2750_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3117__A1 _3341_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3117__B2 _3461_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_567 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1773__A_N _1774_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2953__A _2953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3784__A _3784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput19 la_data_in[22] vssd1 vssd1 vccd1 vccd1 _3784_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_96_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1751__B _2026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2331__A2 _2330_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3024__A _3024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_518 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2863__A _2973_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1982_ _1965_/Y _1834_/X _1959_/B _2007_/B _1981_/X vssd1 vssd1 vccd1 vccd1 _1983_/B
+ sky130_fd_sc_hd__a221oi_4
XFILLER_9_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2603_ _3232_/A vssd1 vssd1 vccd1 vccd1 _2760_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_9_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2534_ _2549_/B vssd1 vssd1 vccd1 vccd1 _2544_/B sky130_fd_sc_hd__clkbuf_1
X_2465_ _2584_/A _2468_/B vssd1 vssd1 vccd1 vccd1 _2465_/X sky130_fd_sc_hd__or2_1
XANTENNA__1942__A _3313_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2396_ _2399_/B vssd1 vssd1 vccd1 vccd1 _2396_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2773__A _2773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3017_ _3017_/A vssd1 vssd1 vccd1 vccd1 _3017_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_434 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3035__B1 _2643_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2013__A _3327_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3779__A _3779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2683__A _2758_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_423 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2250_ _3382_/Q _2250_/B vssd1 vssd1 vccd1 vccd1 _2254_/C sky130_fd_sc_hd__xnor2_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_6 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2304__A2 _1878_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2181_ _2179_/Y _1834_/X _2132_/A _2169_/B _2180_/X vssd1 vssd1 vccd1 vccd1 _2185_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_65_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_559 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_378 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_326 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1815__A1 _3430_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_426 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1965_ _3318_/Q vssd1 vssd1 vccd1 vccd1 _1965_/Y sky130_fd_sc_hd__inv_2
X_1896_ _3409_/Q _1896_/B vssd1 vssd1 vccd1 vccd1 _1910_/B sky130_fd_sc_hd__xnor2_1
X_2517_ _3223_/A _2520_/B vssd1 vssd1 vccd1 vccd1 _2533_/A sky130_fd_sc_hd__and2_1
X_3497_ _3507_/CLK _3497_/D vssd1 vssd1 vccd1 vccd1 _3497_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1672__A _2282_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2448_ _2468_/B vssd1 vssd1 vccd1 vccd1 _2461_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_56_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2379_ _2378_/X input2/X vssd1 vssd1 vccd1 vccd1 _2380_/A sky130_fd_sc_hd__and2b_1
XFILLER_83_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input36_A la_data_in[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1750_ _3443_/Q _2025_/B vssd1 vssd1 vccd1 vccd1 _1816_/A sky130_fd_sc_hd__xnor2_1
XFILLER_11_481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1681_ _1949_/A vssd1 vssd1 vccd1 vccd1 _1682_/A sky130_fd_sc_hd__inv_2
XFILLER_99_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3420_ _3427_/CLK _3420_/D vssd1 vssd1 vccd1 vccd1 _3420_/Q sky130_fd_sc_hd__dfxtp_1
X_3351_ _3512_/CLK _3351_/D vssd1 vssd1 vccd1 vccd1 _3351_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2302_ _2329_/A _2330_/B _2301_/X vssd1 vssd1 vccd1 vccd1 _2335_/B sky130_fd_sc_hd__a21o_1
XFILLER_31_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3282_ _3282_/A vssd1 vssd1 vccd1 vccd1 _3282_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2233_ _3392_/Q _2233_/B vssd1 vssd1 vccd1 vccd1 _2234_/B sky130_fd_sc_hd__xnor2_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2164_ _3370_/Q _2164_/B vssd1 vssd1 vccd1 vccd1 _2167_/C sky130_fd_sc_hd__xnor2_1
XFILLER_93_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2095_ _2094_/Y _1693_/A _2030_/A vssd1 vssd1 vccd1 vccd1 _2095_/X sky130_fd_sc_hd__o21a_1
XANTENNA__3212__A _3508_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1667__A _2389_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2997_ _2997_/A vssd1 vssd1 vccd1 vccd1 _2997_/X sky130_fd_sc_hd__clkbuf_2
X_1948_ _3310_/Q _2301_/B vssd1 vssd1 vccd1 vccd1 _2001_/A sky130_fd_sc_hd__xnor2_1
XFILLER_21_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1879_ _3418_/Q _2052_/B vssd1 vssd1 vccd1 vccd1 _1879_/X sky130_fd_sc_hd__and2b_1
XFILLER_1_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3549_ _3559_/CLK _3549_/D _3284_/Y vssd1 vssd1 vccd1 vccd1 _3549_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_507 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_9_net107_A clkbuf_leaf_9_net107/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3792__A _3792_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3165__C1 _3156_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1715__B1 _1667_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrlbp_macro_250 vssd1 vssd1 vccd1 vccd1 rlbp_macro_250/HI la_data_out[52] sky130_fd_sc_hd__conb_1
XFILLER_67_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrlbp_macro_272 vssd1 vssd1 vccd1 vccd1 rlbp_macro_272/HI la_data_out[74] sky130_fd_sc_hd__conb_1
Xrlbp_macro_261 vssd1 vssd1 vccd1 vccd1 rlbp_macro_261/HI la_data_out[63] sky130_fd_sc_hd__conb_1
Xrlbp_macro_283 vssd1 vssd1 vccd1 vccd1 rlbp_macro_283/HI la_data_out[85] sky130_fd_sc_hd__conb_1
Xrlbp_macro_294 vssd1 vssd1 vccd1 vccd1 rlbp_macro_294/HI la_data_out[96] sky130_fd_sc_hd__conb_1
XFILLER_85_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2920_ _3455_/Q _2910_/X _2919_/X _2915_/X vssd1 vssd1 vccd1 vccd1 _3455_/D sky130_fd_sc_hd__o211a_1
XFILLER_43_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2851_ _2895_/A vssd1 vssd1 vccd1 vccd1 _2851_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2782_ _2782_/A _2782_/B vssd1 vssd1 vccd1 vccd1 _2782_/X sky130_fd_sc_hd__or2_1
X_1802_ _1830_/B _1824_/A _1799_/Y _1801_/X vssd1 vssd1 vccd1 vccd1 _1802_/X sky130_fd_sc_hd__a31o_1
X_1733_ _3293_/Q _3294_/Q vssd1 vssd1 vccd1 vccd1 _1786_/A sky130_fd_sc_hd__or2b_1
XFILLER_7_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3403_ _3404_/CLK _3403_/D vssd1 vssd1 vccd1 vccd1 _3403_/Q sky130_fd_sc_hd__dfxtp_1
X_1664_ _1757_/A vssd1 vssd1 vccd1 vccd1 _2313_/B sky130_fd_sc_hd__clkbuf_4
X_3334_ _3520_/CLK _3334_/D vssd1 vssd1 vccd1 vccd1 _3334_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3265_ _3265_/A vssd1 vssd1 vccd1 vccd1 _3529_/D sky130_fd_sc_hd__clkbuf_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2216_ _3396_/Q vssd1 vssd1 vccd1 vccd1 _2216_/Y sky130_fd_sc_hd__inv_2
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3196_ _3502_/Q _3221_/B vssd1 vssd1 vccd1 vccd1 _3196_/X sky130_fd_sc_hd__or2_1
XFILLER_26_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_495 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2147_ _2173_/B _2175_/A _2144_/Y _2146_/X vssd1 vssd1 vccd1 vccd1 _2147_/X sky130_fd_sc_hd__a31o_1
XFILLER_53_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2078_ _3336_/Q _2078_/B vssd1 vssd1 vccd1 vccd1 _2079_/B sky130_fd_sc_hd__xnor2_1
XFILLER_26_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1844__B _2025_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2673__A1 _3380_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3787__A _3787_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1754__B _2052_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output67_A _3808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2866__A _2975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1770__A _3304_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3050_ _3324_/Q _2477_/A _2751_/A _3408_/Q _3049_/X vssd1 vssd1 vccd1 vccd1 _3059_/A
+ sky130_fd_sc_hd__a221o_1
X_2001_ _2001_/A _2001_/B vssd1 vssd1 vccd1 vccd1 _2003_/C sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_31_net107 _3436_/CLK vssd1 vssd1 vccd1 vccd1 _3435_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_36_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2903_ _2977_/A _2903_/B vssd1 vssd1 vccd1 vccd1 _2903_/X sky130_fd_sc_hd__or2_1
XFILLER_31_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2106__A _3362_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2834_ _2834_/A vssd1 vssd1 vccd1 vccd1 _3158_/A sky130_fd_sc_hd__clkbuf_2
X_2765_ _2765_/A _2765_/B vssd1 vssd1 vccd1 vccd1 _2765_/X sky130_fd_sc_hd__or2_1
X_2696_ _2771_/A _2703_/B vssd1 vssd1 vccd1 vccd1 _2696_/X sky130_fd_sc_hd__or2_1
X_1716_ _3500_/Q _3308_/Q vssd1 vssd1 vccd1 vccd1 _1716_/Y sky130_fd_sc_hd__xnor2_1
X_1647_ _2281_/B vssd1 vssd1 vccd1 vccd1 _2395_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_100_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3317_ _3491_/CLK _3317_/D vssd1 vssd1 vccd1 vccd1 _3317_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3248_ _3521_/Q _3253_/A2 _3239_/X _3247_/X vssd1 vssd1 vccd1 vccd1 _3521_/D sky130_fd_sc_hd__o211a_1
XFILLER_73_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2655__A1 _3373_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3179_ _3243_/A _3183_/B vssd1 vssd1 vccd1 vccd1 _3179_/X sky130_fd_sc_hd__or2_1
XFILLER_39_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3080__A1 _3326_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3080__B2 _3410_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2389__C _2389_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_395 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2646__A1 _3369_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_479 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3071__A1 _3313_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2550_ _3344_/Q _2533_/A _2549_/X _2547_/X vssd1 vssd1 vccd1 vccd1 _3344_/D sky130_fd_sc_hd__o211a_1
Xoutput107 _3516_/CLK vssd1 vssd1 vccd1 vccd1 io_out[21] sky130_fd_sc_hd__clkbuf_1
Xoutput118 _3809_/X vssd1 vssd1 vccd1 vccd1 io_out[32] sky130_fd_sc_hd__buf_2
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput129 _3484_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[7] sky130_fd_sc_hd__buf_2
X_2481_ _2509_/B vssd1 vssd1 vccd1 vccd1 _2491_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_99_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3126__A2 _2996_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3102_ _3424_/Q _2786_/A _2945_/A _3472_/Q vssd1 vssd1 vccd1 vccd1 _3102_/X sky130_fd_sc_hd__a22o_1
X_3033_ _3033_/A vssd1 vssd1 vccd1 vccd1 _3225_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_36_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_126 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3062__B2 _3457_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3062__A1 _3361_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3797_ input7/X vssd1 vssd1 vccd1 vccd1 _3797_/X sky130_fd_sc_hd__clkbuf_1
X_2817_ _3243_/A vssd1 vssd1 vccd1 vccd1 _2968_/A sky130_fd_sc_hd__clkbuf_2
X_2748_ _2983_/A _2870_/B vssd1 vssd1 vccd1 vccd1 _2985_/A sky130_fd_sc_hd__nor2_1
X_2679_ _2679_/A _2679_/B vssd1 vssd1 vccd1 vccd1 _2707_/B sky130_fd_sc_hd__nand2_1
XANTENNA__3117__A2 _2996_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_579 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input66_A wbs_we_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2867__A1 _3439_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2095__A2 _1693_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3044__A1 _3395_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1981_ _1965_/Y _1922_/X _1956_/A vssd1 vssd1 vccd1 vccd1 _1981_/X sky130_fd_sc_hd__o21a_1
XFILLER_9_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2602_ _3358_/Q _2593_/X _2600_/X _2601_/X vssd1 vssd1 vccd1 vccd1 _3358_/D sky130_fd_sc_hd__o211a_1
X_2533_ _2533_/A vssd1 vssd1 vccd1 vccd1 _2533_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2464_ _3186_/A vssd1 vssd1 vccd1 vccd1 _2584_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_68_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2395_ _2395_/A _2395_/B _2395_/C vssd1 vssd1 vccd1 vccd1 _2399_/B sky130_fd_sc_hd__and3_1
XANTENNA__2858__A1 _3435_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1942__B _2281_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3016_ _3418_/Q _2791_/B _2949_/B _3466_/Q _3015_/X vssd1 vssd1 vccd1 vccd1 _3016_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_36_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3035__B2 _3371_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1852__B _2121_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2849__A1 _3432_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2964__A _2964_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_435 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3795__A _3795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3026__B2 _3370_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_16_net107_A clkbuf_2_3__f_net107/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2180_ _2179_/Y _1922_/X _2120_/A vssd1 vssd1 vccd1 vccd1 _2180_/X sky130_fd_sc_hd__o21a_1
XFILLER_65_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2296__D _2330_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1964_ _1946_/A _3544_/Q _1963_/Y vssd1 vssd1 vccd1 vccd1 _3541_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__1937__B _3315_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1895_ _1895_/A _1895_/B vssd1 vssd1 vccd1 vccd1 _1896_/B sky130_fd_sc_hd__xnor2_1
X_2516_ _2516_/A vssd1 vssd1 vccd1 vccd1 _2520_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3496_ _3511_/CLK _3496_/D vssd1 vssd1 vccd1 vccd1 _3496_/Q sky130_fd_sc_hd__dfxtp_1
X_2447_ _3238_/A vssd1 vssd1 vccd1 vccd1 _2572_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_68_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2378_ _2378_/A vssd1 vssd1 vccd1 vccd1 _2378_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_56_335 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2784__A _2943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2231__A2 _1693_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1847__B _2052_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2694__A _2769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input29_A la_data_in[32] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1680_ _3297_/Q vssd1 vssd1 vccd1 vccd1 _1949_/A sky130_fd_sc_hd__buf_2
XANTENNA_output97_A _3295_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3350_ _3512_/CLK _3350_/D vssd1 vssd1 vccd1 vccd1 _3350_/Q sky130_fd_sc_hd__dfxtp_2
X_2301_ _3466_/Q _2301_/B vssd1 vssd1 vccd1 vccd1 _2301_/X sky130_fd_sc_hd__and2b_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3281_ _3281_/A vssd1 vssd1 vccd1 vccd1 _3281_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2232_ _2267_/A _2267_/B _2210_/A vssd1 vssd1 vccd1 vccd1 _2234_/A sky130_fd_sc_hd__a21o_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2163_ _2163_/A _2165_/B vssd1 vssd1 vccd1 vccd1 _2164_/B sky130_fd_sc_hd__xnor2_1
XFILLER_38_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_176 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2094_ _3354_/Q vssd1 vssd1 vccd1 vccd1 _2094_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1948__A _3310_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2996_ _2996_/A vssd1 vssd1 vccd1 vccd1 _2996_/X sky130_fd_sc_hd__buf_2
XFILLER_21_268 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1947_ _3298_/Q vssd1 vssd1 vccd1 vccd1 _2301_/B sky130_fd_sc_hd__clkbuf_4
X_1878_ _2191_/B vssd1 vssd1 vccd1 vccd1 _1878_/X sky130_fd_sc_hd__buf_4
X_3548_ _3559_/CLK _3548_/D _3283_/Y vssd1 vssd1 vccd1 vccd1 _3548_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__1683__A _2295_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3479_ _3529_/CLK _3479_/D vssd1 vssd1 vccd1 vccd1 _3479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3229__A1 _3521_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_519 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2019__A _3332_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_382 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1715__A1 _3497_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2201__B _3398_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrlbp_macro_251 vssd1 vssd1 vccd1 vccd1 rlbp_macro_251/HI la_data_out[53] sky130_fd_sc_hd__conb_1
Xrlbp_macro_240 vssd1 vssd1 vccd1 vccd1 rlbp_macro_240/HI la_data_out[42] sky130_fd_sc_hd__conb_1
Xrlbp_macro_262 vssd1 vssd1 vccd1 vccd1 rlbp_macro_262/HI la_data_out[64] sky130_fd_sc_hd__conb_1
Xrlbp_macro_273 vssd1 vssd1 vccd1 vccd1 rlbp_macro_273/HI la_data_out[75] sky130_fd_sc_hd__conb_1
Xrlbp_macro_284 vssd1 vssd1 vccd1 vccd1 rlbp_macro_284/HI la_data_out[86] sky130_fd_sc_hd__conb_1
Xrlbp_macro_295 vssd1 vssd1 vccd1 vccd1 rlbp_macro_295/HI la_data_out[97] sky130_fd_sc_hd__conb_1
XFILLER_47_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_198 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_31_net107_A _3436_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2850_ _2960_/A _2850_/B vssd1 vssd1 vccd1 vccd1 _2850_/X sky130_fd_sc_hd__or2_1
XANTENNA__1768__A _3304_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1801_ _1800_/X _1775_/B _1772_/B vssd1 vssd1 vccd1 vccd1 _1801_/X sky130_fd_sc_hd__a21o_1
X_2781_ _3415_/Q _2767_/A _2780_/X _2776_/X vssd1 vssd1 vccd1 vccd1 _3415_/D sky130_fd_sc_hd__o211a_1
X_1732_ _2442_/A vssd1 vssd1 vccd1 vccd1 _2381_/B sky130_fd_sc_hd__clkinv_2
XANTENNA__2599__A _3230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1663_ _3305_/Q vssd1 vssd1 vccd1 vccd1 _1757_/A sky130_fd_sc_hd__inv_2
X_3402_ _3404_/CLK _3402_/D vssd1 vssd1 vccd1 vccd1 _3402_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3333_ _3520_/CLK _3333_/D vssd1 vssd1 vccd1 vccd1 _3333_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2111__B _3363_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3264_ _3264_/A _3264_/B vssd1 vssd1 vccd1 vccd1 _3265_/A sky130_fd_sc_hd__and2_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2215_ _3402_/Q vssd1 vssd1 vccd1 vccd1 _2215_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3223__A _3223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3195_ _3225_/A _3195_/B vssd1 vssd1 vccd1 vccd1 _3221_/B sky130_fd_sc_hd__and2_1
X_2146_ _2145_/X _2113_/B _2110_/B vssd1 vssd1 vccd1 vccd1 _2146_/X sky130_fd_sc_hd__a21o_1
XFILLER_81_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2077_ _2080_/A _2080_/B _2054_/X vssd1 vssd1 vccd1 vccd1 _2079_/A sky130_fd_sc_hd__a21oi_1
XFILLER_81_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2307__A_N _1974_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1678__A _2190_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2979_ _3000_/A _2979_/B _2997_/A _3053_/A vssd1 vssd1 vccd1 vccd1 _2981_/C sky130_fd_sc_hd__or4_1
XFILLER_100_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3147__B1 _2679_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2000_ _3323_/Q _2000_/B vssd1 vssd1 vccd1 vccd1 _2000_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_35_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2902_ _3451_/Q _2888_/A _2901_/X _2895_/X vssd1 vssd1 vccd1 vccd1 _3451_/D sky130_fd_sc_hd__o211a_1
XANTENNA__2106__B _2106_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2833_ _3428_/Q _2808_/A _2830_/X _2832_/X vssd1 vssd1 vccd1 vccd1 _3428_/D sky130_fd_sc_hd__o211a_1
X_2764_ _3408_/Q _2753_/X _2762_/X _2763_/X vssd1 vssd1 vccd1 vccd1 _3408_/D sky130_fd_sc_hd__o211a_1
XFILLER_8_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1715_ _3497_/Q _2118_/B _1667_/X _1714_/Y vssd1 vssd1 vccd1 vccd1 _1719_/C sky130_fd_sc_hd__a22o_1
X_2695_ _3386_/Q _2692_/X _2694_/X _2686_/X vssd1 vssd1 vccd1 vccd1 _3386_/D sky130_fd_sc_hd__o211a_1
XANTENNA__3129__B1 _2679_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1646_ _3301_/Q vssd1 vssd1 vccd1 vccd1 _2281_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_6_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1961__A _3309_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3316_ _3491_/CLK _3316_/D vssd1 vssd1 vccd1 vccd1 _3316_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_86_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3247_ input1/X _3256_/B _3256_/C vssd1 vssd1 vccd1 vccd1 _3247_/X sky130_fd_sc_hd__or3_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3178_ _3495_/Q _3173_/X _3177_/X _3171_/X vssd1 vssd1 vccd1 vccd1 _3495_/D sky130_fd_sc_hd__o211a_1
X_2129_ _2129_/A _2129_/B vssd1 vssd1 vccd1 vccd1 _2159_/B sky130_fd_sc_hd__nor2_1
XFILLER_81_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1855__B _2105_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2389__D hold5/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3798__A input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input11_A la_data_in[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1909__A1 _3406_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput108 _3807_/X vssd1 vssd1 vccd1 vccd1 io_out[22] sky130_fd_sc_hd__buf_2
Xoutput119 _3529_/Q vssd1 vssd1 vccd1 vccd1 wbs_ack_o sky130_fd_sc_hd__buf_2
X_2480_ _3225_/A _2480_/B vssd1 vssd1 vccd1 vccd1 _2509_/B sky130_fd_sc_hd__nand2_1
XFILLER_99_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2877__A _2951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput90 _3799_/X vssd1 vssd1 vccd1 vccd1 Pd7_b sky130_fd_sc_hd__buf_2
X_3101_ _3328_/Q _2477_/A _2751_/A _3412_/Q _3100_/X vssd1 vssd1 vccd1 vccd1 _3108_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_68_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3032_ _3478_/Q _2990_/X _3029_/X _3031_/X vssd1 vssd1 vccd1 vccd1 _3478_/D sky130_fd_sc_hd__o211a_1
XFILLER_91_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3047__C1 _3046_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_138 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3062__A2 _3036_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2816_ _3423_/Q _2808_/X _2814_/X _2815_/X vssd1 vssd1 vccd1 vccd1 _3423_/D sky130_fd_sc_hd__o211a_1
X_3796_ input6/X vssd1 vssd1 vccd1 vccd1 _3796_/X sky130_fd_sc_hd__clkbuf_1
X_2747_ _2982_/B _2982_/C _2905_/B _2982_/A vssd1 vssd1 vccd1 vccd1 _2870_/B sky130_fd_sc_hd__or4b_2
X_2678_ _2692_/A vssd1 vssd1 vccd1 vccd1 _2678_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2573__A1 _3350_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1691__A _3306_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input3_A io_in[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_160 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2564__A1 _3347_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input59_A wbs_dat_i[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_255 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1980_ _1945_/X _1988_/B _1979_/X vssd1 vssd1 vccd1 vccd1 _2007_/B sky130_fd_sc_hd__a21o_1
XFILLER_33_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3044__A2 _3041_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2601_ _2654_/A vssd1 vssd1 vccd1 vccd1 _2601_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2532_ _3337_/Q _2518_/X _2531_/X _2523_/X vssd1 vssd1 vccd1 vccd1 _3337_/D sky130_fd_sc_hd__o211a_1
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2463_ _3318_/Q _2446_/X _2461_/X _2462_/X vssd1 vssd1 vccd1 vccd1 _3318_/D sky130_fd_sc_hd__o211a_1
X_2394_ _2394_/A _2394_/B vssd1 vssd1 vccd1 vccd1 _3300_/D sky130_fd_sc_hd__nor2_1
X_3015_ _3358_/Q _2595_/B _2911_/B _3454_/Q vssd1 vssd1 vccd1 vccd1 _3015_/X sky130_fd_sc_hd__a22o_1
XFILLER_71_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3779_ _3779_/A vssd1 vssd1 vccd1 vccd1 _3779_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_79_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_491 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_458 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3026__A2 _2516_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2890__A _2964_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1963_ _1963_/A _1963_/B vssd1 vssd1 vccd1 vccd1 _1963_/Y sky130_fd_sc_hd__nor2_1
X_1894_ _1894_/A _1894_/B vssd1 vssd1 vccd1 vccd1 _1910_/A sky130_fd_sc_hd__xnor2_1
X_3564_ _3564_/CLK _3564_/D _3290_/Y vssd1 vssd1 vccd1 vccd1 _3564_/Q sky130_fd_sc_hd__dfrtp_1
X_2515_ _2996_/A vssd1 vssd1 vccd1 vccd1 _2516_/A sky130_fd_sc_hd__clkbuf_2
X_3495_ _3507_/CLK _3495_/D vssd1 vssd1 vccd1 vccd1 _3495_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2130__A _3359_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2446_ _2446_/A vssd1 vssd1 vccd1 vccd1 _2446_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2377_ _2372_/X _2374_/X _2376_/X vssd1 vssd1 vccd1 vccd1 _2377_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_83_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2024__B _3345_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1863__B _2206_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2975__A _2975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_122 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_196 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_564 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_288 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1981__A2 _1922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1773__B _3447_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3280_ hold2/X vssd1 vssd1 vccd1 vccd1 _3280_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2300_ _3468_/Q vssd1 vssd1 vccd1 vccd1 _2300_/Y sky130_fd_sc_hd__inv_2
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2231_ _2215_/Y _1693_/A _2198_/C _2264_/B _2230_/X vssd1 vssd1 vccd1 vccd1 _2267_/B
+ sky130_fd_sc_hd__a221o_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2162_ _3371_/Q _2162_/B vssd1 vssd1 vccd1 vccd1 _2167_/B sky130_fd_sc_hd__xnor2_1
XFILLER_81_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2093_ _2093_/A _2093_/B _2093_/C _2093_/D vssd1 vssd1 vccd1 vccd1 _2102_/B sky130_fd_sc_hd__and4_1
XFILLER_93_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_14_net107 clkbuf_2_3__f_net107/X vssd1 vssd1 vccd1 vccd1 _3404_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_65_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2109__B _2309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_391 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_372 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1730__A_N _2373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1949__B_N _3309_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_564 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1948__B _2301_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2125__A _3357_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2995_ _3417_/Q _2786_/A _2945_/A _3465_/Q _2994_/X vssd1 vssd1 vccd1 vccd1 _3005_/A
+ sky130_fd_sc_hd__a221o_1
X_1946_ _1946_/A _1983_/A _3544_/Q _1945_/X vssd1 vssd1 vccd1 vccd1 _1963_/A sky130_fd_sc_hd__or4b_1
XFILLER_9_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1877_ _3300_/Q vssd1 vssd1 vccd1 vccd1 _2191_/B sky130_fd_sc_hd__clkbuf_2
X_3547_ _3547_/D _2362_/X vssd1 vssd1 vccd1 vccd1 _3549_/D sky130_fd_sc_hd__dlxtn_1
XFILLER_88_236 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3478_ _3529_/CLK _3478_/D vssd1 vssd1 vccd1 vccd1 _3478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2795__A _3230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2429_ _2559_/A _2441_/B vssd1 vssd1 vccd1 vccd1 _2429_/X sky130_fd_sc_hd__or2_1
XFILLER_44_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2035__A _3350_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3165__A1 _3490_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1715__A2 _2118_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input41_A wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrlbp_macro_241 vssd1 vssd1 vccd1 vccd1 rlbp_macro_241/HI la_data_out[43] sky130_fd_sc_hd__conb_1
Xrlbp_macro_230 vssd1 vssd1 vccd1 vccd1 rlbp_macro_230/HI la_data_out[32] sky130_fd_sc_hd__conb_1
XFILLER_79_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrlbp_macro_252 vssd1 vssd1 vccd1 vccd1 rlbp_macro_252/HI la_data_out[54] sky130_fd_sc_hd__conb_1
Xrlbp_macro_263 vssd1 vssd1 vccd1 vccd1 rlbp_macro_263/HI la_data_out[65] sky130_fd_sc_hd__conb_1
Xrlbp_macro_274 vssd1 vssd1 vccd1 vccd1 rlbp_macro_274/HI la_data_out[76] sky130_fd_sc_hd__conb_1
Xrlbp_macro_285 vssd1 vssd1 vccd1 vccd1 rlbp_macro_285/HI la_data_out[87] sky130_fd_sc_hd__conb_1
Xrlbp_macro_296 vssd1 vssd1 vccd1 vccd1 rlbp_macro_296/HI la_data_out[98] sky130_fd_sc_hd__conb_1
XFILLER_47_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2109__A_N _3364_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1800_ _2145_/A _3448_/Q vssd1 vssd1 vccd1 vccd1 _1800_/X sky130_fd_sc_hd__or2b_1
X_2780_ _2780_/A _2782_/B vssd1 vssd1 vccd1 vccd1 _2780_/X sky130_fd_sc_hd__or2_1
X_1731_ hold1/X _2373_/A _2375_/A vssd1 vssd1 vccd1 vccd1 _2442_/A sky130_fd_sc_hd__a21oi_4
X_1662_ _3511_/Q _2115_/B _1657_/Y _3504_/Q _1661_/X vssd1 vssd1 vccd1 vccd1 _1686_/B
+ sky130_fd_sc_hd__a221o_1
X_3401_ _3404_/CLK _3401_/D vssd1 vssd1 vccd1 vccd1 _3401_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3332_ _3332_/CLK _3332_/D vssd1 vssd1 vccd1 vccd1 _3332_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_1_net107 _3494_/CLK vssd1 vssd1 vccd1 vccd1 _3507_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_98_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3263_ _3528_/Q _1707_/A _3264_/A _3262_/X vssd1 vssd1 vccd1 vccd1 _3528_/D sky130_fd_sc_hd__o211a_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2214_ _3555_/D _2189_/Y _2213_/X _2189_/B vssd1 vssd1 vccd1 vccd1 _3556_/D sky130_fd_sc_hd__o22ai_1
X_3194_ _2559_/A _3191_/X _3193_/Y _3184_/X vssd1 vssd1 vccd1 vccd1 _3501_/D sky130_fd_sc_hd__o211a_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2145_ _2145_/A _3364_/Q vssd1 vssd1 vccd1 vccd1 _2145_/X sky130_fd_sc_hd__or2b_1
XFILLER_93_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_456 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2076_ _3334_/Q _2073_/Y _2074_/X _2075_/Y vssd1 vssd1 vccd1 vccd1 _2076_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2978_ _3476_/Q _2962_/A _2977_/X _2971_/X vssd1 vssd1 vccd1 vccd1 _3476_/D sky130_fd_sc_hd__o211a_1
X_1929_ _3415_/Q _1929_/B vssd1 vssd1 vccd1 vccd1 _1930_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__1694__A _3510_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3147__A1 _3380_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1869__A _3427_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3138__A1 _3415_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1779__A _3451_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2901_ _2975_/A _2903_/B vssd1 vssd1 vccd1 vccd1 _2901_/X sky130_fd_sc_hd__or2_1
XFILLER_31_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2832_ _2895_/A vssd1 vssd1 vccd1 vccd1 _2832_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2763_ _2815_/A vssd1 vssd1 vccd1 vccd1 _2763_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2585__C1 _2580_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1714_ _3491_/Q vssd1 vssd1 vccd1 vccd1 _1714_/Y sky130_fd_sc_hd__inv_2
X_2694_ _2769_/A _2703_/B vssd1 vssd1 vccd1 vccd1 _2694_/X sky130_fd_sc_hd__or2_1
X_1645_ _2405_/B vssd1 vssd1 vccd1 vccd1 _1645_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1961__B _2046_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3315_ _3491_/CLK _3315_/D vssd1 vssd1 vccd1 vccd1 _3315_/Q sky130_fd_sc_hd__dfxtp_1
X_3246_ _3262_/C vssd1 vssd1 vccd1 vccd1 _3256_/C sky130_fd_sc_hd__clkbuf_1
XANTENNA__3234__A _3234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3177_ _3241_/A _3183_/B vssd1 vssd1 vccd1 vccd1 _3177_/X sky130_fd_sc_hd__or2_1
XFILLER_39_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2128_ _3360_/Q _2191_/B vssd1 vssd1 vccd1 vccd1 _2129_/B sky130_fd_sc_hd__and2b_1
X_2059_ _3349_/Q _1794_/X vssd1 vssd1 vccd1 vccd1 _2059_/X sky130_fd_sc_hd__or2b_1
XFILLER_54_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1871__B _2046_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2983__A _2983_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_283 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2223__A _3397_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput109 _3521_/Q vssd1 vssd1 vccd1 vccd1 io_out[23] sky130_fd_sc_hd__buf_2
Xoutput80 _3789_/X vssd1 vssd1 vccd1 vccd1 Pd2_b sky130_fd_sc_hd__buf_2
Xoutput91 _3800_/X vssd1 vssd1 vccd1 vccd1 Pd8_a sky130_fd_sc_hd__buf_2
X_3100_ _3448_/Q _3017_/X _3018_/X _3496_/Q vssd1 vssd1 vccd1 vccd1 _3100_/X sky130_fd_sc_hd__a22o_1
XFILLER_83_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3031_ _3184_/A vssd1 vssd1 vccd1 vccd1 _3031_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2815_ _2815_/A vssd1 vssd1 vccd1 vccd1 _2815_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3795_ _3795_/A vssd1 vssd1 vccd1 vccd1 _3795_/X sky130_fd_sc_hd__clkbuf_1
X_2746_ _3404_/Q _2728_/A _2745_/X _2743_/X vssd1 vssd1 vccd1 vccd1 _3404_/D sky130_fd_sc_hd__o211a_1
XFILLER_8_390 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2677_ _2788_/A _2679_/B vssd1 vssd1 vccd1 vccd1 _2692_/A sky130_fd_sc_hd__and2_1
XANTENNA__1972__A _3313_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3229_ _3521_/Q _3224_/X _3227_/X _3228_/X vssd1 vssd1 vccd1 vccd1 _3513_/D sky130_fd_sc_hd__o211a_1
XFILLER_46_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_172 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1866__B _2042_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2043__A _3355_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_312 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output110_A _3522_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2600_ _2758_/A _2610_/B vssd1 vssd1 vccd1 vccd1 _2600_/X sky130_fd_sc_hd__or2_1
X_2531_ _2568_/A _2531_/B vssd1 vssd1 vccd1 vccd1 _2531_/X sky130_fd_sc_hd__or2_1
XFILLER_5_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2462_ _3264_/A vssd1 vssd1 vccd1 vccd1 _2462_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2393_ _2395_/B _2395_/C _2397_/A vssd1 vssd1 vccd1 vccd1 _2394_/B sky130_fd_sc_hd__o21ai_1
XFILLER_56_507 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3014_ _3155_/A vssd1 vssd1 vccd1 vccd1 _3121_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_83_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3778_ _3778_/A vssd1 vssd1 vccd1 vccd1 _3778_/X sky130_fd_sc_hd__clkbuf_1
X_2729_ _2745_/B vssd1 vssd1 vccd1 vccd1 _2739_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_59_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_378 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1877__A _3300_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_60 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2501__A _2566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_25_net107_A _3436_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1962_ _2003_/B _1962_/B _2019_/B _1995_/C vssd1 vssd1 vccd1 vccd1 _1963_/B sky130_fd_sc_hd__or4_1
X_1893_ _3414_/Q _1893_/B vssd1 vssd1 vccd1 vccd1 _1894_/B sky130_fd_sc_hd__xnor2_1
X_3563_ _3564_/CLK _3563_/D _3289_/Y vssd1 vssd1 vccd1 vccd1 _3563_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_37_net107 _3494_/CLK vssd1 vssd1 vccd1 vccd1 _3322_/CLK sky130_fd_sc_hd__clkbuf_16
X_2514_ _2552_/A _3006_/A vssd1 vssd1 vccd1 vccd1 _2996_/A sky130_fd_sc_hd__nor2_1
X_3494_ _3494_/CLK _3494_/D vssd1 vssd1 vccd1 vccd1 _3494_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2130__B _2389_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2445_ _3313_/Q _2425_/X _2441_/X _2444_/X vssd1 vssd1 vccd1 vccd1 _3313_/D sky130_fd_sc_hd__o211a_1
XFILLER_84_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2376_ _3282_/A vssd1 vssd1 vccd1 vccd1 _2376_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_29_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1697__A _2026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_540 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_576 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2038__A_N _2206_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2230_ _2215_/Y _1922_/X _2229_/Y vssd1 vssd1 vccd1 vccd1 _2230_/X sky130_fd_sc_hd__o21a_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_462 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2161_ _2161_/A _2161_/B vssd1 vssd1 vccd1 vccd1 _2162_/B sky130_fd_sc_hd__xnor2_1
XFILLER_65_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2092_ _2092_/A _2092_/B vssd1 vssd1 vccd1 vccd1 _2093_/D sky130_fd_sc_hd__xnor2_1
XFILLER_0_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_576 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2994_ _3357_/Q _2979_/B _2985_/C _3453_/Q vssd1 vssd1 vccd1 vccd1 _2994_/X sky130_fd_sc_hd__a22o_1
XANTENNA__2125__B _2295_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1945_ _2011_/A _2015_/B _1945_/C vssd1 vssd1 vccd1 vccd1 _1945_/X sky130_fd_sc_hd__and3_1
X_1876_ _3420_/Q vssd1 vssd1 vccd1 vccd1 _1876_/Y sky130_fd_sc_hd__inv_2
X_3546_ _3546_/D _2362_/X vssd1 vssd1 vccd1 vccd1 _3548_/D sky130_fd_sc_hd__dlxtn_1
XANTENNA__2141__A _3361_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3477_ _3529_/CLK _3477_/D vssd1 vssd1 vccd1 vccd1 _3477_/Q sky130_fd_sc_hd__dfxtp_1
X_2428_ _2468_/B vssd1 vssd1 vccd1 vccd1 _2441_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_84_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2359_ _3543_/Q _3544_/Q vssd1 vssd1 vccd1 vccd1 _2360_/A sky130_fd_sc_hd__and2_1
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2035__B _2106_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2051__A _3348_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_20_net107 clkbuf_2_3__f_net107/X vssd1 vssd1 vccd1 vccd1 _3414_/CLK sky130_fd_sc_hd__clkbuf_16
Xrlbp_macro_231 vssd1 vssd1 vccd1 vccd1 rlbp_macro_231/HI la_data_out[33] sky130_fd_sc_hd__conb_1
Xrlbp_macro_242 vssd1 vssd1 vccd1 vccd1 rlbp_macro_242/HI la_data_out[44] sky130_fd_sc_hd__conb_1
Xrlbp_macro_220 vssd1 vssd1 vccd1 vccd1 rlbp_macro_220/HI la_data_out[22] sky130_fd_sc_hd__conb_1
XFILLER_0_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrlbp_macro_275 vssd1 vssd1 vccd1 vccd1 rlbp_macro_275/HI la_data_out[77] sky130_fd_sc_hd__conb_1
Xrlbp_macro_253 vssd1 vssd1 vccd1 vccd1 rlbp_macro_253/HI la_data_out[55] sky130_fd_sc_hd__conb_1
Xrlbp_macro_264 vssd1 vssd1 vccd1 vccd1 rlbp_macro_264/HI la_data_out[66] sky130_fd_sc_hd__conb_1
XFILLER_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input34_A la_data_in[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrlbp_macro_297 vssd1 vssd1 vccd1 vccd1 rlbp_macro_297/HI la_data_out[99] sky130_fd_sc_hd__conb_1
Xrlbp_macro_286 vssd1 vssd1 vccd1 vccd1 rlbp_macro_286/HI la_data_out[88] sky130_fd_sc_hd__conb_1
XFILLER_47_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1730_ _2373_/A _2378_/A vssd1 vssd1 vccd1 vccd1 _2375_/A sky130_fd_sc_hd__and2b_1
XFILLER_7_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1661_ _3508_/Q _2405_/A vssd1 vssd1 vccd1 vccd1 _1661_/X sky130_fd_sc_hd__xor2_1
X_3400_ _3400_/CLK _3400_/D vssd1 vssd1 vccd1 vccd1 _3400_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_98_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3331_ _3486_/CLK _3331_/D vssd1 vssd1 vccd1 vccd1 _3331_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3262_ _3527_/Q _3262_/B _3262_/C vssd1 vssd1 vccd1 vccd1 _3262_/X sky130_fd_sc_hd__or3_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_518 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2213_ _2213_/A _2213_/B _2233_/B _2213_/D vssd1 vssd1 vccd1 vccd1 _2213_/X sky130_fd_sc_hd__and4_1
XFILLER_78_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3193_ _3193_/A _3202_/B vssd1 vssd1 vccd1 vccd1 _3193_/Y sky130_fd_sc_hd__nand2_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2144_ _2141_/X _2142_/X _2143_/X vssd1 vssd1 vccd1 vccd1 _2144_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_38_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2075_ _2074_/B _2074_/C _3333_/Q vssd1 vssd1 vccd1 vccd1 _2075_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_53_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_370 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_468 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3092__B2 _3411_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3092__A1 _3327_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2977_ _2977_/A _2977_/B vssd1 vssd1 vccd1 vccd1 _2977_/X sky130_fd_sc_hd__or2_1
X_1928_ _1928_/A _1928_/B vssd1 vssd1 vccd1 vccd1 _1929_/B sky130_fd_sc_hd__xor2_1
X_1859_ _3424_/Q _2309_/A vssd1 vssd1 vccd1 vccd1 _1860_/B sky130_fd_sc_hd__and2b_1
XFILLER_1_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3529_ _3529_/CLK _3529_/D vssd1 vssd1 vccd1 vccd1 _3529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_240 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_402 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1869__B _2292_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2046__A _3345_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1779__B _2292_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2900_ _3450_/Q _2888_/X _2899_/X _2895_/X vssd1 vssd1 vccd1 vccd1 _3450_/D sky130_fd_sc_hd__o211a_1
XFILLER_45_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2831_ _3199_/A vssd1 vssd1 vccd1 vccd1 _2895_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__1795__A _3445_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2762_ _2762_/A _2765_/B vssd1 vssd1 vccd1 vccd1 _2762_/X sky130_fd_sc_hd__or2_1
X_1713_ _3497_/Q _2118_/B _1673_/Y _3494_/Q vssd1 vssd1 vccd1 vccd1 _1719_/B sky130_fd_sc_hd__a2bb2o_1
X_2693_ _2707_/B vssd1 vssd1 vccd1 vccd1 _2703_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__3129__A2 _3036_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1644_ _1774_/B vssd1 vssd1 vccd1 vccd1 _2405_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_98_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1713__A2_N _2118_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3314_ _3491_/CLK _3314_/D vssd1 vssd1 vccd1 vccd1 _3314_/Q sky130_fd_sc_hd__dfxtp_1
X_3245_ _3262_/B vssd1 vssd1 vccd1 vccd1 _3256_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_58_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3176_ _3494_/Q _3173_/X _3175_/X _3171_/X vssd1 vssd1 vccd1 vccd1 _3494_/D sky130_fd_sc_hd__o211a_1
XFILLER_39_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2127_ _2191_/B _3360_/Q vssd1 vssd1 vccd1 vccd1 _2129_/A sky130_fd_sc_hd__and2b_1
XFILLER_66_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2058_ _2057_/Y _2405_/A _2040_/B vssd1 vssd1 vccd1 vccd1 _2058_/X sky130_fd_sc_hd__o21a_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3065__A1 _3325_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3065__B2 _3409_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2313__B _2313_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_295 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3160__A _3160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput70 _3779_/X vssd1 vssd1 vccd1 vccd1 OTA_sh_c sky130_fd_sc_hd__buf_2
Xoutput81 _3790_/X vssd1 vssd1 vccd1 vccd1 Pd3_a sky130_fd_sc_hd__buf_2
Xoutput92 _3801_/X vssd1 vssd1 vccd1 vccd1 Pd8_b sky130_fd_sc_hd__buf_2
XFILLER_95_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_2_net107_A _3494_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3030_ _3199_/A vssd1 vssd1 vccd1 vccd1 _3184_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_63_210 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_295 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2270__A2 _2213_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2814_ _2966_/A _2824_/B vssd1 vssd1 vccd1 vccd1 _2814_/X sky130_fd_sc_hd__or2_1
X_3794_ _3794_/A vssd1 vssd1 vccd1 vccd1 _3794_/X sky130_fd_sc_hd__clkbuf_1
X_2745_ _2782_/A _2745_/B vssd1 vssd1 vccd1 vccd1 _2745_/X sky130_fd_sc_hd__or2_1
XFILLER_11_18 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2676_ _2676_/A vssd1 vssd1 vccd1 vccd1 _2679_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__3245__A _3262_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3228_ _3251_/A vssd1 vssd1 vccd1 vccd1 _3228_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1836__A2 _1834_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3159_ _3173_/A vssd1 vssd1 vccd1 vccd1 _3159_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3038__A1 _3359_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3038__B2 _3455_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_184 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2043__B _2291_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3201__A1 _2563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2530_ _3336_/Q _2518_/X _2529_/X _2523_/X vssd1 vssd1 vccd1 vccd1 _3336_/D sky130_fd_sc_hd__o211a_1
X_2461_ _2582_/A _2461_/B vssd1 vssd1 vccd1 vccd1 _2461_/X sky130_fd_sc_hd__or2_1
X_2392_ _2395_/B _2395_/C vssd1 vssd1 vccd1 vccd1 _2394_/A sky130_fd_sc_hd__and2_1
XFILLER_68_324 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_519 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3013_ _3477_/Q _2990_/X _3012_/X _2971_/X vssd1 vssd1 vccd1 vccd1 _3477_/D sky130_fd_sc_hd__o211a_1
XANTENNA__2128__B _2191_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1967__B _2301_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2728_ _2728_/A vssd1 vssd1 vccd1 vccd1 _2728_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2659_ _3374_/Q _2656_/X _2658_/X _2654_/X vssd1 vssd1 vccd1 vccd1 _3374_/D sky130_fd_sc_hd__o211a_1
XFILLER_86_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_454 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3259__A1 _3526_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2038__B _3351_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3533_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input64_A wbs_sel_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2305__B_N _1794_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_460 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1961_ _3309_/Q _2046_/B vssd1 vssd1 vccd1 vccd1 _1995_/C sky130_fd_sc_hd__nor2_1
X_1892_ _1911_/A _1911_/B _1851_/A vssd1 vssd1 vccd1 vccd1 _1894_/A sky130_fd_sc_hd__a21o_1
XANTENNA__2899__A _2973_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3562_ _3562_/D _2368_/X vssd1 vssd1 vccd1 vccd1 _3564_/D sky130_fd_sc_hd__dlxtn_1
X_2513_ _2513_/A vssd1 vssd1 vccd1 vccd1 _3006_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_5_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3493_ _3511_/CLK _3493_/D vssd1 vssd1 vccd1 vccd1 _3493_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2444_ _3264_/A vssd1 vssd1 vccd1 vccd1 _2444_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2375_ _2375_/A vssd1 vssd1 vccd1 vccd1 _3282_/A sky130_fd_sc_hd__buf_2
XFILLER_83_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1972__B_N _2105_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_552 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1888__A _2145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_588 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1718__A1 _3489_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2160_ _2160_/A _2160_/B vssd1 vssd1 vccd1 vccd1 _2167_/A sky130_fd_sc_hd__xnor2_1
XFILLER_78_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2091_ _3340_/Q _2091_/B vssd1 vssd1 vccd1 vccd1 _2092_/B sky130_fd_sc_hd__xnor2_1
XFILLER_38_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2993_ _2993_/A vssd1 vssd1 vccd1 vccd1 _2993_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1944_ _1988_/A _1991_/B vssd1 vssd1 vccd1 vccd1 _1945_/C sky130_fd_sc_hd__and2_1
XFILLER_9_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1875_ _1875_/A vssd1 vssd1 vccd1 vccd1 _3536_/D sky130_fd_sc_hd__clkbuf_1
X_3545_ _3545_/D _2362_/X vssd1 vssd1 vccd1 vccd1 _3545_/Q sky130_fd_sc_hd__dlxtn_1
X_3476_ _3476_/CLK _3476_/D vssd1 vssd1 vccd1 vccd1 _3476_/Q sky130_fd_sc_hd__dfxtp_1
X_2427_ _2427_/A _2834_/A vssd1 vssd1 vccd1 vccd1 _2468_/B sky130_fd_sc_hd__or2b_1
XFILLER_69_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2358_ _2358_/A vssd1 vssd1 vccd1 vccd1 _2358_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_84_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2289_ _2289_/A _2289_/B vssd1 vssd1 vccd1 vccd1 _2343_/A sky130_fd_sc_hd__nor2_1
XFILLER_84_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_127 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_547 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrlbp_macro_210 vssd1 vssd1 vccd1 vccd1 rlbp_macro_210/HI la_data_out[12] sky130_fd_sc_hd__conb_1
Xrlbp_macro_232 vssd1 vssd1 vccd1 vccd1 rlbp_macro_232/HI la_data_out[34] sky130_fd_sc_hd__conb_1
Xrlbp_macro_221 vssd1 vssd1 vccd1 vccd1 rlbp_macro_221/HI la_data_out[23] sky130_fd_sc_hd__conb_1
Xrlbp_macro_243 vssd1 vssd1 vccd1 vccd1 rlbp_macro_243/HI la_data_out[45] sky130_fd_sc_hd__conb_1
Xrlbp_macro_254 vssd1 vssd1 vccd1 vccd1 rlbp_macro_254/HI la_data_out[56] sky130_fd_sc_hd__conb_1
Xrlbp_macro_265 vssd1 vssd1 vccd1 vccd1 rlbp_macro_265/HI la_data_out[67] sky130_fd_sc_hd__conb_1
Xrlbp_macro_276 vssd1 vssd1 vccd1 vccd1 rlbp_macro_276/HI la_data_out[78] sky130_fd_sc_hd__conb_1
XFILLER_85_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrlbp_macro_287 vssd1 vssd1 vccd1 vccd1 rlbp_macro_287/HI la_data_out[89] sky130_fd_sc_hd__conb_1
Xrlbp_macro_298 vssd1 vssd1 vccd1 vccd1 rlbp_macro_298/HI la_data_out[100] sky130_fd_sc_hd__conb_1
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input27_A la_data_in[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2507__A _2584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1660_ _2037_/B vssd1 vssd1 vccd1 vccd1 _2405_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__1784__C _1840_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output95_A _3804_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3330_ _3332_/CLK _3330_/D vssd1 vssd1 vccd1 vccd1 _3330_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3261_ _3527_/Q _1707_/A _3251_/X _3260_/X vssd1 vssd1 vccd1 vccd1 _3527_/D sky130_fd_sc_hd__o211a_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2212_ _2212_/A _2212_/B _2267_/A _2251_/C vssd1 vssd1 vccd1 vccd1 _2213_/D sky130_fd_sc_hd__and4_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3192_ _3207_/A vssd1 vssd1 vccd1 vccd1 _3202_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_2143_ _1796_/X _3362_/Q vssd1 vssd1 vccd1 vccd1 _2143_/X sky130_fd_sc_hd__and2b_1
XANTENNA__3801__A _3801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2074_ _3333_/Q _2074_/B _2074_/C vssd1 vssd1 vccd1 vccd1 _2074_/X sky130_fd_sc_hd__and3_1
XFILLER_53_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2136__B _2389_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1975__B _3314_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2976_ _3475_/Q _2962_/A _2975_/X _2971_/X vssd1 vssd1 vccd1 vccd1 _3475_/D sky130_fd_sc_hd__o211a_1
X_1927_ _1927_/A _1927_/B vssd1 vssd1 vccd1 vccd1 _1930_/C sky130_fd_sc_hd__xnor2_1
X_1858_ _2145_/A _3424_/Q vssd1 vssd1 vccd1 vccd1 _1860_/A sky130_fd_sc_hd__and2b_1
XFILLER_89_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1789_ _3442_/Q _2389_/B vssd1 vssd1 vccd1 vccd1 _1789_/X sky130_fd_sc_hd__and2b_1
XANTENNA__1991__A _3326_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3528_ _3528_/CLK _3528_/D vssd1 vssd1 vccd1 vccd1 _3528_/Q sky130_fd_sc_hd__dfxtp_1
X_3459_ _3462_/CLK _3459_/D vssd1 vssd1 vccd1 vccd1 _3459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_400 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_127 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2327__A _3456_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2046__B _2046_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3158__A _3158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2997__A _2997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_2_1__f_net107 clkbuf_0_net107/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_9_net107/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_48_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_6 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2830_ _2977_/A _2830_/B vssd1 vssd1 vccd1 vccd1 _2830_/X sky130_fd_sc_hd__or2_1
XFILLER_31_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2761_ _3407_/Q _2753_/X _2760_/X _2743_/X vssd1 vssd1 vccd1 vccd1 _3407_/D sky130_fd_sc_hd__o211a_1
XFILLER_31_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2692_ _2692_/A vssd1 vssd1 vccd1 vccd1 _2692_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1712_ _1757_/A vssd1 vssd1 vccd1 vccd1 _2118_/B sky130_fd_sc_hd__buf_2
XANTENNA__2585__A1 _3355_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1643_ _3303_/Q vssd1 vssd1 vccd1 vccd1 _1774_/B sky130_fd_sc_hd__buf_2
XANTENNA__2337__A1 _3454_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3313_ _3322_/CLK _3313_/D vssd1 vssd1 vccd1 vccd1 _3313_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3244_ _3528_/Q _3224_/A _3243_/X _3239_/X vssd1 vssd1 vccd1 vccd1 _3520_/D sky130_fd_sc_hd__o211a_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3175_ _3238_/A _3183_/B vssd1 vssd1 vccd1 vccd1 _3175_/X sky130_fd_sc_hd__or2_1
XFILLER_81_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2126_ _3368_/Q _2294_/B vssd1 vssd1 vccd1 vccd1 _2183_/B sky130_fd_sc_hd__xor2_1
X_2057_ _3352_/Q vssd1 vssd1 vccd1 vccd1 _2057_/Y sky130_fd_sc_hd__inv_2
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2959_ _3468_/Q _2948_/X _2957_/X _2958_/X vssd1 vssd1 vccd1 vccd1 _3468_/D sky130_fd_sc_hd__o211a_1
XFILLER_41_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2610__A _2765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_528 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2057__A _3352_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3160__B _3160_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1896__A _3409_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2567__A1 _3348_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_19_net107_A clkbuf_2_3__f_net107/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2319__A1 _2339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2520__A _2679_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput82 _3791_/X vssd1 vssd1 vccd1 vccd1 Pd3_b sky130_fd_sc_hd__buf_2
Xoutput93 _3802_/X vssd1 vssd1 vccd1 vccd1 Pd9_a sky130_fd_sc_hd__buf_2
Xoutput71 _3780_/X vssd1 vssd1 vccd1 vccd1 Pd10_a sky130_fd_sc_hd__buf_2
XANTENNA_hold5_A hold5/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_288 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_182 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2813_ _3241_/A vssd1 vssd1 vccd1 vccd1 _2966_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_31_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3793_ _3793_/A vssd1 vssd1 vccd1 vccd1 _3793_/X sky130_fd_sc_hd__clkbuf_1
X_2744_ _3403_/Q _2728_/A _2741_/X _2743_/X vssd1 vssd1 vccd1 vccd1 _3403_/D sky130_fd_sc_hd__o211a_1
X_2675_ _3053_/A vssd1 vssd1 vccd1 vccd1 _2676_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_98_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3227_ _3227_/A _3236_/B vssd1 vssd1 vccd1 vccd1 _3227_/X sky130_fd_sc_hd__or2_1
XFILLER_67_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3158_ _3158_/A _3160_/B vssd1 vssd1 vccd1 vccd1 _3173_/A sky130_fd_sc_hd__and2_1
XFILLER_94_391 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2109_ _3364_/Q _2309_/A vssd1 vssd1 vccd1 vccd1 _2110_/B sky130_fd_sc_hd__and2b_1
XFILLER_15_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3089_ _3387_/Q _2676_/A _3033_/A _3527_/Q vssd1 vssd1 vccd1 vccd1 _3089_/X sky130_fd_sc_hd__a22o_1
XFILLER_54_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _1748_/A0 sky130_fd_sc_hd__clkbuf_16
XANTENNA__3038__A2 _3036_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2340__A _3461_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2721__A1 _3394_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2460_ _3183_/A vssd1 vssd1 vccd1 vccd1 _2582_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_96_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2391_ _2395_/C _2391_/B vssd1 vssd1 vccd1 vccd1 _3299_/D sky130_fd_sc_hd__nor2_1
XFILLER_3_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3012_ _3012_/A _3012_/B vssd1 vssd1 vccd1 vccd1 _3012_/X sky130_fd_sc_hd__or2_1
XFILLER_91_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_7_net107 clkbuf_leaf_9_net107/A vssd1 vssd1 vccd1 vccd1 _3520_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_20_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2727_ _3397_/Q _2713_/X _2726_/X _2718_/X vssd1 vssd1 vccd1 vccd1 _3397_/D sky130_fd_sc_hd__o211a_1
XANTENNA__3256__A _3524_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2658_ _2769_/A _2666_/B vssd1 vssd1 vccd1 vccd1 _2658_/X sky130_fd_sc_hd__or2_1
X_2589_ _2983_/A _2709_/B vssd1 vssd1 vccd1 vccd1 _2979_/B sky130_fd_sc_hd__nor2_1
XFILLER_101_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input1_A CMP vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_556 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2054__B _2190_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2942__A1 _3464_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3166__A _3232_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input57_A wbs_dat_i[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2229__B _2313_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_34_net107_A _3494_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1960_ _3320_/Q _2294_/B vssd1 vssd1 vccd1 vccd1 _2019_/B sky130_fd_sc_hd__xor2_1
X_1891_ _1873_/B _1895_/B _1890_/X vssd1 vssd1 vccd1 vccd1 _1911_/B sky130_fd_sc_hd__a21o_1
XFILLER_41_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3561_ _3561_/D _2368_/X vssd1 vssd1 vccd1 vccd1 _3563_/D sky130_fd_sc_hd__dlxtn_1
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2512_ _2512_/A _2512_/B _2512_/C _2551_/A vssd1 vssd1 vccd1 vccd1 _2513_/A sky130_fd_sc_hd__or4_1
X_3492_ _3511_/CLK _3492_/D vssd1 vssd1 vccd1 vccd1 _3492_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3804__A _3804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2443_ _3199_/A vssd1 vssd1 vccd1 vccd1 _3264_/A sky130_fd_sc_hd__buf_2
XFILLER_68_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2374_ _3281_/A vssd1 vssd1 vccd1 vccd1 _2374_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_68_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2061__A_N _1974_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2924__A1 _3457_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2049__B _2049_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3101__A1 _3328_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_564 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3101__B2 _3412_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_372 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1718__A2 _2295_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1797__B_N _1796_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2090_ _2087_/A _2087_/B _2040_/B vssd1 vssd1 vccd1 vccd1 _2092_/A sky130_fd_sc_hd__a21oi_1
XFILLER_17_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1798__B _3446_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2992_ _3155_/A vssd1 vssd1 vccd1 vccd1 _3012_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_34_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1943_ _3314_/Q _3302_/Q vssd1 vssd1 vccd1 vccd1 _1991_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__2703__A _2778_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1874_ _1874_/A _1874_/B vssd1 vssd1 vccd1 vccd1 _1875_/A sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_0_net107_A _1749_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3544_ _3544_/CLK _3544_/D _3279_/Y vssd1 vssd1 vccd1 vccd1 _3544_/Q sky130_fd_sc_hd__dfrtp_1
X_3475_ _3476_/CLK _3475_/D vssd1 vssd1 vccd1 vccd1 _3475_/Q sky130_fd_sc_hd__dfxtp_1
X_2426_ _3227_/A vssd1 vssd1 vccd1 vccd1 _2559_/A sky130_fd_sc_hd__buf_2
XFILLER_57_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2357_ _3539_/Q _3538_/Q vssd1 vssd1 vccd1 vccd1 _2358_/A sky130_fd_sc_hd__and2_1
XFILLER_84_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2288_ _3471_/Q _2288_/B vssd1 vssd1 vccd1 vccd1 _2289_/B sky130_fd_sc_hd__and2b_1
XANTENNA__1989__A _3325_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2613__A _3238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrlbp_macro_200 vssd1 vssd1 vccd1 vccd1 rlbp_macro_200/HI la_data_out[2] sky130_fd_sc_hd__conb_1
Xrlbp_macro_211 vssd1 vssd1 vccd1 vccd1 rlbp_macro_211/HI la_data_out[13] sky130_fd_sc_hd__conb_1
Xrlbp_macro_233 vssd1 vssd1 vccd1 vccd1 rlbp_macro_233/HI la_data_out[35] sky130_fd_sc_hd__conb_1
Xrlbp_macro_222 vssd1 vssd1 vccd1 vccd1 rlbp_macro_222/HI la_data_out[24] sky130_fd_sc_hd__conb_1
Xrlbp_macro_244 vssd1 vssd1 vccd1 vccd1 rlbp_macro_244/HI la_data_out[46] sky130_fd_sc_hd__conb_1
Xrlbp_macro_255 vssd1 vssd1 vccd1 vccd1 rlbp_macro_255/HI la_data_out[57] sky130_fd_sc_hd__conb_1
Xrlbp_macro_266 vssd1 vssd1 vccd1 vccd1 rlbp_macro_266/HI la_data_out[68] sky130_fd_sc_hd__conb_1
XFILLER_94_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrlbp_macro_277 vssd1 vssd1 vccd1 vccd1 rlbp_macro_277/HI la_data_out[79] sky130_fd_sc_hd__conb_1
Xrlbp_macro_288 vssd1 vssd1 vccd1 vccd1 rlbp_macro_288/HI la_data_out[90] sky130_fd_sc_hd__conb_1
Xrlbp_macro_299 vssd1 vssd1 vccd1 vccd1 rlbp_macro_299/HI la_data_out[101] sky130_fd_sc_hd__conb_1
XFILLER_90_404 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2523__A _2566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3260_ _3526_/Q _3262_/B _3262_/C vssd1 vssd1 vccd1 vccd1 _3260_/X sky130_fd_sc_hd__or3_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2211_ _3393_/Q _2295_/B vssd1 vssd1 vccd1 vccd1 _2251_/C sky130_fd_sc_hd__or2_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3191_ _3207_/A vssd1 vssd1 vccd1 vccd1 _3191_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2142_ _3362_/Q _1796_/X vssd1 vssd1 vccd1 vccd1 _2142_/X sky130_fd_sc_hd__or2b_1
XFILLER_15_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2073_ _2073_/A _2074_/B vssd1 vssd1 vccd1 vccd1 _2073_/Y sky130_fd_sc_hd__xnor2_1
X_2975_ _2975_/A _2977_/B vssd1 vssd1 vccd1 vccd1 _2975_/X sky130_fd_sc_hd__or2_1
X_1926_ _3416_/Q _1926_/B vssd1 vssd1 vccd1 vccd1 _1927_/B sky130_fd_sc_hd__xnor2_1
XFILLER_30_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1857_ _1895_/A _1898_/B vssd1 vssd1 vccd1 vccd1 _1865_/A sky130_fd_sc_hd__and2_1
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3527_ _3528_/CLK _3527_/D vssd1 vssd1 vccd1 vccd1 _3527_/Q sky130_fd_sc_hd__dfxtp_1
X_1788_ _3444_/Q vssd1 vssd1 vccd1 vccd1 _1788_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3264__A _3264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3458_ _3474_/CLK _3458_/D vssd1 vssd1 vccd1 vccd1 _3458_/Q sky130_fd_sc_hd__dfxtp_1
X_3389_ _3392_/CLK _3389_/D vssd1 vssd1 vccd1 vccd1 _3389_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_57_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2409_ _2407_/A _2407_/B _2408_/Y _2397_/X vssd1 vssd1 vccd1 vccd1 _3305_/D sky130_fd_sc_hd__o211a_1
XFILLER_29_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1967__A_N _3310_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3158__B _3160_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_492 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2760_ _2760_/A _2765_/B vssd1 vssd1 vccd1 vccd1 _2760_/X sky130_fd_sc_hd__or2_1
XFILLER_12_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2691_ _3385_/Q _2678_/X _2690_/X _2686_/X vssd1 vssd1 vccd1 vccd1 _3385_/D sky130_fd_sc_hd__o211a_1
X_1711_ _3499_/Q _1654_/A _1657_/Y _3492_/Q _1710_/X vssd1 vssd1 vccd1 vccd1 _1719_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_6_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3312_ _3322_/CLK _3312_/D vssd1 vssd1 vccd1 vccd1 _3312_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3243_ _3243_/A _3243_/B vssd1 vssd1 vccd1 vccd1 _3243_/X sky130_fd_sc_hd__or2_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3174_ _3188_/B vssd1 vssd1 vccd1 vccd1 _3183_/B sky130_fd_sc_hd__clkbuf_1
X_2125_ _3357_/Q _2295_/B vssd1 vssd1 vccd1 vccd1 _2125_/Y sky130_fd_sc_hd__nor2_1
XFILLER_81_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2056_ _2051_/Y _1878_/X _2033_/C _2080_/B _2055_/X vssd1 vssd1 vccd1 vccd1 _2068_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_54_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2958_ _2971_/A vssd1 vssd1 vccd1 vccd1 _2958_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1909_ _3406_/Q _1900_/Y _1903_/Y _1906_/Y _1908_/Y vssd1 vssd1 vccd1 vccd1 _1910_/D
+ sky130_fd_sc_hd__o2111ai_1
X_2889_ _2903_/B vssd1 vssd1 vccd1 vccd1 _2899_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_89_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3289__B1 _3282_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_407 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2972__C1 _2971_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput83 _3792_/X vssd1 vssd1 vccd1 vccd1 Pd4_a sky130_fd_sc_hd__buf_2
Xoutput94 _3803_/X vssd1 vssd1 vccd1 vccd1 Pd9_b sky130_fd_sc_hd__buf_2
Xoutput72 _3781_/X vssd1 vssd1 vccd1 vccd1 Pd10_b sky130_fd_sc_hd__buf_2
XFILLER_95_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_256 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3792_ _3792_/A vssd1 vssd1 vccd1 vccd1 _3792_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2812_ _3422_/Q _2808_/X _2811_/X _2797_/X vssd1 vssd1 vccd1 vccd1 _3422_/D sky130_fd_sc_hd__o211a_1
X_2743_ _2815_/A vssd1 vssd1 vccd1 vccd1 _2743_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2711__A _2711_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2674_ _3006_/A _2709_/B vssd1 vssd1 vccd1 vccd1 _3053_/A sky130_fd_sc_hd__nor2_1
XFILLER_101_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3226_ _3243_/B vssd1 vssd1 vccd1 vccd1 _3236_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_67_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3157_ _3488_/Q _3074_/A _3155_/X _3156_/X vssd1 vssd1 vccd1 vccd1 _3488_/D sky130_fd_sc_hd__o211a_1
XFILLER_27_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2108_ _2309_/A _3364_/Q vssd1 vssd1 vccd1 vccd1 _2110_/A sky130_fd_sc_hd__and2b_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1997__A _3324_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3088_ _3423_/Q _2787_/A _2946_/A _3471_/Q _3087_/X vssd1 vssd1 vccd1 vccd1 _3088_/X
+ sky130_fd_sc_hd__a221o_1
X_2039_ _3351_/Q _2288_/B vssd1 vssd1 vccd1 vccd1 _2040_/B sky130_fd_sc_hd__and2b_1
XFILLER_35_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_495 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2621__A _3243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2485__A1 _3322_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3131__C1 _3130_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_204 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1700__A _2389_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_26_net107 _3436_/CLK vssd1 vssd1 vccd1 vccd1 _3464_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_41_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2531__A _2568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2390_ _1667_/X _2385_/X _2397_/A vssd1 vssd1 vccd1 vccd1 _2391_/B sky130_fd_sc_hd__o21ai_1
XFILLER_3_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3011_ _3309_/Q _2993_/X _3005_/X _3010_/X vssd1 vssd1 vccd1 vccd1 _3012_/B sky130_fd_sc_hd__a211o_1
XFILLER_36_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2726_ _2765_/A _2726_/B vssd1 vssd1 vccd1 vccd1 _2726_/X sky130_fd_sc_hd__or2_1
XANTENNA__2441__A _2568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2657_ _2672_/B vssd1 vssd1 vccd1 vccd1 _2666_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__2059__B_N _1794_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2588_ _2982_/A _2982_/C _2905_/B _2982_/B vssd1 vssd1 vccd1 vccd1 _2709_/B sky130_fd_sc_hd__or4b_2
XFILLER_99_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3209_ _2572_/A _3207_/X _3208_/Y _3200_/X vssd1 vssd1 vccd1 vccd1 _3506_/D sky130_fd_sc_hd__o211a_1
XFILLER_55_543 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_568 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_59 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_292 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3544__RESET_B _3279_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2351__A _3463_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1902__B1 _3405_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1890_ _1918_/B _1914_/A _1887_/Y _1889_/X vssd1 vssd1 vccd1 vccd1 _1890_/X sky130_fd_sc_hd__a31o_1
X_3560_ _3560_/D _2368_/X vssd1 vssd1 vccd1 vccd1 _3560_/Q sky130_fd_sc_hd__dlxtn_1
X_2511_ _2511_/A vssd1 vssd1 vccd1 vccd1 _2551_/A sky130_fd_sc_hd__inv_2
XFILLER_5_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3491_ _3491_/CLK _3491_/D vssd1 vssd1 vccd1 vccd1 _3491_/Q sky130_fd_sc_hd__dfxtp_1
X_2442_ _2442_/A vssd1 vssd1 vccd1 vccd1 _3199_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_45_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2373_ _2373_/A vssd1 vssd1 vccd1 vccd1 _3281_/A sky130_fd_sc_hd__buf_2
XFILLER_83_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2709_ _3002_/A _2709_/B vssd1 vssd1 vccd1 vccd1 _3041_/A sky130_fd_sc_hd__nor2_1
XFILLER_99_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_576 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_395 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2860__A1 _3436_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_398 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3177__A _3241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2991_ _2427_/A _2988_/A _3264_/B vssd1 vssd1 vccd1 vccd1 _3155_/A sky130_fd_sc_hd__a21bo_1
XFILLER_61_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1942_ _3313_/Q _2281_/B vssd1 vssd1 vccd1 vccd1 _1988_/A sky130_fd_sc_hd__xnor2_1
X_1873_ _1873_/A _1873_/B _1926_/B _1873_/D vssd1 vssd1 vccd1 vccd1 _1874_/B sky130_fd_sc_hd__nand4_1
X_3543_ _3544_/CLK _3543_/D _3278_/Y vssd1 vssd1 vccd1 vccd1 _3543_/Q sky130_fd_sc_hd__dfrtp_1
X_3474_ _3474_/CLK _3474_/D vssd1 vssd1 vccd1 vccd1 _3474_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2425_ _2446_/A vssd1 vssd1 vccd1 vccd1 _2425_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_clkbuf_0_wb_clk_i_A wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2356_ _2356_/A vssd1 vssd1 vccd1 vccd1 _2356_/X sky130_fd_sc_hd__clkbuf_1
X_2287_ _2206_/B _3471_/Q vssd1 vssd1 vccd1 vccd1 _2289_/A sky130_fd_sc_hd__and2b_1
XFILLER_29_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2166__A _3369_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrlbp_macro_212 vssd1 vssd1 vccd1 vccd1 rlbp_macro_212/HI la_data_out[14] sky130_fd_sc_hd__conb_1
Xrlbp_macro_223 vssd1 vssd1 vccd1 vccd1 rlbp_macro_223/HI la_data_out[25] sky130_fd_sc_hd__conb_1
Xrlbp_macro_201 vssd1 vssd1 vccd1 vccd1 rlbp_macro_201/HI la_data_out[3] sky130_fd_sc_hd__conb_1
Xrlbp_macro_234 vssd1 vssd1 vccd1 vccd1 rlbp_macro_234/HI la_data_out[36] sky130_fd_sc_hd__conb_1
Xrlbp_macro_245 vssd1 vssd1 vccd1 vccd1 rlbp_macro_245/HI la_data_out[47] sky130_fd_sc_hd__conb_1
Xrlbp_macro_256 vssd1 vssd1 vccd1 vccd1 rlbp_macro_256/HI la_data_out[58] sky130_fd_sc_hd__conb_1
Xrlbp_macro_267 vssd1 vssd1 vccd1 vccd1 rlbp_macro_267/HI la_data_out[69] sky130_fd_sc_hd__conb_1
Xrlbp_macro_289 vssd1 vssd1 vccd1 vccd1 rlbp_macro_289/HI la_data_out[91] sky130_fd_sc_hd__conb_1
Xrlbp_macro_278 vssd1 vssd1 vccd1 vccd1 rlbp_macro_278/HI la_data_out[80] sky130_fd_sc_hd__conb_1
XFILLER_87_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3010__A1 _3321_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3010__B2 _3405_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2210_ _2210_/A _2210_/B vssd1 vssd1 vccd1 vccd1 _2267_/A sky130_fd_sc_hd__nor2_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3190_ _3225_/A _3195_/B vssd1 vssd1 vccd1 vccd1 _3207_/A sky130_fd_sc_hd__nand2_1
X_2141_ _3361_/Q _1794_/X vssd1 vssd1 vccd1 vccd1 _2141_/X sky130_fd_sc_hd__or2b_1
XFILLER_38_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2072_ _2072_/A _2072_/B vssd1 vssd1 vccd1 vccd1 _2083_/C sky130_fd_sc_hd__xnor2_1
XFILLER_81_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3077__B2 _3526_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_376 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1769__A_N _2145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2974_ _3474_/Q _2962_/X _2973_/X _2971_/X vssd1 vssd1 vccd1 vccd1 _3474_/D sky130_fd_sc_hd__o211a_1
X_1925_ _1928_/A _1928_/B _1870_/A vssd1 vssd1 vccd1 vccd1 _1927_/A sky130_fd_sc_hd__a21oi_1
X_1856_ _3422_/Q _2106_/B vssd1 vssd1 vccd1 vccd1 _1898_/B sky130_fd_sc_hd__xnor2_1
X_1787_ _1787_/A vssd1 vssd1 vccd1 vccd1 _3291_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3001__A1 _3345_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3001__B2 _3429_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3526_ _3528_/CLK _3526_/D vssd1 vssd1 vccd1 vccd1 _3526_/Q sky130_fd_sc_hd__dfxtp_1
X_3457_ _3464_/CLK _3457_/D vssd1 vssd1 vccd1 vccd1 _3457_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3388_ _3392_/CLK _3388_/D vssd1 vssd1 vccd1 vccd1 _3388_/Q sky130_fd_sc_hd__dfxtp_1
X_2408_ _2412_/C vssd1 vssd1 vccd1 vccd1 _2408_/Y sky130_fd_sc_hd__inv_2
X_2339_ _2339_/A _2339_/B vssd1 vssd1 vccd1 vccd1 _2341_/B sky130_fd_sc_hd__xor2_1
XANTENNA__3280__A hold2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3068__B2 _3525_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2624__A _3181_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3240__A1 _3526_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input32_A la_data_in[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3190__A _3225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3231__A1 _3522_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2690_ _2765_/A _2690_/B vssd1 vssd1 vccd1 vccd1 _2690_/X sky130_fd_sc_hd__or2_1
X_1710_ _3496_/Q _2037_/B vssd1 vssd1 vccd1 vccd1 _1710_/X sky130_fd_sc_hd__xor2_1
X_3311_ _3322_/CLK _3311_/D vssd1 vssd1 vccd1 vccd1 _3311_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3242_ _3527_/Q _3224_/A _3241_/X _3239_/X vssd1 vssd1 vccd1 vccd1 _3519_/D sky130_fd_sc_hd__o211a_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3173_ _3173_/A vssd1 vssd1 vccd1 vccd1 _3173_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2709__A _3002_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2124_ _2389_/C _3357_/Q vssd1 vssd1 vccd1 vccd1 _2165_/B sky130_fd_sc_hd__or2b_1
XFILLER_66_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_427 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2055_ _2051_/Y _1698_/A _2054_/X vssd1 vssd1 vccd1 vccd1 _2055_/X sky130_fd_sc_hd__o21a_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2444__A _3264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3222__A1 _2586_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2957_ _2957_/A _2960_/B vssd1 vssd1 vccd1 vccd1 _2957_/X sky130_fd_sc_hd__or2_1
XFILLER_41_18 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1908_ _3407_/Q _1908_/B vssd1 vssd1 vccd1 vccd1 _1908_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__2430__C1 _2370_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2888_ _2888_/A vssd1 vssd1 vccd1 vccd1 _2888_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1839_ _1837_/A _1837_/B _1780_/A vssd1 vssd1 vccd1 vccd1 _1841_/A sky130_fd_sc_hd__a21oi_1
XFILLER_1_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3509_ _3511_/CLK _3509_/D vssd1 vssd1 vccd1 vccd1 _3509_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3289__A1 hold2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_58 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput84 _3793_/X vssd1 vssd1 vccd1 vccd1 Pd4_b sky130_fd_sc_hd__buf_2
Xoutput73 _3782_/X vssd1 vssd1 vccd1 vccd1 Pd11_a sky130_fd_sc_hd__buf_2
XFILLER_95_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput95 _3804_/X vssd1 vssd1 vccd1 vccd1 SH_out_c sky130_fd_sc_hd__buf_2
XFILLER_0_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2529__A _2565_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3791_ _3791_/A vssd1 vssd1 vccd1 vccd1 _3791_/X sky130_fd_sc_hd__clkbuf_1
X_2811_ _2964_/A _2824_/B vssd1 vssd1 vccd1 vccd1 _2811_/X sky130_fd_sc_hd__or2_1
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2742_ _2742_/A vssd1 vssd1 vccd1 vccd1 _2815_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2673_ _3380_/Q _2656_/A _2672_/X _2668_/X vssd1 vssd1 vccd1 vccd1 _3380_/D sky130_fd_sc_hd__o211a_1
X_3225_ _3225_/A _3225_/B vssd1 vssd1 vccd1 vccd1 _3243_/B sky130_fd_sc_hd__nand2_1
XANTENNA__3140__B1 _2595_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3156_ _3184_/A vssd1 vssd1 vccd1 vccd1 _3156_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_27_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2107_ _2155_/A _2153_/B vssd1 vssd1 vccd1 vccd1 _2114_/A sky130_fd_sc_hd__and2_1
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3087_ _3363_/Q _3036_/X _3037_/X _3459_/Q vssd1 vssd1 vccd1 vccd1 _3087_/X sky130_fd_sc_hd__a22o_1
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2038_ _2206_/B _3351_/Q vssd1 vssd1 vccd1 vccd1 _2040_/A sky130_fd_sc_hd__and2b_1
XFILLER_42_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2112__A_N _3363_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_216 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3010_ _3321_/Q _2480_/B _2754_/B _3405_/Q _3009_/X vssd1 vssd1 vccd1 vccd1 _3010_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_64_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1684__B1 _2046_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2722__A _2760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2725_ _3396_/Q _2713_/X _2724_/X _2718_/X vssd1 vssd1 vccd1 vccd1 _3396_/D sky130_fd_sc_hd__o211a_1
X_2656_ _2656_/A vssd1 vssd1 vccd1 vccd1 _2656_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_99_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2587_ _3356_/Q _2570_/A _2586_/X _2580_/X vssd1 vssd1 vccd1 vccd1 _3356_/D sky130_fd_sc_hd__o211a_1
XANTENNA__3272__B input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3208_ _3208_/A _3219_/B vssd1 vssd1 vccd1 vccd1 _3208_/Y sky130_fd_sc_hd__nand2_1
XFILLER_67_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_32_net107 _3436_/CLK vssd1 vssd1 vccd1 vccd1 _3452_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__1675__B1 _1667_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3139_ _3391_/Q _3053_/X _2945_/A _3475_/Q vssd1 vssd1 vccd1 vccd1 _3139_/X sky130_fd_sc_hd__a22o_1
XFILLER_82_330 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_555 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output101_A _3540_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2542__A _2578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2510_ _3332_/Q _2493_/A _2509_/X _2501_/X vssd1 vssd1 vccd1 vccd1 _3332_/D sky130_fd_sc_hd__o211a_1
X_3490_ _3511_/CLK _3490_/D vssd1 vssd1 vccd1 vccd1 _3490_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2441_ _2568_/A _2441_/B vssd1 vssd1 vccd1 vccd1 _2441_/X sky130_fd_sc_hd__or2_1
XFILLER_5_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2372_ hold2/X vssd1 vssd1 vccd1 vccd1 _2372_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2717__A _2756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2452__A _2574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2708_ _3392_/Q _2692_/A _2707_/X _2699_/X vssd1 vssd1 vccd1 vccd1 _3392_/D sky130_fd_sc_hd__o211a_1
X_2639_ _2997_/A vssd1 vssd1 vccd1 vccd1 _2640_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_99_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2627__A _3183_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_12 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input62_A wbs_dat_i[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1706__A _3262_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_522 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_503 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2990_ _3074_/A vssd1 vssd1 vccd1 vccd1 _2990_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_61_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1941_ _1941_/A _1941_/B vssd1 vssd1 vccd1 vccd1 _2015_/B sky130_fd_sc_hd__nor2_1
X_1872_ _3539_/Q _3538_/Q _1928_/A _1901_/C vssd1 vssd1 vccd1 vccd1 _1873_/D sky130_fd_sc_hd__and4b_1
XANTENNA__3013__C1 _2971_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3542_ _3542_/D _2360_/X vssd1 vssd1 vccd1 vccd1 _3544_/D sky130_fd_sc_hd__dlxtn_1
X_3473_ _3474_/CLK _3473_/D vssd1 vssd1 vccd1 vccd1 _3473_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2424_ _2427_/A _3225_/A vssd1 vssd1 vccd1 vccd1 _2446_/A sky130_fd_sc_hd__nor2b_1
X_2355_ _3294_/Q _3293_/Q vssd1 vssd1 vccd1 vccd1 _2356_/A sky130_fd_sc_hd__and2_1
XFILLER_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2286_ _2286_/A _2286_/B vssd1 vssd1 vccd1 vccd1 _2347_/B sky130_fd_sc_hd__nor2_1
XFILLER_84_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2447__A _3238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_35 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3809_ input1/X vssd1 vssd1 vccd1 vccd1 _3809_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_69_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrlbp_macro_213 vssd1 vssd1 vccd1 vccd1 rlbp_macro_213/HI la_data_out[15] sky130_fd_sc_hd__conb_1
Xrlbp_macro_224 vssd1 vssd1 vccd1 vccd1 rlbp_macro_224/HI la_data_out[26] sky130_fd_sc_hd__conb_1
Xrlbp_macro_202 vssd1 vssd1 vccd1 vccd1 rlbp_macro_202/HI la_data_out[4] sky130_fd_sc_hd__conb_1
Xrlbp_macro_235 vssd1 vssd1 vccd1 vccd1 rlbp_macro_235/HI la_data_out[37] sky130_fd_sc_hd__conb_1
Xrlbp_macro_246 vssd1 vssd1 vccd1 vccd1 rlbp_macro_246/HI la_data_out[48] sky130_fd_sc_hd__conb_1
Xrlbp_macro_257 vssd1 vssd1 vccd1 vccd1 rlbp_macro_257/HI la_data_out[59] sky130_fd_sc_hd__conb_1
XFILLER_0_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrlbp_macro_268 vssd1 vssd1 vccd1 vccd1 rlbp_macro_268/HI la_data_out[70] sky130_fd_sc_hd__conb_1
Xrlbp_macro_279 vssd1 vssd1 vccd1 vccd1 rlbp_macro_279/HI la_data_out[81] sky130_fd_sc_hd__conb_1
XFILLER_87_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3188__A _3188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2820__A _3181_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_6 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2140_ _2161_/A _2159_/B _2161_/B _2139_/Y vssd1 vssd1 vccd1 vccd1 _2155_/B sky130_fd_sc_hd__a31o_1
XFILLER_66_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2071_ _3338_/Q _2071_/B vssd1 vssd1 vccd1 vccd1 _2072_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_clkbuf_leaf_5_net107_A clkbuf_leaf_9_net107/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2973_ _2973_/A _2973_/B vssd1 vssd1 vccd1 vccd1 _2973_/X sky130_fd_sc_hd__or2_1
X_1924_ _1921_/Y _1834_/X _1854_/D _1911_/B _1923_/X vssd1 vssd1 vccd1 vccd1 _1928_/B
+ sky130_fd_sc_hd__a221o_1
X_1855_ _3421_/Q _2105_/B vssd1 vssd1 vccd1 vccd1 _1895_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__2730__A _2769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1786_ _1786_/A _1786_/B vssd1 vssd1 vccd1 vccd1 _1787_/A sky130_fd_sc_hd__and2_1
X_3525_ _3528_/CLK _3525_/D vssd1 vssd1 vccd1 vccd1 _3525_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3456_ _3464_/CLK _3456_/D vssd1 vssd1 vccd1 vccd1 _3456_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3387_ _3387_/CLK _3387_/D vssd1 vssd1 vccd1 vccd1 _3387_/Q sky130_fd_sc_hd__dfxtp_1
X_2407_ _2407_/A _2407_/B vssd1 vssd1 vccd1 vccd1 _2412_/C sky130_fd_sc_hd__and2_1
X_2338_ _2338_/A _2338_/B _2338_/C _2338_/D vssd1 vssd1 vccd1 vccd1 _2352_/B sky130_fd_sc_hd__or4_1
X_2269_ _2269_/A _2269_/B _2269_/C _2269_/D vssd1 vssd1 vccd1 vccd1 _2269_/X sky130_fd_sc_hd__or4_1
XANTENNA__2177__A _3375_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3068__A2 _3053_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_480 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input25_A la_data_in[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3190__B _3195_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1703__B _2294_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1793__A2 _2395_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3310_ _3322_/CLK _3310_/D vssd1 vssd1 vccd1 vccd1 _3310_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3241_ _3241_/A _3243_/B vssd1 vssd1 vccd1 vccd1 _3241_/X sky130_fd_sc_hd__or2_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3172_ _3493_/Q _3159_/X _3170_/X _3171_/X vssd1 vssd1 vccd1 vccd1 _3493_/D sky130_fd_sc_hd__o211a_1
XFILLER_39_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2123_ _3358_/Q _2389_/B vssd1 vssd1 vccd1 vccd1 _2163_/A sky130_fd_sc_hd__xnor2_1
XFILLER_66_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2709__B _2709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2054_ _3347_/Q _2190_/B vssd1 vssd1 vccd1 vccd1 _2054_/X sky130_fd_sc_hd__and2b_1
XFILLER_54_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_480 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1886__A_N _1796_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0_net107 _1749_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0_net107/X sky130_fd_sc_hd__clkbuf_16
XFILLER_10_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2956_ _3467_/Q _2948_/X _2955_/X _2939_/X vssd1 vssd1 vccd1 vccd1 _3467_/D sky130_fd_sc_hd__o211a_1
X_1907_ _1907_/A _1907_/B vssd1 vssd1 vccd1 vccd1 _1908_/B sky130_fd_sc_hd__xor2_1
X_2887_ _3445_/Q _2874_/X _2886_/X _2882_/X vssd1 vssd1 vccd1 vccd1 _3445_/D sky130_fd_sc_hd__o211a_1
X_1838_ _3439_/Q _1838_/B vssd1 vssd1 vccd1 vccd1 _1842_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__2460__A _3183_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1769_ _2145_/A _3448_/Q vssd1 vssd1 vccd1 vccd1 _1772_/A sky130_fd_sc_hd__and2b_1
X_3508_ _3511_/CLK _3508_/D vssd1 vssd1 vccd1 vccd1 _3508_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3289__A2 _3281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3439_ _3440_/CLK _3439_/D vssd1 vssd1 vccd1 vccd1 _3439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3538__RESET_B _3276_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2370__A _2742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput85 _3794_/X vssd1 vssd1 vccd1 vccd1 Pd5_a sky130_fd_sc_hd__buf_2
Xoutput74 _3783_/X vssd1 vssd1 vccd1 vccd1 Pd11_b sky130_fd_sc_hd__buf_2
Xoutput96 _3535_/Q vssd1 vssd1 vccd1 vccd1 Sh sky130_fd_sc_hd__buf_2
XFILLER_95_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1714__A _3491_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3790_ _3790_/A vssd1 vssd1 vccd1 vccd1 _3790_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_31_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2810_ _2830_/B vssd1 vssd1 vccd1 vccd1 _2824_/B sky130_fd_sc_hd__clkbuf_1
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2741_ _2780_/A _2745_/B vssd1 vssd1 vccd1 vccd1 _2741_/X sky130_fd_sc_hd__or2_1
XFILLER_31_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2672_ _2782_/A _2672_/B vssd1 vssd1 vccd1 vccd1 _2672_/X sky130_fd_sc_hd__or2_1
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3224_ _3224_/A vssd1 vssd1 vccd1 vccd1 _3224_/X sky130_fd_sc_hd__dlymetal6s2s_1
.ends

