magic
tech sky130B
magscale 1 2
timestamp 1662149813
<< viali >>
rect 9413 33541 9447 33575
rect 1685 33473 1719 33507
rect 2237 33473 2271 33507
rect 20085 33473 20119 33507
rect 25789 33473 25823 33507
rect 32137 33473 32171 33507
rect 37289 33473 37323 33507
rect 1501 33269 1535 33303
rect 9505 33269 9539 33303
rect 1501 33065 1535 33099
rect 9137 33065 9171 33099
rect 11805 32929 11839 32963
rect 1685 32861 1719 32895
rect 11529 32861 11563 32895
rect 2237 32725 2271 32759
rect 3341 32385 3375 32419
rect 6745 32385 6779 32419
rect 11796 32385 11830 32419
rect 17417 32385 17451 32419
rect 17693 32385 17727 32419
rect 3617 32317 3651 32351
rect 6469 32317 6503 32351
rect 11529 32317 11563 32351
rect 2605 32181 2639 32215
rect 7481 32181 7515 32215
rect 10885 32181 10919 32215
rect 12909 32181 12943 32215
rect 16681 32181 16715 32215
rect 2881 31977 2915 32011
rect 6653 31977 6687 32011
rect 26065 31977 26099 32011
rect 29009 31977 29043 32011
rect 2237 31909 2271 31943
rect 11529 31909 11563 31943
rect 16405 31909 16439 31943
rect 18337 31909 18371 31943
rect 20913 31909 20947 31943
rect 22385 31909 22419 31943
rect 22845 31909 22879 31943
rect 12541 31841 12575 31875
rect 21373 31841 21407 31875
rect 23857 31841 23891 31875
rect 1685 31773 1719 31807
rect 2697 31773 2731 31807
rect 6469 31773 6503 31807
rect 9137 31773 9171 31807
rect 12265 31773 12299 31807
rect 16221 31773 16255 31807
rect 17325 31773 17359 31807
rect 17601 31773 17635 31807
rect 20729 31773 20763 31807
rect 21649 31773 21683 31807
rect 23581 31773 23615 31807
rect 25053 31773 25087 31807
rect 25329 31773 25363 31807
rect 27997 31773 28031 31807
rect 28273 31773 28307 31807
rect 1501 31637 1535 31671
rect 8953 31637 8987 31671
rect 2697 31433 2731 31467
rect 6745 31433 6779 31467
rect 8033 31433 8067 31467
rect 11897 31433 11931 31467
rect 15209 31433 15243 31467
rect 16865 31433 16899 31467
rect 20453 31433 20487 31467
rect 22017 31433 22051 31467
rect 29285 31433 29319 31467
rect 2881 31297 2915 31331
rect 6561 31297 6595 31331
rect 8769 31297 8803 31331
rect 9045 31297 9079 31331
rect 11713 31297 11747 31331
rect 15025 31297 15059 31331
rect 15853 31297 15887 31331
rect 16037 31297 16071 31331
rect 16681 31297 16715 31331
rect 20269 31297 20303 31331
rect 21833 31297 21867 31331
rect 28549 31297 28583 31331
rect 3065 31229 3099 31263
rect 3525 31229 3559 31263
rect 6377 31229 6411 31263
rect 14841 31229 14875 31263
rect 15669 31229 15703 31263
rect 19625 31229 19659 31263
rect 20085 31229 20119 31263
rect 28273 31229 28307 31263
rect 4997 30889 5031 30923
rect 8953 30889 8987 30923
rect 15577 30889 15611 30923
rect 21373 30889 21407 30923
rect 24777 30889 24811 30923
rect 25421 30889 25455 30923
rect 28641 30889 28675 30923
rect 29561 30889 29595 30923
rect 3985 30753 4019 30787
rect 1685 30685 1719 30719
rect 4261 30685 4295 30719
rect 9137 30685 9171 30719
rect 9321 30685 9355 30719
rect 21005 30685 21039 30719
rect 21189 30685 21223 30719
rect 24593 30685 24627 30719
rect 25237 30685 25271 30719
rect 28825 30685 28859 30719
rect 29745 30685 29779 30719
rect 21833 30617 21867 30651
rect 1501 30549 1535 30583
rect 9873 30549 9907 30583
rect 4261 30345 4295 30379
rect 11897 30345 11931 30379
rect 3433 30209 3467 30243
rect 3617 30209 3651 30243
rect 4077 30209 4111 30243
rect 11713 30209 11747 30243
rect 24777 30209 24811 30243
rect 3249 30141 3283 30175
rect 11529 30141 11563 30175
rect 24501 30141 24535 30175
rect 12449 30005 12483 30039
rect 25513 30005 25547 30039
rect 2605 29801 2639 29835
rect 11805 29801 11839 29835
rect 25145 29801 25179 29835
rect 28733 29801 28767 29835
rect 24777 29665 24811 29699
rect 2789 29597 2823 29631
rect 12541 29597 12575 29631
rect 12817 29597 12851 29631
rect 24961 29597 24995 29631
rect 28457 29597 28491 29631
rect 28549 29597 28583 29631
rect 25605 29529 25639 29563
rect 29561 29529 29595 29563
rect 3893 29461 3927 29495
rect 12817 29257 12851 29291
rect 24777 29257 24811 29291
rect 29101 29257 29135 29291
rect 31401 29257 31435 29291
rect 32689 29257 32723 29291
rect 1685 29121 1719 29155
rect 11805 29121 11839 29155
rect 13001 29121 13035 29155
rect 15853 29121 15887 29155
rect 17509 29121 17543 29155
rect 24961 29121 24995 29155
rect 28917 29121 28951 29155
rect 31309 29121 31343 29155
rect 32597 29121 32631 29155
rect 11529 29053 11563 29087
rect 15669 29053 15703 29087
rect 17233 29053 17267 29087
rect 28733 29053 28767 29087
rect 1501 28985 1535 29019
rect 2145 28985 2179 29019
rect 2973 28985 3007 29019
rect 16037 28985 16071 29019
rect 18245 28985 18279 29019
rect 13461 28917 13495 28951
rect 12541 28713 12575 28747
rect 16865 28713 16899 28747
rect 34805 28713 34839 28747
rect 20085 28645 20119 28679
rect 14381 28577 14415 28611
rect 21005 28577 21039 28611
rect 9137 28509 9171 28543
rect 12265 28509 12299 28543
rect 12357 28509 12391 28543
rect 13185 28509 13219 28543
rect 14105 28509 14139 28543
rect 16681 28509 16715 28543
rect 20269 28509 20303 28543
rect 20729 28509 20763 28543
rect 22017 28509 22051 28543
rect 31585 28441 31619 28475
rect 8953 28373 8987 28407
rect 13001 28373 13035 28407
rect 15485 28373 15519 28407
rect 32321 28373 32355 28407
rect 24961 28169 24995 28203
rect 29193 28169 29227 28203
rect 19073 28101 19107 28135
rect 19625 28101 19659 28135
rect 1685 28033 1719 28067
rect 8401 28033 8435 28067
rect 21005 28033 21039 28067
rect 21281 28033 21315 28067
rect 24777 28033 24811 28067
rect 28181 28033 28215 28067
rect 28457 28033 28491 28067
rect 34345 28033 34379 28067
rect 35173 28033 35207 28067
rect 35357 28033 35391 28067
rect 35817 28033 35851 28067
rect 8125 27965 8159 27999
rect 24593 27965 24627 27999
rect 34161 27965 34195 27999
rect 34989 27965 35023 27999
rect 12909 27897 12943 27931
rect 20269 27897 20303 27931
rect 1501 27829 1535 27863
rect 2237 27829 2271 27863
rect 9137 27829 9171 27863
rect 13461 27829 13495 27863
rect 19717 27829 19751 27863
rect 24133 27829 24167 27863
rect 34529 27829 34563 27863
rect 36001 27829 36035 27863
rect 8953 27625 8987 27659
rect 21005 27625 21039 27659
rect 6101 27557 6135 27591
rect 24777 27557 24811 27591
rect 31677 27557 31711 27591
rect 2697 27421 2731 27455
rect 5089 27421 5123 27455
rect 5365 27421 5399 27455
rect 6745 27421 6779 27455
rect 6929 27421 6963 27455
rect 9137 27421 9171 27455
rect 9321 27421 9355 27455
rect 19993 27421 20027 27455
rect 20177 27421 20211 27455
rect 20361 27421 20395 27455
rect 20821 27421 20855 27455
rect 28549 27421 28583 27455
rect 28641 27421 28675 27455
rect 34989 27421 35023 27455
rect 35633 27421 35667 27455
rect 35909 27421 35943 27455
rect 36737 27421 36771 27455
rect 24961 27353 24995 27387
rect 2881 27285 2915 27319
rect 6561 27285 6595 27319
rect 9873 27285 9907 27319
rect 19441 27285 19475 27319
rect 28825 27285 28859 27319
rect 35173 27285 35207 27319
rect 2513 27081 2547 27115
rect 5549 27081 5583 27115
rect 24133 27081 24167 27115
rect 28549 27081 28583 27115
rect 3249 26945 3283 26979
rect 3525 26945 3559 26979
rect 5733 26945 5767 26979
rect 7849 26945 7883 26979
rect 23949 26945 23983 26979
rect 28733 26945 28767 26979
rect 31309 26945 31343 26979
rect 31401 26945 31435 26979
rect 32965 26945 32999 26979
rect 35909 26945 35943 26979
rect 36737 26945 36771 26979
rect 33241 26877 33275 26911
rect 35633 26877 35667 26911
rect 7665 26741 7699 26775
rect 15485 26741 15519 26775
rect 20545 26741 20579 26775
rect 31585 26741 31619 26775
rect 32219 26741 32253 26775
rect 2881 26537 2915 26571
rect 8401 26537 8435 26571
rect 19257 26537 19291 26571
rect 31861 26537 31895 26571
rect 2237 26469 2271 26503
rect 7389 26401 7423 26435
rect 14933 26401 14967 26435
rect 1685 26333 1719 26367
rect 2421 26333 2455 26367
rect 3065 26333 3099 26367
rect 3157 26333 3191 26367
rect 3801 26333 3835 26367
rect 7665 26333 7699 26367
rect 12357 26333 12391 26367
rect 15117 26333 15151 26367
rect 15761 26333 15795 26367
rect 16037 26333 16071 26367
rect 19441 26333 19475 26367
rect 24869 26333 24903 26367
rect 31677 26333 31711 26367
rect 19625 26265 19659 26299
rect 1501 26197 1535 26231
rect 12173 26197 12207 26231
rect 15301 26197 15335 26231
rect 16773 26197 16807 26231
rect 25053 26197 25087 26231
rect 7757 25993 7791 26027
rect 15945 25993 15979 26027
rect 25789 25993 25823 26027
rect 7573 25857 7607 25891
rect 11989 25857 12023 25891
rect 15761 25857 15795 25891
rect 25053 25857 25087 25891
rect 25973 25857 26007 25891
rect 28457 25857 28491 25891
rect 7389 25789 7423 25823
rect 11713 25789 11747 25823
rect 25329 25789 25363 25823
rect 26157 25789 26191 25823
rect 27077 25789 27111 25823
rect 2605 25653 2639 25687
rect 12725 25653 12759 25687
rect 24317 25653 24351 25687
rect 28273 25653 28307 25687
rect 12265 25449 12299 25483
rect 24409 25449 24443 25483
rect 12633 25313 12667 25347
rect 15577 25313 15611 25347
rect 21833 25313 21867 25347
rect 1685 25245 1719 25279
rect 12449 25245 12483 25279
rect 15853 25245 15887 25279
rect 20821 25245 20855 25279
rect 21005 25245 21039 25279
rect 22109 25245 22143 25279
rect 24593 25245 24627 25279
rect 27537 25245 27571 25279
rect 27813 25245 27847 25279
rect 1501 25109 1535 25143
rect 2237 25109 2271 25143
rect 16589 25109 16623 25143
rect 20269 25109 20303 25143
rect 21189 25109 21223 25143
rect 22845 25109 22879 25143
rect 28549 25109 28583 25143
rect 15945 24905 15979 24939
rect 28365 24905 28399 24939
rect 12725 24769 12759 24803
rect 13461 24769 13495 24803
rect 14933 24769 14967 24803
rect 15117 24769 15151 24803
rect 15301 24769 15335 24803
rect 15761 24769 15795 24803
rect 19993 24769 20027 24803
rect 21833 24769 21867 24803
rect 28549 24769 28583 24803
rect 32965 24769 32999 24803
rect 33609 24769 33643 24803
rect 28733 24701 28767 24735
rect 20177 24633 20211 24667
rect 12817 24565 12851 24599
rect 14473 24565 14507 24599
rect 22017 24565 22051 24599
rect 33149 24565 33183 24599
rect 33793 24565 33827 24599
rect 28457 24225 28491 24259
rect 3065 24157 3099 24191
rect 3801 24157 3835 24191
rect 3985 24157 4019 24191
rect 4169 24157 4203 24191
rect 4629 24157 4663 24191
rect 8953 24157 8987 24191
rect 9229 24157 9263 24191
rect 19441 24157 19475 24191
rect 19901 24157 19935 24191
rect 20085 24157 20119 24191
rect 20269 24157 20303 24191
rect 20913 24157 20947 24191
rect 28641 24157 28675 24191
rect 32873 24157 32907 24191
rect 33149 24157 33183 24191
rect 33977 24157 34011 24191
rect 31125 24089 31159 24123
rect 31769 24089 31803 24123
rect 3249 24021 3283 24055
rect 20729 24021 20763 24055
rect 28825 24021 28859 24055
rect 31217 24021 31251 24055
rect 8033 23817 8067 23851
rect 8493 23817 8527 23851
rect 28733 23817 28767 23851
rect 29193 23817 29227 23851
rect 32965 23817 32999 23851
rect 13461 23749 13495 23783
rect 1685 23681 1719 23715
rect 3617 23681 3651 23715
rect 3893 23681 3927 23715
rect 7849 23681 7883 23715
rect 9229 23681 9263 23715
rect 13277 23681 13311 23715
rect 16865 23681 16899 23715
rect 20637 23681 20671 23715
rect 20913 23681 20947 23715
rect 27997 23681 28031 23715
rect 29377 23681 29411 23715
rect 31309 23681 31343 23715
rect 32781 23681 32815 23715
rect 34805 23681 34839 23715
rect 35633 23681 35667 23715
rect 35909 23681 35943 23715
rect 36737 23681 36771 23715
rect 9505 23613 9539 23647
rect 27721 23613 27755 23647
rect 31585 23613 31619 23647
rect 32597 23613 32631 23647
rect 34161 23613 34195 23647
rect 34621 23613 34655 23647
rect 30297 23545 30331 23579
rect 1501 23477 1535 23511
rect 2881 23477 2915 23511
rect 9965 23477 9999 23511
rect 13921 23477 13955 23511
rect 16681 23477 16715 23511
rect 19901 23477 19935 23511
rect 34989 23477 35023 23511
rect 9873 23273 9907 23307
rect 15393 23273 15427 23307
rect 35725 23273 35759 23307
rect 5549 23137 5583 23171
rect 31217 23137 31251 23171
rect 5733 23069 5767 23103
rect 9045 23069 9079 23103
rect 9229 23069 9263 23103
rect 9413 23069 9447 23103
rect 10057 23069 10091 23103
rect 15577 23069 15611 23103
rect 16037 23069 16071 23103
rect 16313 23069 16347 23103
rect 30941 23069 30975 23103
rect 35541 23069 35575 23103
rect 5917 22933 5951 22967
rect 17049 22933 17083 22967
rect 3893 22729 3927 22763
rect 9965 22729 9999 22763
rect 16681 22729 16715 22763
rect 3157 22593 3191 22627
rect 3341 22593 3375 22627
rect 7021 22593 7055 22627
rect 10149 22593 10183 22627
rect 12633 22593 12667 22627
rect 12817 22593 12851 22627
rect 13461 22593 13495 22627
rect 16865 22593 16899 22627
rect 17049 22593 17083 22627
rect 17509 22593 17543 22627
rect 25697 22593 25731 22627
rect 7205 22525 7239 22559
rect 12449 22525 12483 22559
rect 1409 22389 1443 22423
rect 2973 22389 3007 22423
rect 6837 22389 6871 22423
rect 13277 22389 13311 22423
rect 25881 22389 25915 22423
rect 10793 22185 10827 22219
rect 11805 22185 11839 22219
rect 13277 22049 13311 22083
rect 14749 22049 14783 22083
rect 24409 22049 24443 22083
rect 5825 21981 5859 22015
rect 6929 21981 6963 22015
rect 11161 21981 11195 22015
rect 11621 21981 11655 22015
rect 13001 21981 13035 22015
rect 15025 21981 15059 22015
rect 23673 21981 23707 22015
rect 24685 21981 24719 22015
rect 25973 21981 26007 22015
rect 26249 21981 26283 22015
rect 27077 21981 27111 22015
rect 10977 21913 11011 21947
rect 6009 21845 6043 21879
rect 7113 21845 7147 21879
rect 12265 21845 12299 21879
rect 23857 21845 23891 21879
rect 25421 21845 25455 21879
rect 18981 21641 19015 21675
rect 22385 21641 22419 21675
rect 23673 21641 23707 21675
rect 25329 21641 25363 21675
rect 3065 21505 3099 21539
rect 18797 21505 18831 21539
rect 19901 21505 19935 21539
rect 22201 21505 22235 21539
rect 23489 21505 23523 21539
rect 25145 21505 25179 21539
rect 34069 21505 34103 21539
rect 34529 21505 34563 21539
rect 34713 21505 34747 21539
rect 23305 21437 23339 21471
rect 24961 21437 24995 21471
rect 2881 21301 2915 21335
rect 20085 21301 20119 21335
rect 34897 21301 34931 21335
rect 19993 20961 20027 20995
rect 1685 20893 1719 20927
rect 2973 20893 3007 20927
rect 3249 20893 3283 20927
rect 6009 20893 6043 20927
rect 6285 20893 6319 20927
rect 6745 20893 6779 20927
rect 7021 20893 7055 20927
rect 20269 20893 20303 20927
rect 29745 20893 29779 20927
rect 30573 20893 30607 20927
rect 36001 20893 36035 20927
rect 1501 20757 1535 20791
rect 2237 20757 2271 20791
rect 5273 20757 5307 20791
rect 7757 20757 7791 20791
rect 19257 20757 19291 20791
rect 21005 20757 21039 20791
rect 29929 20757 29963 20791
rect 30389 20757 30423 20791
rect 36185 20757 36219 20791
rect 1777 20553 1811 20587
rect 7757 20553 7791 20587
rect 19809 20553 19843 20587
rect 30205 20553 30239 20587
rect 8309 20485 8343 20519
rect 18337 20485 18371 20519
rect 16957 20417 16991 20451
rect 19625 20417 19659 20451
rect 29561 20417 29595 20451
rect 30389 20417 30423 20451
rect 30573 20417 30607 20451
rect 33149 20417 33183 20451
rect 33333 20417 33367 20451
rect 34253 20417 34287 20451
rect 34437 20417 34471 20451
rect 35081 20417 35115 20451
rect 17233 20349 17267 20383
rect 19441 20349 19475 20383
rect 29377 20349 29411 20383
rect 29745 20349 29779 20383
rect 34069 20349 34103 20383
rect 9597 20213 9631 20247
rect 33517 20213 33551 20247
rect 35265 20213 35299 20247
rect 6653 20009 6687 20043
rect 14841 20009 14875 20043
rect 16865 20009 16899 20043
rect 17325 19941 17359 19975
rect 15117 19873 15151 19907
rect 15853 19873 15887 19907
rect 20637 19873 20671 19907
rect 21097 19873 21131 19907
rect 1685 19805 1719 19839
rect 6469 19805 6503 19839
rect 15209 19805 15243 19839
rect 16129 19805 16163 19839
rect 17509 19805 17543 19839
rect 21281 19805 21315 19839
rect 29653 19805 29687 19839
rect 29929 19805 29963 19839
rect 33885 19805 33919 19839
rect 35725 19805 35759 19839
rect 36001 19805 36035 19839
rect 2237 19737 2271 19771
rect 14749 19737 14783 19771
rect 1501 19669 1535 19703
rect 15393 19669 15427 19703
rect 21465 19669 21499 19703
rect 30665 19669 30699 19703
rect 34069 19669 34103 19703
rect 36737 19669 36771 19703
rect 17049 19465 17083 19499
rect 25513 19465 25547 19499
rect 30665 19465 30699 19499
rect 33977 19465 34011 19499
rect 10701 19397 10735 19431
rect 3433 19329 3467 19363
rect 7113 19329 7147 19363
rect 10057 19329 10091 19363
rect 10149 19329 10183 19363
rect 16865 19329 16899 19363
rect 22017 19329 22051 19363
rect 25329 19329 25363 19363
rect 25973 19329 26007 19363
rect 29653 19329 29687 19363
rect 29929 19329 29963 19363
rect 34713 19329 34747 19363
rect 34989 19329 35023 19363
rect 3249 19261 3283 19295
rect 4077 19261 4111 19295
rect 16681 19261 16715 19295
rect 26157 19193 26191 19227
rect 3617 19125 3651 19159
rect 6929 19125 6963 19159
rect 21833 19125 21867 19159
rect 7389 18921 7423 18955
rect 10057 18921 10091 18955
rect 20913 18921 20947 18955
rect 26249 18921 26283 18955
rect 10609 18785 10643 18819
rect 24409 18785 24443 18819
rect 3985 18717 4019 18751
rect 6377 18717 6411 18751
rect 6653 18717 6687 18751
rect 9873 18717 9907 18751
rect 21649 18717 21683 18751
rect 21925 18717 21959 18751
rect 24593 18717 24627 18751
rect 25237 18717 25271 18751
rect 25513 18717 25547 18751
rect 36645 18717 36679 18751
rect 36921 18717 36955 18751
rect 10885 18649 10919 18683
rect 3801 18581 3835 18615
rect 12357 18581 12391 18615
rect 24777 18581 24811 18615
rect 37657 18581 37691 18615
rect 6929 18377 6963 18411
rect 13001 18377 13035 18411
rect 25421 18377 25455 18411
rect 7849 18309 7883 18343
rect 14105 18309 14139 18343
rect 1685 18241 1719 18275
rect 3617 18241 3651 18275
rect 3893 18241 3927 18275
rect 7113 18241 7147 18275
rect 13645 18241 13679 18275
rect 14381 18241 14415 18275
rect 14565 18241 14599 18275
rect 25237 18241 25271 18275
rect 7297 18173 7331 18207
rect 9597 18173 9631 18207
rect 14197 18173 14231 18207
rect 1501 18037 1535 18071
rect 2145 18037 2179 18071
rect 2881 18037 2915 18071
rect 14289 18037 14323 18071
rect 9321 17833 9355 17867
rect 14749 17833 14783 17867
rect 4629 17697 4663 17731
rect 15393 17697 15427 17731
rect 4905 17629 4939 17663
rect 9137 17629 9171 17663
rect 14749 17629 14783 17663
rect 14933 17629 14967 17663
rect 24685 17629 24719 17663
rect 24961 17629 24995 17663
rect 26985 17629 27019 17663
rect 27077 17629 27111 17663
rect 27261 17629 27295 17663
rect 28089 17629 28123 17663
rect 8953 17561 8987 17595
rect 7481 17493 7515 17527
rect 28273 17493 28307 17527
rect 17601 17289 17635 17323
rect 17785 17289 17819 17323
rect 18981 17289 19015 17323
rect 22477 17289 22511 17323
rect 27445 17289 27479 17323
rect 18613 17221 18647 17255
rect 18829 17221 18863 17255
rect 22109 17221 22143 17255
rect 22309 17221 22343 17255
rect 1685 17153 1719 17187
rect 2237 17153 2271 17187
rect 28825 17153 28859 17187
rect 29101 17153 29135 17187
rect 32597 17153 32631 17187
rect 33057 17153 33091 17187
rect 33241 17153 33275 17187
rect 35817 17153 35851 17187
rect 18153 17017 18187 17051
rect 29837 17017 29871 17051
rect 1501 16949 1535 16983
rect 17785 16949 17819 16983
rect 18797 16949 18831 16983
rect 22293 16949 22327 16983
rect 33425 16949 33459 16983
rect 36001 16949 36035 16983
rect 4721 16745 4755 16779
rect 11897 16745 11931 16779
rect 21649 16745 21683 16779
rect 35081 16745 35115 16779
rect 2237 16677 2271 16711
rect 6193 16677 6227 16711
rect 16129 16677 16163 16711
rect 36737 16677 36771 16711
rect 3249 16609 3283 16643
rect 9781 16609 9815 16643
rect 12081 16609 12115 16643
rect 19809 16609 19843 16643
rect 20085 16609 20119 16643
rect 21097 16609 21131 16643
rect 22845 16609 22879 16643
rect 22937 16609 22971 16643
rect 2973 16541 3007 16575
rect 3985 16541 4019 16575
rect 4169 16541 4203 16575
rect 7021 16541 7055 16575
rect 10057 16541 10091 16575
rect 12173 16541 12207 16575
rect 22661 16541 22695 16575
rect 32505 16541 32539 16575
rect 33977 16541 34011 16575
rect 34713 16541 34747 16575
rect 34897 16541 34931 16575
rect 35725 16541 35759 16575
rect 36001 16541 36035 16575
rect 6377 16473 6411 16507
rect 11897 16473 11931 16507
rect 15853 16473 15887 16507
rect 21281 16473 21315 16507
rect 21373 16473 21407 16507
rect 23029 16473 23063 16507
rect 3801 16405 3835 16439
rect 7113 16405 7147 16439
rect 11345 16405 11379 16439
rect 12357 16405 12391 16439
rect 16313 16405 16347 16439
rect 21465 16405 21499 16439
rect 22753 16405 22787 16439
rect 32689 16405 32723 16439
rect 34161 16405 34195 16439
rect 2973 16201 3007 16235
rect 10517 16201 10551 16235
rect 11529 16201 11563 16235
rect 19809 16201 19843 16235
rect 25881 16201 25915 16235
rect 35909 16201 35943 16235
rect 7849 16133 7883 16167
rect 12265 16133 12299 16167
rect 2789 16065 2823 16099
rect 10241 16065 10275 16099
rect 19625 16065 19659 16099
rect 26065 16065 26099 16099
rect 26157 16065 26191 16099
rect 26341 16065 26375 16099
rect 26433 16065 26467 16099
rect 29745 16065 29779 16099
rect 35725 16065 35759 16099
rect 10149 15997 10183 16031
rect 10333 15997 10367 16031
rect 11713 15997 11747 16031
rect 11805 15997 11839 16031
rect 29561 15997 29595 16031
rect 12265 15929 12299 15963
rect 29009 15929 29043 15963
rect 34529 15929 34563 15963
rect 9137 15861 9171 15895
rect 29929 15861 29963 15895
rect 9873 15657 9907 15691
rect 24501 15657 24535 15691
rect 30757 15657 30791 15691
rect 37473 15657 37507 15691
rect 9137 15589 9171 15623
rect 11437 15589 11471 15623
rect 14105 15589 14139 15623
rect 2237 15521 2271 15555
rect 29745 15521 29779 15555
rect 36461 15521 36495 15555
rect 1685 15453 1719 15487
rect 11621 15453 11655 15487
rect 14381 15453 14415 15487
rect 14565 15453 14599 15487
rect 14841 15453 14875 15487
rect 15117 15453 15151 15487
rect 30021 15453 30055 15487
rect 36737 15453 36771 15487
rect 9137 15385 9171 15419
rect 9597 15385 9631 15419
rect 24685 15385 24719 15419
rect 24869 15385 24903 15419
rect 1501 15317 1535 15351
rect 9689 15317 9723 15351
rect 18797 15113 18831 15147
rect 26249 15113 26283 15147
rect 30021 15113 30055 15147
rect 35541 15113 35575 15147
rect 25881 15045 25915 15079
rect 10425 14977 10459 15011
rect 16037 14977 16071 15011
rect 17785 14977 17819 15011
rect 18981 14977 19015 15011
rect 25789 14977 25823 15011
rect 26065 14977 26099 15011
rect 30205 14977 30239 15011
rect 32873 14977 32907 15011
rect 34805 14977 34839 15011
rect 10149 14909 10183 14943
rect 15761 14909 15795 14943
rect 17509 14909 17543 14943
rect 26985 14909 27019 14943
rect 27261 14909 27295 14943
rect 34529 14909 34563 14943
rect 33057 14841 33091 14875
rect 8861 14773 8895 14807
rect 26985 14569 27019 14603
rect 31309 14569 31343 14603
rect 31493 14569 31527 14603
rect 33701 14569 33735 14603
rect 9965 14433 9999 14467
rect 15209 14433 15243 14467
rect 16497 14433 16531 14467
rect 17877 14433 17911 14467
rect 21833 14433 21867 14467
rect 22318 14433 22352 14467
rect 31217 14433 31251 14467
rect 1685 14365 1719 14399
rect 2145 14365 2179 14399
rect 5457 14365 5491 14399
rect 9689 14365 9723 14399
rect 15485 14365 15519 14399
rect 16773 14365 16807 14399
rect 18153 14365 18187 14399
rect 22109 14365 22143 14399
rect 26801 14365 26835 14399
rect 31125 14365 31159 14399
rect 31953 14365 31987 14399
rect 33517 14365 33551 14399
rect 5733 14297 5767 14331
rect 1501 14229 1535 14263
rect 7205 14229 7239 14263
rect 22201 14229 22235 14263
rect 22477 14229 22511 14263
rect 32137 14229 32171 14263
rect 7757 14025 7791 14059
rect 8401 14025 8435 14059
rect 22201 14025 22235 14059
rect 22477 14025 22511 14059
rect 23489 14025 23523 14059
rect 32505 14025 32539 14059
rect 22318 13957 22352 13991
rect 23305 13957 23339 13991
rect 26985 13957 27019 13991
rect 7849 13889 7883 13923
rect 17601 13889 17635 13923
rect 22109 13889 22143 13923
rect 27169 13889 27203 13923
rect 27261 13889 27295 13923
rect 32321 13889 32355 13923
rect 17877 13821 17911 13855
rect 21833 13821 21867 13855
rect 22937 13821 22971 13855
rect 26341 13821 26375 13855
rect 31493 13821 31527 13855
rect 32137 13821 32171 13855
rect 23305 13685 23339 13719
rect 27261 13685 27295 13719
rect 27445 13685 27479 13719
rect 6377 13481 6411 13515
rect 11529 13481 11563 13515
rect 21097 13481 21131 13515
rect 21281 13481 21315 13515
rect 7205 13413 7239 13447
rect 12357 13413 12391 13447
rect 25053 13413 25087 13447
rect 17785 13345 17819 13379
rect 19257 13345 19291 13379
rect 6561 13277 6595 13311
rect 7389 13277 7423 13311
rect 8033 13277 8067 13311
rect 9321 13277 9355 13311
rect 12173 13277 12207 13311
rect 16865 13277 16899 13311
rect 17049 13277 17083 13311
rect 17509 13277 17543 13311
rect 19533 13277 19567 13311
rect 22017 13277 22051 13311
rect 22201 13277 22235 13311
rect 22477 13277 22511 13311
rect 16957 13209 16991 13243
rect 20913 13209 20947 13243
rect 24869 13209 24903 13243
rect 7849 13141 7883 13175
rect 9137 13141 9171 13175
rect 21113 13141 21147 13175
rect 22661 13141 22695 13175
rect 3525 12937 3559 12971
rect 21925 12937 21959 12971
rect 27185 12937 27219 12971
rect 30665 12937 30699 12971
rect 31585 12937 31619 12971
rect 33517 12937 33551 12971
rect 2237 12869 2271 12903
rect 19257 12869 19291 12903
rect 26985 12869 27019 12903
rect 31217 12869 31251 12903
rect 31422 12869 31456 12903
rect 32137 12869 32171 12903
rect 32337 12869 32371 12903
rect 1685 12801 1719 12835
rect 3433 12801 3467 12835
rect 3709 12801 3743 12835
rect 14197 12801 14231 12835
rect 18613 12801 18647 12835
rect 19349 12801 19383 12835
rect 21833 12801 21867 12835
rect 22017 12801 22051 12835
rect 23765 12801 23799 12835
rect 33333 12801 33367 12835
rect 34621 12801 34655 12835
rect 35357 12801 35391 12835
rect 35633 12801 35667 12835
rect 14013 12733 14047 12767
rect 14105 12733 14139 12767
rect 14289 12733 14323 12767
rect 18429 12733 18463 12767
rect 23949 12665 23983 12699
rect 32505 12665 32539 12699
rect 1501 12597 1535 12631
rect 2973 12597 3007 12631
rect 3709 12597 3743 12631
rect 4261 12597 4295 12631
rect 13277 12597 13311 12631
rect 13829 12597 13863 12631
rect 14841 12597 14875 12631
rect 17969 12597 18003 12631
rect 20177 12597 20211 12631
rect 26341 12597 26375 12631
rect 27169 12597 27203 12631
rect 27353 12597 27387 12631
rect 31401 12597 31435 12631
rect 32321 12597 32355 12631
rect 34805 12597 34839 12631
rect 36369 12597 36403 12631
rect 5595 12393 5629 12427
rect 31953 12393 31987 12427
rect 15209 12325 15243 12359
rect 3801 12257 3835 12291
rect 13553 12257 13587 12291
rect 14381 12257 14415 12291
rect 14749 12257 14783 12291
rect 35817 12257 35851 12291
rect 3065 12189 3099 12223
rect 4169 12189 4203 12223
rect 9413 12189 9447 12223
rect 9873 12189 9907 12223
rect 13277 12189 13311 12223
rect 14289 12189 14323 12223
rect 25053 12189 25087 12223
rect 27353 12189 27387 12223
rect 36093 12189 36127 12223
rect 2421 12053 2455 12087
rect 3157 12053 3191 12087
rect 9229 12053 9263 12087
rect 14105 12053 14139 12087
rect 14565 12053 14599 12087
rect 14657 12053 14691 12087
rect 25237 12053 25271 12087
rect 27169 12053 27203 12087
rect 36829 12053 36863 12087
rect 3801 11849 3835 11883
rect 6469 11849 6503 11883
rect 8585 11849 8619 11883
rect 12725 11849 12759 11883
rect 14473 11849 14507 11883
rect 14565 11849 14599 11883
rect 13185 11781 13219 11815
rect 1685 11713 1719 11747
rect 2881 11713 2915 11747
rect 3433 11713 3467 11747
rect 3617 11713 3651 11747
rect 6561 11713 6595 11747
rect 10793 11713 10827 11747
rect 14197 11713 14231 11747
rect 14657 11713 14691 11747
rect 15117 11713 15151 11747
rect 18061 11713 18095 11747
rect 18245 11713 18279 11747
rect 26985 11713 27019 11747
rect 27261 11713 27295 11747
rect 28457 11713 28491 11747
rect 28733 11713 28767 11747
rect 3341 11645 3375 11679
rect 10517 11645 10551 11679
rect 12909 11577 12943 11611
rect 14197 11577 14231 11611
rect 1501 11509 1535 11543
rect 2237 11509 2271 11543
rect 9045 11509 9079 11543
rect 14289 11509 14323 11543
rect 18061 11509 18095 11543
rect 27997 11509 28031 11543
rect 29469 11509 29503 11543
rect 10057 11305 10091 11339
rect 13553 11305 13587 11339
rect 16497 11305 16531 11339
rect 24593 11305 24627 11339
rect 26985 11305 27019 11339
rect 31677 11305 31711 11339
rect 32505 11305 32539 11339
rect 14749 11237 14783 11271
rect 24777 11237 24811 11271
rect 32689 11237 32723 11271
rect 31033 11169 31067 11203
rect 10149 11101 10183 11135
rect 14565 11101 14599 11135
rect 16497 11101 16531 11135
rect 16773 11101 16807 11135
rect 26801 11101 26835 11135
rect 17325 11033 17359 11067
rect 24409 11033 24443 11067
rect 24625 11033 24659 11067
rect 31493 11033 31527 11067
rect 31693 11033 31727 11067
rect 32321 11033 32355 11067
rect 32521 11033 32555 11067
rect 16681 10965 16715 10999
rect 31861 10965 31895 10999
rect 18061 10761 18095 10795
rect 22937 10761 22971 10795
rect 32137 10761 32171 10795
rect 33241 10761 33275 10795
rect 35817 10761 35851 10795
rect 7097 10693 7131 10727
rect 7297 10693 7331 10727
rect 18245 10693 18279 10727
rect 18429 10693 18463 10727
rect 22293 10693 22327 10727
rect 22477 10693 22511 10727
rect 18153 10625 18187 10659
rect 33057 10625 33091 10659
rect 33701 10625 33735 10659
rect 34805 10625 34839 10659
rect 35081 10625 35115 10659
rect 6929 10421 6963 10455
rect 7113 10421 7147 10455
rect 17877 10421 17911 10455
rect 18981 10421 19015 10455
rect 33885 10421 33919 10455
rect 36553 10217 36587 10251
rect 16037 10081 16071 10115
rect 16313 10081 16347 10115
rect 35541 10081 35575 10115
rect 1685 10013 1719 10047
rect 4905 10013 4939 10047
rect 27445 10013 27479 10047
rect 35817 10013 35851 10047
rect 2237 9945 2271 9979
rect 1501 9877 1535 9911
rect 4721 9877 4755 9911
rect 27261 9877 27295 9911
rect 7205 9605 7239 9639
rect 22109 9537 22143 9571
rect 22937 9537 22971 9571
rect 24409 9537 24443 9571
rect 21833 9469 21867 9503
rect 6929 9401 6963 9435
rect 3249 9333 3283 9367
rect 6745 9333 6779 9367
rect 24593 9333 24627 9367
rect 31033 9333 31067 9367
rect 2881 9129 2915 9163
rect 22017 9129 22051 9163
rect 22661 9129 22695 9163
rect 22845 9129 22879 9163
rect 31401 9129 31435 9163
rect 32045 9061 32079 9095
rect 2237 8993 2271 9027
rect 21097 8993 21131 9027
rect 23305 8993 23339 9027
rect 27445 8993 27479 9027
rect 1685 8925 1719 8959
rect 6653 8925 6687 8959
rect 20913 8925 20947 8959
rect 22017 8925 22051 8959
rect 27169 8925 27203 8959
rect 30573 8925 30607 8959
rect 31217 8925 31251 8959
rect 2697 8857 2731 8891
rect 3893 8857 3927 8891
rect 22477 8857 22511 8891
rect 22693 8857 22727 8891
rect 1501 8789 1535 8823
rect 2897 8789 2931 8823
rect 3065 8789 3099 8823
rect 6561 8789 6595 8823
rect 7389 8789 7423 8823
rect 26433 8789 26467 8823
rect 30757 8789 30791 8823
rect 4997 8585 5031 8619
rect 7005 8585 7039 8619
rect 8099 8585 8133 8619
rect 8861 8585 8895 8619
rect 9413 8585 9447 8619
rect 19073 8585 19107 8619
rect 19809 8585 19843 8619
rect 30481 8585 30515 8619
rect 31401 8585 31435 8619
rect 2881 8517 2915 8551
rect 3097 8517 3131 8551
rect 7205 8517 7239 8551
rect 8309 8517 8343 8551
rect 20637 8517 20671 8551
rect 20821 8517 20855 8551
rect 23581 8517 23615 8551
rect 23797 8517 23831 8551
rect 30021 8517 30055 8551
rect 31033 8517 31067 8551
rect 31233 8517 31267 8551
rect 32137 8517 32171 8551
rect 32337 8517 32371 8551
rect 3709 8449 3743 8483
rect 13185 8449 13219 8483
rect 17785 8449 17819 8483
rect 19257 8449 19291 8483
rect 22293 8449 22327 8483
rect 26985 8449 27019 8483
rect 27905 8449 27939 8483
rect 17509 8381 17543 8415
rect 22017 8381 22051 8415
rect 27629 8381 27663 8415
rect 4445 8313 4479 8347
rect 6837 8313 6871 8347
rect 7941 8313 7975 8347
rect 18521 8313 18555 8347
rect 23029 8313 23063 8347
rect 23949 8313 23983 8347
rect 27169 8313 27203 8347
rect 28641 8313 28675 8347
rect 32505 8313 32539 8347
rect 3065 8245 3099 8279
rect 3249 8245 3283 8279
rect 3893 8245 3927 8279
rect 7021 8245 7055 8279
rect 8125 8245 8159 8279
rect 13093 8245 13127 8279
rect 23765 8245 23799 8279
rect 31217 8245 31251 8279
rect 32321 8245 32355 8279
rect 6377 8041 6411 8075
rect 23489 8041 23523 8075
rect 31125 8041 31159 8075
rect 31861 8041 31895 8075
rect 27905 7973 27939 8007
rect 9137 7905 9171 7939
rect 11805 7905 11839 7939
rect 13553 7905 13587 7939
rect 3065 7837 3099 7871
rect 3801 7837 3835 7871
rect 4077 7837 4111 7871
rect 14105 7837 14139 7871
rect 27721 7837 27755 7871
rect 30941 7837 30975 7871
rect 33793 7837 33827 7871
rect 34713 7837 34747 7871
rect 35725 7837 35759 7871
rect 36001 7837 36035 7871
rect 6561 7769 6595 7803
rect 9413 7769 9447 7803
rect 12081 7769 12115 7803
rect 3249 7701 3283 7735
rect 4813 7701 4847 7735
rect 6193 7701 6227 7735
rect 6361 7701 6395 7735
rect 7573 7701 7607 7735
rect 10885 7701 10919 7735
rect 14197 7701 14231 7735
rect 30389 7701 30423 7735
rect 33977 7701 34011 7735
rect 34897 7701 34931 7735
rect 36737 7701 36771 7735
rect 7389 7497 7423 7531
rect 9965 7497 9999 7531
rect 11713 7497 11747 7531
rect 12173 7497 12207 7531
rect 30865 7497 30899 7531
rect 36461 7497 36495 7531
rect 30665 7429 30699 7463
rect 1685 7361 1719 7395
rect 2237 7361 2271 7395
rect 9873 7361 9907 7395
rect 12725 7361 12759 7395
rect 18245 7361 18279 7395
rect 35725 7361 35759 7395
rect 13001 7293 13035 7327
rect 14473 7293 14507 7327
rect 17969 7293 18003 7327
rect 35449 7293 35483 7327
rect 17693 7225 17727 7259
rect 1501 7157 1535 7191
rect 6929 7157 6963 7191
rect 18061 7157 18095 7191
rect 30113 7157 30147 7191
rect 30849 7157 30883 7191
rect 31033 7157 31067 7191
rect 25789 6953 25823 6987
rect 30481 6953 30515 6987
rect 31401 6953 31435 6987
rect 19257 6817 19291 6851
rect 6929 6749 6963 6783
rect 17969 6749 18003 6783
rect 18429 6749 18463 6783
rect 19533 6749 19567 6783
rect 26525 6749 26559 6783
rect 26801 6749 26835 6783
rect 32045 6749 32079 6783
rect 34713 6749 34747 6783
rect 31217 6681 31251 6715
rect 6745 6613 6779 6647
rect 17785 6613 17819 6647
rect 18521 6613 18555 6647
rect 31417 6613 31451 6647
rect 31585 6613 31619 6647
rect 32229 6613 32263 6647
rect 34897 6613 34931 6647
rect 31493 6409 31527 6443
rect 33149 6409 33183 6443
rect 36461 6409 36495 6443
rect 18981 6341 19015 6375
rect 1685 6273 1719 6307
rect 2145 6273 2179 6307
rect 3617 6273 3651 6307
rect 3893 6273 3927 6307
rect 32137 6273 32171 6307
rect 32413 6273 32447 6307
rect 35725 6273 35759 6307
rect 35449 6205 35483 6239
rect 19165 6137 19199 6171
rect 1501 6069 1535 6103
rect 2881 6069 2915 6103
rect 30849 6069 30883 6103
rect 28365 5865 28399 5899
rect 19993 5797 20027 5831
rect 23213 5797 23247 5831
rect 22477 5729 22511 5763
rect 22937 5729 22971 5763
rect 6193 5661 6227 5695
rect 20177 5661 20211 5695
rect 22201 5661 22235 5695
rect 27353 5661 27387 5695
rect 27629 5661 27663 5695
rect 6377 5525 6411 5559
rect 23397 5525 23431 5559
rect 22477 5321 22511 5355
rect 26985 5321 27019 5355
rect 19441 5253 19475 5287
rect 6377 5185 6411 5219
rect 6653 5185 6687 5219
rect 20085 5185 20119 5219
rect 20453 5185 20487 5219
rect 22385 5185 22419 5219
rect 22569 5185 22603 5219
rect 27169 5185 27203 5219
rect 20269 5117 20303 5151
rect 19625 5049 19659 5083
rect 7389 4981 7423 5015
rect 20177 4981 20211 5015
rect 2881 4777 2915 4811
rect 19441 4777 19475 4811
rect 20269 4777 20303 4811
rect 22937 4777 22971 4811
rect 19993 4709 20027 4743
rect 26801 4709 26835 4743
rect 22569 4641 22603 4675
rect 28181 4641 28215 4675
rect 1685 4573 1719 4607
rect 6101 4573 6135 4607
rect 7757 4573 7791 4607
rect 14841 4573 14875 4607
rect 15117 4573 15151 4607
rect 15577 4573 15611 4607
rect 15761 4573 15795 4607
rect 19533 4573 19567 4607
rect 20269 4573 20303 4607
rect 20361 4573 20395 4607
rect 26709 4573 26743 4607
rect 27629 4573 27663 4607
rect 28089 4573 28123 4607
rect 28273 4573 28307 4607
rect 15025 4505 15059 4539
rect 22937 4505 22971 4539
rect 27353 4505 27387 4539
rect 1501 4437 1535 4471
rect 5917 4437 5951 4471
rect 7573 4437 7607 4471
rect 14657 4437 14691 4471
rect 15577 4437 15611 4471
rect 23121 4437 23155 4471
rect 3157 4233 3191 4267
rect 7481 4233 7515 4267
rect 27261 4233 27295 4267
rect 27429 4233 27463 4267
rect 19625 4165 19659 4199
rect 27629 4165 27663 4199
rect 2513 4097 2547 4131
rect 3893 4097 3927 4131
rect 5549 4097 5583 4131
rect 5825 4097 5859 4131
rect 6469 4097 6503 4131
rect 6745 4097 6779 4131
rect 10241 4097 10275 4131
rect 14013 4097 14047 4131
rect 14289 4097 14323 4131
rect 18337 4097 18371 4131
rect 20269 4097 20303 4131
rect 20453 4097 20487 4131
rect 23489 4097 23523 4131
rect 28089 4097 28123 4131
rect 28365 4097 28399 4131
rect 2329 4029 2363 4063
rect 4169 4029 4203 4063
rect 10517 4029 10551 4063
rect 14105 4029 14139 4063
rect 18061 4029 18095 4063
rect 9505 3961 9539 3995
rect 14197 3961 14231 3995
rect 19073 3961 19107 3995
rect 2697 3893 2731 3927
rect 4813 3893 4847 3927
rect 13829 3893 13863 3927
rect 14933 3893 14967 3927
rect 19717 3893 19751 3927
rect 20269 3893 20303 3927
rect 23673 3893 23707 3927
rect 27445 3893 27479 3927
rect 11529 3689 11563 3723
rect 15117 3689 15151 3723
rect 16773 3689 16807 3723
rect 21373 3689 21407 3723
rect 32413 3689 32447 3723
rect 36829 3689 36863 3723
rect 11989 3621 12023 3655
rect 13001 3621 13035 3655
rect 21189 3621 21223 3655
rect 31401 3621 31435 3655
rect 32229 3621 32263 3655
rect 36645 3621 36679 3655
rect 10517 3553 10551 3587
rect 14657 3553 14691 3587
rect 21557 3553 21591 3587
rect 26893 3553 26927 3587
rect 30205 3553 30239 3587
rect 31493 3553 31527 3587
rect 31585 3553 31619 3587
rect 32597 3553 32631 3587
rect 1685 3485 1719 3519
rect 2881 3485 2915 3519
rect 10793 3485 10827 3519
rect 12173 3485 12207 3519
rect 12449 3485 12483 3519
rect 14381 3485 14415 3519
rect 14565 3485 14599 3519
rect 14749 3485 14783 3519
rect 14841 3485 14875 3519
rect 16589 3485 16623 3519
rect 16681 3485 16715 3519
rect 21373 3485 21407 3519
rect 27169 3485 27203 3519
rect 27997 3485 28031 3519
rect 28457 3485 28491 3519
rect 31309 3485 31343 3519
rect 31769 3485 31803 3519
rect 32413 3485 32447 3519
rect 36829 3485 36863 3519
rect 36921 3485 36955 3519
rect 12357 3417 12391 3451
rect 16865 3417 16899 3451
rect 21649 3417 21683 3451
rect 29837 3417 29871 3451
rect 30021 3417 30055 3451
rect 32689 3417 32723 3451
rect 37105 3417 37139 3451
rect 1501 3349 1535 3383
rect 2697 3349 2731 3383
rect 16405 3349 16439 3383
rect 23489 3349 23523 3383
rect 31033 3349 31067 3383
rect 38117 3349 38151 3383
rect 2145 3145 2179 3179
rect 4997 3145 5031 3179
rect 14473 3145 14507 3179
rect 37933 3145 37967 3179
rect 14197 3077 14231 3111
rect 14565 3077 14599 3111
rect 31585 3077 31619 3111
rect 2881 3009 2915 3043
rect 23489 3009 23523 3043
rect 24317 3009 24351 3043
rect 24593 3009 24627 3043
rect 31309 3009 31343 3043
rect 31401 3009 31435 3043
rect 38117 3009 38151 3043
rect 14381 2941 14415 2975
rect 36737 2941 36771 2975
rect 3433 2873 3467 2907
rect 31309 2873 31343 2907
rect 2697 2805 2731 2839
rect 12817 2805 12851 2839
rect 13737 2805 13771 2839
rect 14289 2805 14323 2839
rect 17601 2805 17635 2839
rect 19993 2805 20027 2839
rect 28365 2805 28399 2839
rect 32137 2805 32171 2839
rect 34529 2805 34563 2839
rect 37289 2805 37323 2839
rect 13093 2601 13127 2635
rect 14289 2601 14323 2635
rect 16681 2601 16715 2635
rect 17693 2601 17727 2635
rect 19257 2601 19291 2635
rect 20269 2601 20303 2635
rect 21833 2601 21867 2635
rect 22477 2601 22511 2635
rect 23673 2601 23707 2635
rect 28641 2601 28675 2635
rect 29837 2601 29871 2635
rect 31033 2601 31067 2635
rect 32321 2601 32355 2635
rect 33241 2601 33275 2635
rect 34713 2601 34747 2635
rect 35817 2601 35851 2635
rect 37289 2601 37323 2635
rect 37933 2601 37967 2635
rect 3985 2533 4019 2567
rect 15485 2533 15519 2567
rect 1685 2397 1719 2431
rect 2421 2397 2455 2431
rect 3801 2397 3835 2431
rect 4813 2397 4847 2431
rect 5825 2397 5859 2431
rect 7205 2397 7239 2431
rect 8401 2397 8435 2431
rect 9597 2397 9631 2431
rect 11989 2397 12023 2431
rect 12909 2397 12943 2431
rect 14105 2397 14139 2431
rect 14841 2397 14875 2431
rect 15301 2397 15335 2431
rect 16129 2397 16163 2431
rect 16865 2397 16899 2431
rect 17877 2397 17911 2431
rect 19441 2397 19475 2431
rect 20085 2397 20119 2431
rect 22017 2397 22051 2431
rect 22661 2397 22695 2431
rect 23121 2397 23155 2431
rect 23857 2397 23891 2431
rect 25145 2397 25179 2431
rect 25605 2397 25639 2431
rect 27537 2397 27571 2431
rect 28457 2397 28491 2431
rect 29653 2397 29687 2431
rect 30297 2397 30331 2431
rect 30849 2397 30883 2431
rect 31493 2397 31527 2431
rect 32137 2397 32171 2431
rect 33425 2397 33459 2431
rect 33885 2397 33919 2431
rect 34897 2397 34931 2431
rect 35633 2397 35667 2431
rect 36277 2397 36311 2431
rect 37473 2397 37507 2431
rect 38117 2397 38151 2431
rect 10149 2329 10183 2363
rect 1501 2261 1535 2295
rect 2237 2261 2271 2295
rect 3249 2261 3283 2295
rect 4629 2261 4663 2295
rect 5641 2261 5675 2295
rect 7021 2261 7055 2295
rect 8217 2261 8251 2295
rect 9413 2261 9447 2295
rect 11805 2261 11839 2295
rect 18705 2261 18739 2295
rect 21189 2261 21223 2295
rect 24961 2261 24995 2295
rect 27353 2261 27387 2295
<< metal1 >>
rect 1104 33754 38824 33776
rect 1104 33702 10398 33754
rect 10450 33702 10462 33754
rect 10514 33702 10526 33754
rect 10578 33702 10590 33754
rect 10642 33702 10654 33754
rect 10706 33702 19846 33754
rect 19898 33702 19910 33754
rect 19962 33702 19974 33754
rect 20026 33702 20038 33754
rect 20090 33702 20102 33754
rect 20154 33702 29294 33754
rect 29346 33702 29358 33754
rect 29410 33702 29422 33754
rect 29474 33702 29486 33754
rect 29538 33702 29550 33754
rect 29602 33702 38824 33754
rect 1104 33680 38824 33702
rect 8570 33532 8576 33584
rect 8628 33572 8634 33584
rect 9122 33572 9128 33584
rect 8628 33544 9128 33572
rect 8628 33532 8634 33544
rect 9122 33532 9128 33544
rect 9180 33572 9186 33584
rect 9401 33575 9459 33581
rect 9401 33572 9413 33575
rect 9180 33544 9413 33572
rect 9180 33532 9186 33544
rect 9401 33541 9413 33544
rect 9447 33541 9459 33575
rect 9401 33535 9459 33541
rect 1673 33507 1731 33513
rect 1673 33473 1685 33507
rect 1719 33504 1731 33507
rect 2225 33507 2283 33513
rect 2225 33504 2237 33507
rect 1719 33476 2237 33504
rect 1719 33473 1731 33476
rect 1673 33467 1731 33473
rect 2225 33473 2237 33476
rect 2271 33504 2283 33507
rect 14090 33504 14096 33516
rect 2271 33476 14096 33504
rect 2271 33473 2283 33476
rect 2225 33467 2283 33473
rect 14090 33464 14096 33476
rect 14148 33464 14154 33516
rect 20073 33507 20131 33513
rect 20073 33473 20085 33507
rect 20119 33504 20131 33507
rect 20254 33504 20260 33516
rect 20119 33476 20260 33504
rect 20119 33473 20131 33476
rect 20073 33467 20131 33473
rect 20254 33464 20260 33476
rect 20312 33464 20318 33516
rect 25774 33504 25780 33516
rect 25735 33476 25780 33504
rect 25774 33464 25780 33476
rect 25832 33464 25838 33516
rect 31754 33464 31760 33516
rect 31812 33504 31818 33516
rect 32125 33507 32183 33513
rect 32125 33504 32137 33507
rect 31812 33476 32137 33504
rect 31812 33464 31818 33476
rect 32125 33473 32137 33476
rect 32171 33473 32183 33507
rect 32125 33467 32183 33473
rect 37090 33464 37096 33516
rect 37148 33504 37154 33516
rect 37277 33507 37335 33513
rect 37277 33504 37289 33507
rect 37148 33476 37289 33504
rect 37148 33464 37154 33476
rect 37277 33473 37289 33476
rect 37323 33473 37335 33507
rect 37277 33467 37335 33473
rect 1486 33300 1492 33312
rect 1447 33272 1492 33300
rect 1486 33260 1492 33272
rect 1544 33260 1550 33312
rect 9398 33260 9404 33312
rect 9456 33300 9462 33312
rect 9493 33303 9551 33309
rect 9493 33300 9505 33303
rect 9456 33272 9505 33300
rect 9456 33260 9462 33272
rect 9493 33269 9505 33272
rect 9539 33269 9551 33303
rect 9493 33263 9551 33269
rect 1104 33210 38824 33232
rect 1104 33158 5674 33210
rect 5726 33158 5738 33210
rect 5790 33158 5802 33210
rect 5854 33158 5866 33210
rect 5918 33158 5930 33210
rect 5982 33158 15122 33210
rect 15174 33158 15186 33210
rect 15238 33158 15250 33210
rect 15302 33158 15314 33210
rect 15366 33158 15378 33210
rect 15430 33158 24570 33210
rect 24622 33158 24634 33210
rect 24686 33158 24698 33210
rect 24750 33158 24762 33210
rect 24814 33158 24826 33210
rect 24878 33158 34018 33210
rect 34070 33158 34082 33210
rect 34134 33158 34146 33210
rect 34198 33158 34210 33210
rect 34262 33158 34274 33210
rect 34326 33158 38824 33210
rect 1104 33136 38824 33158
rect 1394 33056 1400 33108
rect 1452 33096 1458 33108
rect 1489 33099 1547 33105
rect 1489 33096 1501 33099
rect 1452 33068 1501 33096
rect 1452 33056 1458 33068
rect 1489 33065 1501 33068
rect 1535 33065 1547 33099
rect 9122 33096 9128 33108
rect 9083 33068 9128 33096
rect 1489 33059 1547 33065
rect 9122 33056 9128 33068
rect 9180 33056 9186 33108
rect 9030 32920 9036 32972
rect 9088 32960 9094 32972
rect 11793 32963 11851 32969
rect 11793 32960 11805 32963
rect 9088 32932 11805 32960
rect 9088 32920 9094 32932
rect 11793 32929 11805 32932
rect 11839 32929 11851 32963
rect 11793 32923 11851 32929
rect 1673 32895 1731 32901
rect 1673 32861 1685 32895
rect 1719 32892 1731 32895
rect 11517 32895 11575 32901
rect 1719 32864 2268 32892
rect 1719 32861 1731 32864
rect 1673 32855 1731 32861
rect 2240 32768 2268 32864
rect 11517 32861 11529 32895
rect 11563 32892 11575 32895
rect 12526 32892 12532 32904
rect 11563 32864 12532 32892
rect 11563 32861 11575 32864
rect 11517 32855 11575 32861
rect 12526 32852 12532 32864
rect 12584 32852 12590 32904
rect 2222 32756 2228 32768
rect 2183 32728 2228 32756
rect 2222 32716 2228 32728
rect 2280 32716 2286 32768
rect 1104 32666 38824 32688
rect 1104 32614 10398 32666
rect 10450 32614 10462 32666
rect 10514 32614 10526 32666
rect 10578 32614 10590 32666
rect 10642 32614 10654 32666
rect 10706 32614 19846 32666
rect 19898 32614 19910 32666
rect 19962 32614 19974 32666
rect 20026 32614 20038 32666
rect 20090 32614 20102 32666
rect 20154 32614 29294 32666
rect 29346 32614 29358 32666
rect 29410 32614 29422 32666
rect 29474 32614 29486 32666
rect 29538 32614 29550 32666
rect 29602 32614 38824 32666
rect 1104 32592 38824 32614
rect 2222 32512 2228 32564
rect 2280 32552 2286 32564
rect 12894 32552 12900 32564
rect 2280 32524 12900 32552
rect 2280 32512 2286 32524
rect 12894 32512 12900 32524
rect 12952 32512 12958 32564
rect 9030 32484 9036 32496
rect 6472 32456 9036 32484
rect 3326 32416 3332 32428
rect 3287 32388 3332 32416
rect 3326 32376 3332 32388
rect 3384 32376 3390 32428
rect 3605 32351 3663 32357
rect 3605 32317 3617 32351
rect 3651 32348 3663 32351
rect 3970 32348 3976 32360
rect 3651 32320 3976 32348
rect 3651 32317 3663 32320
rect 3605 32311 3663 32317
rect 3970 32308 3976 32320
rect 4028 32348 4034 32360
rect 6472 32357 6500 32456
rect 9030 32444 9036 32456
rect 9088 32444 9094 32496
rect 17218 32444 17224 32496
rect 17276 32484 17282 32496
rect 17276 32456 17724 32484
rect 17276 32444 17282 32456
rect 6638 32376 6644 32428
rect 6696 32416 6702 32428
rect 11790 32425 11796 32428
rect 6733 32419 6791 32425
rect 6733 32416 6745 32419
rect 6696 32388 6745 32416
rect 6696 32376 6702 32388
rect 6733 32385 6745 32388
rect 6779 32385 6791 32419
rect 6733 32379 6791 32385
rect 11784 32379 11796 32425
rect 11848 32416 11854 32428
rect 11848 32388 11884 32416
rect 11790 32376 11796 32379
rect 11848 32376 11854 32388
rect 16390 32376 16396 32428
rect 16448 32416 16454 32428
rect 17696 32425 17724 32456
rect 17405 32419 17463 32425
rect 17405 32416 17417 32419
rect 16448 32388 17417 32416
rect 16448 32376 16454 32388
rect 17405 32385 17417 32388
rect 17451 32385 17463 32419
rect 17405 32379 17463 32385
rect 17681 32419 17739 32425
rect 17681 32385 17693 32419
rect 17727 32385 17739 32419
rect 17681 32379 17739 32385
rect 6457 32351 6515 32357
rect 6457 32348 6469 32351
rect 4028 32320 6469 32348
rect 4028 32308 4034 32320
rect 6457 32317 6469 32320
rect 6503 32317 6515 32351
rect 11517 32351 11575 32357
rect 11517 32348 11529 32351
rect 6457 32311 6515 32317
rect 10888 32320 11529 32348
rect 10888 32224 10916 32320
rect 11517 32317 11529 32320
rect 11563 32317 11575 32351
rect 11517 32311 11575 32317
rect 1762 32172 1768 32224
rect 1820 32212 1826 32224
rect 2593 32215 2651 32221
rect 2593 32212 2605 32215
rect 1820 32184 2605 32212
rect 1820 32172 1826 32184
rect 2593 32181 2605 32184
rect 2639 32212 2651 32215
rect 4982 32212 4988 32224
rect 2639 32184 4988 32212
rect 2639 32181 2651 32184
rect 2593 32175 2651 32181
rect 4982 32172 4988 32184
rect 5040 32212 5046 32224
rect 7469 32215 7527 32221
rect 7469 32212 7481 32215
rect 5040 32184 7481 32212
rect 5040 32172 5046 32184
rect 7469 32181 7481 32184
rect 7515 32212 7527 32215
rect 8018 32212 8024 32224
rect 7515 32184 8024 32212
rect 7515 32181 7527 32184
rect 7469 32175 7527 32181
rect 8018 32172 8024 32184
rect 8076 32172 8082 32224
rect 10870 32212 10876 32224
rect 10831 32184 10876 32212
rect 10870 32172 10876 32184
rect 10928 32172 10934 32224
rect 12894 32212 12900 32224
rect 12855 32184 12900 32212
rect 12894 32172 12900 32184
rect 12952 32172 12958 32224
rect 16669 32215 16727 32221
rect 16669 32181 16681 32215
rect 16715 32212 16727 32215
rect 18322 32212 18328 32224
rect 16715 32184 18328 32212
rect 16715 32181 16727 32184
rect 16669 32175 16727 32181
rect 18322 32172 18328 32184
rect 18380 32212 18386 32224
rect 22370 32212 22376 32224
rect 18380 32184 22376 32212
rect 18380 32172 18386 32184
rect 22370 32172 22376 32184
rect 22428 32172 22434 32224
rect 1104 32122 38824 32144
rect 1104 32070 5674 32122
rect 5726 32070 5738 32122
rect 5790 32070 5802 32122
rect 5854 32070 5866 32122
rect 5918 32070 5930 32122
rect 5982 32070 15122 32122
rect 15174 32070 15186 32122
rect 15238 32070 15250 32122
rect 15302 32070 15314 32122
rect 15366 32070 15378 32122
rect 15430 32070 24570 32122
rect 24622 32070 24634 32122
rect 24686 32070 24698 32122
rect 24750 32070 24762 32122
rect 24814 32070 24826 32122
rect 24878 32070 34018 32122
rect 34070 32070 34082 32122
rect 34134 32070 34146 32122
rect 34198 32070 34210 32122
rect 34262 32070 34274 32122
rect 34326 32070 38824 32122
rect 1104 32048 38824 32070
rect 2869 32011 2927 32017
rect 2869 31977 2881 32011
rect 2915 32008 2927 32011
rect 3326 32008 3332 32020
rect 2915 31980 3332 32008
rect 2915 31977 2927 31980
rect 2869 31971 2927 31977
rect 3326 31968 3332 31980
rect 3384 31968 3390 32020
rect 6638 32008 6644 32020
rect 6599 31980 6644 32008
rect 6638 31968 6644 31980
rect 6696 31968 6702 32020
rect 18782 32008 18788 32020
rect 6886 31980 18788 32008
rect 2225 31943 2283 31949
rect 2225 31909 2237 31943
rect 2271 31940 2283 31943
rect 6886 31940 6914 31980
rect 18782 31968 18788 31980
rect 18840 31968 18846 32020
rect 23474 32008 23480 32020
rect 21376 31980 23480 32008
rect 2271 31912 6914 31940
rect 2271 31909 2283 31912
rect 2225 31903 2283 31909
rect 1673 31807 1731 31813
rect 1673 31773 1685 31807
rect 1719 31804 1731 31807
rect 2240 31804 2268 31903
rect 8018 31900 8024 31952
rect 8076 31940 8082 31952
rect 11514 31940 11520 31952
rect 8076 31912 11520 31940
rect 8076 31900 8082 31912
rect 11514 31900 11520 31912
rect 11572 31900 11578 31952
rect 16390 31940 16396 31952
rect 16351 31912 16396 31940
rect 16390 31900 16396 31912
rect 16448 31900 16454 31952
rect 18322 31940 18328 31952
rect 18283 31912 18328 31940
rect 18322 31900 18328 31912
rect 18380 31900 18386 31952
rect 20901 31943 20959 31949
rect 20901 31909 20913 31943
rect 20947 31909 20959 31943
rect 20901 31903 20959 31909
rect 12526 31832 12532 31884
rect 12584 31872 12590 31884
rect 12584 31844 12629 31872
rect 12584 31832 12590 31844
rect 2682 31804 2688 31816
rect 1719 31776 2268 31804
rect 2643 31776 2688 31804
rect 1719 31773 1731 31776
rect 1673 31767 1731 31773
rect 2682 31764 2688 31776
rect 2740 31764 2746 31816
rect 6454 31804 6460 31816
rect 6415 31776 6460 31804
rect 6454 31764 6460 31776
rect 6512 31764 6518 31816
rect 9122 31804 9128 31816
rect 9083 31776 9128 31804
rect 9122 31764 9128 31776
rect 9180 31764 9186 31816
rect 12250 31804 12256 31816
rect 12211 31776 12256 31804
rect 12250 31764 12256 31776
rect 12308 31764 12314 31816
rect 16206 31804 16212 31816
rect 16167 31776 16212 31804
rect 16206 31764 16212 31776
rect 16264 31764 16270 31816
rect 17218 31764 17224 31816
rect 17276 31804 17282 31816
rect 17313 31807 17371 31813
rect 17313 31804 17325 31807
rect 17276 31776 17325 31804
rect 17276 31764 17282 31776
rect 17313 31773 17325 31776
rect 17359 31773 17371 31807
rect 17586 31804 17592 31816
rect 17547 31776 17592 31804
rect 17313 31767 17371 31773
rect 17586 31764 17592 31776
rect 17644 31764 17650 31816
rect 20714 31804 20720 31816
rect 20675 31776 20720 31804
rect 20714 31764 20720 31776
rect 20772 31764 20778 31816
rect 20916 31804 20944 31903
rect 21376 31881 21404 31980
rect 23474 31968 23480 31980
rect 23532 32008 23538 32020
rect 23532 31980 23888 32008
rect 23532 31968 23538 31980
rect 22370 31940 22376 31952
rect 22331 31912 22376 31940
rect 22370 31900 22376 31912
rect 22428 31940 22434 31952
rect 22833 31943 22891 31949
rect 22833 31940 22845 31943
rect 22428 31912 22845 31940
rect 22428 31900 22434 31912
rect 22833 31909 22845 31912
rect 22879 31909 22891 31943
rect 22833 31903 22891 31909
rect 23860 31881 23888 31980
rect 25406 31968 25412 32020
rect 25464 32008 25470 32020
rect 26053 32011 26111 32017
rect 26053 32008 26065 32011
rect 25464 31980 26065 32008
rect 25464 31968 25470 31980
rect 26053 31977 26065 31980
rect 26099 32008 26111 32011
rect 28994 32008 29000 32020
rect 26099 31980 29000 32008
rect 26099 31977 26111 31980
rect 26053 31971 26111 31977
rect 28994 31968 29000 31980
rect 29052 31968 29058 32020
rect 21361 31875 21419 31881
rect 21361 31841 21373 31875
rect 21407 31841 21419 31875
rect 21361 31835 21419 31841
rect 23845 31875 23903 31881
rect 23845 31841 23857 31875
rect 23891 31841 23903 31875
rect 23845 31835 23903 31841
rect 21637 31807 21695 31813
rect 21637 31804 21649 31807
rect 20916 31776 21312 31804
rect 21284 31736 21312 31776
rect 21468 31776 21649 31804
rect 21468 31736 21496 31776
rect 21637 31773 21649 31776
rect 21683 31773 21695 31807
rect 21637 31767 21695 31773
rect 22094 31764 22100 31816
rect 22152 31804 22158 31816
rect 23569 31807 23627 31813
rect 23569 31804 23581 31807
rect 22152 31776 23581 31804
rect 22152 31764 22158 31776
rect 23569 31773 23581 31776
rect 23615 31773 23627 31807
rect 25038 31804 25044 31816
rect 24999 31776 25044 31804
rect 23569 31767 23627 31773
rect 25038 31764 25044 31776
rect 25096 31764 25102 31816
rect 25314 31804 25320 31816
rect 25275 31776 25320 31804
rect 25314 31764 25320 31776
rect 25372 31764 25378 31816
rect 27985 31807 28043 31813
rect 27985 31773 27997 31807
rect 28031 31773 28043 31807
rect 28258 31804 28264 31816
rect 28219 31776 28264 31804
rect 27985 31767 28043 31773
rect 21284 31708 21496 31736
rect 25056 31736 25084 31764
rect 28000 31736 28028 31767
rect 28258 31764 28264 31776
rect 28316 31764 28322 31816
rect 28166 31736 28172 31748
rect 25056 31708 28172 31736
rect 28166 31696 28172 31708
rect 28224 31696 28230 31748
rect 1486 31668 1492 31680
rect 1447 31640 1492 31668
rect 1486 31628 1492 31640
rect 1544 31628 1550 31680
rect 8754 31628 8760 31680
rect 8812 31668 8818 31680
rect 8941 31671 8999 31677
rect 8941 31668 8953 31671
rect 8812 31640 8953 31668
rect 8812 31628 8818 31640
rect 8941 31637 8953 31640
rect 8987 31637 8999 31671
rect 8941 31631 8999 31637
rect 1104 31578 38824 31600
rect 1104 31526 10398 31578
rect 10450 31526 10462 31578
rect 10514 31526 10526 31578
rect 10578 31526 10590 31578
rect 10642 31526 10654 31578
rect 10706 31526 19846 31578
rect 19898 31526 19910 31578
rect 19962 31526 19974 31578
rect 20026 31526 20038 31578
rect 20090 31526 20102 31578
rect 20154 31526 29294 31578
rect 29346 31526 29358 31578
rect 29410 31526 29422 31578
rect 29474 31526 29486 31578
rect 29538 31526 29550 31578
rect 29602 31526 38824 31578
rect 1104 31504 38824 31526
rect 2682 31464 2688 31476
rect 2643 31436 2688 31464
rect 2682 31424 2688 31436
rect 2740 31424 2746 31476
rect 6454 31424 6460 31476
rect 6512 31464 6518 31476
rect 6733 31467 6791 31473
rect 6733 31464 6745 31467
rect 6512 31436 6745 31464
rect 6512 31424 6518 31436
rect 6733 31433 6745 31436
rect 6779 31433 6791 31467
rect 8018 31464 8024 31476
rect 7979 31436 8024 31464
rect 6733 31427 6791 31433
rect 8018 31424 8024 31436
rect 8076 31424 8082 31476
rect 11885 31467 11943 31473
rect 11885 31433 11897 31467
rect 11931 31464 11943 31467
rect 12250 31464 12256 31476
rect 11931 31436 12256 31464
rect 11931 31433 11943 31436
rect 11885 31427 11943 31433
rect 12250 31424 12256 31436
rect 12308 31424 12314 31476
rect 15197 31467 15255 31473
rect 15197 31433 15209 31467
rect 15243 31464 15255 31467
rect 16206 31464 16212 31476
rect 15243 31436 16212 31464
rect 15243 31433 15255 31436
rect 15197 31427 15255 31433
rect 16206 31424 16212 31436
rect 16264 31424 16270 31476
rect 16853 31467 16911 31473
rect 16853 31433 16865 31467
rect 16899 31464 16911 31467
rect 17586 31464 17592 31476
rect 16899 31436 17592 31464
rect 16899 31433 16911 31436
rect 16853 31427 16911 31433
rect 17586 31424 17592 31436
rect 17644 31424 17650 31476
rect 20441 31467 20499 31473
rect 20441 31433 20453 31467
rect 20487 31464 20499 31467
rect 20714 31464 20720 31476
rect 20487 31436 20720 31464
rect 20487 31433 20499 31436
rect 20441 31427 20499 31433
rect 20714 31424 20720 31436
rect 20772 31424 20778 31476
rect 22005 31467 22063 31473
rect 22005 31433 22017 31467
rect 22051 31464 22063 31467
rect 22094 31464 22100 31476
rect 22051 31436 22100 31464
rect 22051 31433 22063 31436
rect 22005 31427 22063 31433
rect 22094 31424 22100 31436
rect 22152 31424 22158 31476
rect 28994 31424 29000 31476
rect 29052 31464 29058 31476
rect 29273 31467 29331 31473
rect 29273 31464 29285 31467
rect 29052 31436 29285 31464
rect 29052 31424 29058 31436
rect 29273 31433 29285 31436
rect 29319 31433 29331 31467
rect 29273 31427 29331 31433
rect 15856 31368 20300 31396
rect 15856 31340 15884 31368
rect 2869 31331 2927 31337
rect 2869 31297 2881 31331
rect 2915 31328 2927 31331
rect 3418 31328 3424 31340
rect 2915 31300 3424 31328
rect 2915 31297 2927 31300
rect 2869 31291 2927 31297
rect 3418 31288 3424 31300
rect 3476 31328 3482 31340
rect 6546 31328 6552 31340
rect 3476 31300 6552 31328
rect 3476 31288 3482 31300
rect 6546 31288 6552 31300
rect 6604 31288 6610 31340
rect 8754 31328 8760 31340
rect 8715 31300 8760 31328
rect 8754 31288 8760 31300
rect 8812 31288 8818 31340
rect 9030 31328 9036 31340
rect 8991 31300 9036 31328
rect 9030 31288 9036 31300
rect 9088 31288 9094 31340
rect 11698 31328 11704 31340
rect 11659 31300 11704 31328
rect 11698 31288 11704 31300
rect 11756 31288 11762 31340
rect 15013 31331 15071 31337
rect 15013 31297 15025 31331
rect 15059 31328 15071 31331
rect 15838 31328 15844 31340
rect 15059 31300 15844 31328
rect 15059 31297 15071 31300
rect 15013 31291 15071 31297
rect 15838 31288 15844 31300
rect 15896 31288 15902 31340
rect 20272 31337 20300 31368
rect 16025 31331 16083 31337
rect 16025 31297 16037 31331
rect 16071 31328 16083 31331
rect 16669 31331 16727 31337
rect 16669 31328 16681 31331
rect 16071 31300 16681 31328
rect 16071 31297 16083 31300
rect 16025 31291 16083 31297
rect 16669 31297 16681 31300
rect 16715 31297 16727 31331
rect 16669 31291 16727 31297
rect 20257 31331 20315 31337
rect 20257 31297 20269 31331
rect 20303 31328 20315 31331
rect 21174 31328 21180 31340
rect 20303 31300 21180 31328
rect 20303 31297 20315 31300
rect 20257 31291 20315 31297
rect 21174 31288 21180 31300
rect 21232 31288 21238 31340
rect 21358 31288 21364 31340
rect 21416 31328 21422 31340
rect 21821 31331 21879 31337
rect 21821 31328 21833 31331
rect 21416 31300 21833 31328
rect 21416 31288 21422 31300
rect 21821 31297 21833 31300
rect 21867 31297 21879 31331
rect 21821 31291 21879 31297
rect 28537 31331 28595 31337
rect 28537 31297 28549 31331
rect 28583 31328 28595 31331
rect 29546 31328 29552 31340
rect 28583 31300 29552 31328
rect 28583 31297 28595 31300
rect 28537 31291 28595 31297
rect 29546 31288 29552 31300
rect 29604 31288 29610 31340
rect 3053 31263 3111 31269
rect 3053 31229 3065 31263
rect 3099 31260 3111 31263
rect 3142 31260 3148 31272
rect 3099 31232 3148 31260
rect 3099 31229 3111 31232
rect 3053 31223 3111 31229
rect 3142 31220 3148 31232
rect 3200 31260 3206 31272
rect 3513 31263 3571 31269
rect 3513 31260 3525 31263
rect 3200 31232 3525 31260
rect 3200 31220 3206 31232
rect 3513 31229 3525 31232
rect 3559 31229 3571 31263
rect 3513 31223 3571 31229
rect 6365 31263 6423 31269
rect 6365 31229 6377 31263
rect 6411 31260 6423 31263
rect 6914 31260 6920 31272
rect 6411 31232 6920 31260
rect 6411 31229 6423 31232
rect 6365 31223 6423 31229
rect 6914 31220 6920 31232
rect 6972 31220 6978 31272
rect 13170 31220 13176 31272
rect 13228 31260 13234 31272
rect 14829 31263 14887 31269
rect 14829 31260 14841 31263
rect 13228 31232 14841 31260
rect 13228 31220 13234 31232
rect 14829 31229 14841 31232
rect 14875 31229 14887 31263
rect 15654 31260 15660 31272
rect 15615 31232 15660 31260
rect 14829 31223 14887 31229
rect 15654 31220 15660 31232
rect 15712 31220 15718 31272
rect 19518 31220 19524 31272
rect 19576 31260 19582 31272
rect 19613 31263 19671 31269
rect 19613 31260 19625 31263
rect 19576 31232 19625 31260
rect 19576 31220 19582 31232
rect 19613 31229 19625 31232
rect 19659 31260 19671 31263
rect 20073 31263 20131 31269
rect 20073 31260 20085 31263
rect 19659 31232 20085 31260
rect 19659 31229 19671 31232
rect 19613 31223 19671 31229
rect 20073 31229 20085 31232
rect 20119 31229 20131 31263
rect 20073 31223 20131 31229
rect 28166 31220 28172 31272
rect 28224 31260 28230 31272
rect 28261 31263 28319 31269
rect 28261 31260 28273 31263
rect 28224 31232 28273 31260
rect 28224 31220 28230 31232
rect 28261 31229 28273 31232
rect 28307 31229 28319 31263
rect 28261 31223 28319 31229
rect 1104 31034 38824 31056
rect 1104 30982 5674 31034
rect 5726 30982 5738 31034
rect 5790 30982 5802 31034
rect 5854 30982 5866 31034
rect 5918 30982 5930 31034
rect 5982 30982 15122 31034
rect 15174 30982 15186 31034
rect 15238 30982 15250 31034
rect 15302 30982 15314 31034
rect 15366 30982 15378 31034
rect 15430 30982 24570 31034
rect 24622 30982 24634 31034
rect 24686 30982 24698 31034
rect 24750 30982 24762 31034
rect 24814 30982 24826 31034
rect 24878 30982 34018 31034
rect 34070 30982 34082 31034
rect 34134 30982 34146 31034
rect 34198 30982 34210 31034
rect 34262 30982 34274 31034
rect 34326 30982 38824 31034
rect 1104 30960 38824 30982
rect 4982 30920 4988 30932
rect 4943 30892 4988 30920
rect 4982 30880 4988 30892
rect 5040 30880 5046 30932
rect 8941 30923 8999 30929
rect 8941 30889 8953 30923
rect 8987 30920 8999 30923
rect 9122 30920 9128 30932
rect 8987 30892 9128 30920
rect 8987 30889 8999 30892
rect 8941 30883 8999 30889
rect 9122 30880 9128 30892
rect 9180 30880 9186 30932
rect 15565 30923 15623 30929
rect 15565 30889 15577 30923
rect 15611 30920 15623 30923
rect 15654 30920 15660 30932
rect 15611 30892 15660 30920
rect 15611 30889 15623 30892
rect 15565 30883 15623 30889
rect 15654 30880 15660 30892
rect 15712 30880 15718 30932
rect 21358 30920 21364 30932
rect 21319 30892 21364 30920
rect 21358 30880 21364 30892
rect 21416 30880 21422 30932
rect 24765 30923 24823 30929
rect 24765 30889 24777 30923
rect 24811 30920 24823 30923
rect 25038 30920 25044 30932
rect 24811 30892 25044 30920
rect 24811 30889 24823 30892
rect 24765 30883 24823 30889
rect 25038 30880 25044 30892
rect 25096 30880 25102 30932
rect 25314 30880 25320 30932
rect 25372 30920 25378 30932
rect 25409 30923 25467 30929
rect 25409 30920 25421 30923
rect 25372 30892 25421 30920
rect 25372 30880 25378 30892
rect 25409 30889 25421 30892
rect 25455 30889 25467 30923
rect 25409 30883 25467 30889
rect 28258 30880 28264 30932
rect 28316 30920 28322 30932
rect 28629 30923 28687 30929
rect 28629 30920 28641 30923
rect 28316 30892 28641 30920
rect 28316 30880 28322 30892
rect 28629 30889 28641 30892
rect 28675 30889 28687 30923
rect 29546 30920 29552 30932
rect 29507 30892 29552 30920
rect 28629 30883 28687 30889
rect 29546 30880 29552 30892
rect 29604 30880 29610 30932
rect 3970 30784 3976 30796
rect 3931 30756 3976 30784
rect 3970 30744 3976 30756
rect 4028 30744 4034 30796
rect 6914 30744 6920 30796
rect 6972 30784 6978 30796
rect 12710 30784 12716 30796
rect 6972 30756 12716 30784
rect 6972 30744 6978 30756
rect 12710 30744 12716 30756
rect 12768 30784 12774 30796
rect 13170 30784 13176 30796
rect 12768 30756 13176 30784
rect 12768 30744 12774 30756
rect 13170 30744 13176 30756
rect 13228 30744 13234 30796
rect 23934 30784 23940 30796
rect 22066 30756 23940 30784
rect 1670 30716 1676 30728
rect 1631 30688 1676 30716
rect 1670 30676 1676 30688
rect 1728 30676 1734 30728
rect 4246 30716 4252 30728
rect 4207 30688 4252 30716
rect 4246 30676 4252 30688
rect 4304 30676 4310 30728
rect 6546 30676 6552 30728
rect 6604 30716 6610 30728
rect 9125 30719 9183 30725
rect 9125 30716 9137 30719
rect 6604 30688 9137 30716
rect 6604 30676 6610 30688
rect 9125 30685 9137 30688
rect 9171 30685 9183 30719
rect 9125 30679 9183 30685
rect 9309 30719 9367 30725
rect 9309 30685 9321 30719
rect 9355 30716 9367 30719
rect 9858 30716 9864 30728
rect 9355 30688 9864 30716
rect 9355 30685 9367 30688
rect 9309 30679 9367 30685
rect 9140 30648 9168 30679
rect 9858 30676 9864 30688
rect 9916 30676 9922 30728
rect 20806 30676 20812 30728
rect 20864 30716 20870 30728
rect 20993 30719 21051 30725
rect 20993 30716 21005 30719
rect 20864 30688 21005 30716
rect 20864 30676 20870 30688
rect 20993 30685 21005 30688
rect 21039 30685 21051 30719
rect 21174 30716 21180 30728
rect 21135 30688 21180 30716
rect 20993 30679 21051 30685
rect 11790 30648 11796 30660
rect 9140 30620 11796 30648
rect 11790 30608 11796 30620
rect 11848 30608 11854 30660
rect 21008 30648 21036 30679
rect 21174 30676 21180 30688
rect 21232 30676 21238 30728
rect 21821 30651 21879 30657
rect 21821 30648 21833 30651
rect 21008 30620 21833 30648
rect 21821 30617 21833 30620
rect 21867 30648 21879 30651
rect 22066 30648 22094 30756
rect 23934 30744 23940 30756
rect 23992 30744 23998 30796
rect 24486 30676 24492 30728
rect 24544 30716 24550 30728
rect 24581 30719 24639 30725
rect 24581 30716 24593 30719
rect 24544 30688 24593 30716
rect 24544 30676 24550 30688
rect 24581 30685 24593 30688
rect 24627 30685 24639 30719
rect 25222 30716 25228 30728
rect 25183 30688 25228 30716
rect 24581 30679 24639 30685
rect 25222 30676 25228 30688
rect 25280 30676 25286 30728
rect 28810 30716 28816 30728
rect 28771 30688 28816 30716
rect 28810 30676 28816 30688
rect 28868 30676 28874 30728
rect 29730 30716 29736 30728
rect 29691 30688 29736 30716
rect 29730 30676 29736 30688
rect 29788 30676 29794 30728
rect 21867 30620 22094 30648
rect 21867 30617 21879 30620
rect 21821 30611 21879 30617
rect 1486 30580 1492 30592
rect 1447 30552 1492 30580
rect 1486 30540 1492 30552
rect 1544 30540 1550 30592
rect 9858 30580 9864 30592
rect 9819 30552 9864 30580
rect 9858 30540 9864 30552
rect 9916 30540 9922 30592
rect 1104 30490 38824 30512
rect 1104 30438 10398 30490
rect 10450 30438 10462 30490
rect 10514 30438 10526 30490
rect 10578 30438 10590 30490
rect 10642 30438 10654 30490
rect 10706 30438 19846 30490
rect 19898 30438 19910 30490
rect 19962 30438 19974 30490
rect 20026 30438 20038 30490
rect 20090 30438 20102 30490
rect 20154 30438 29294 30490
rect 29346 30438 29358 30490
rect 29410 30438 29422 30490
rect 29474 30438 29486 30490
rect 29538 30438 29550 30490
rect 29602 30438 38824 30490
rect 1104 30416 38824 30438
rect 4246 30376 4252 30388
rect 4207 30348 4252 30376
rect 4246 30336 4252 30348
rect 4304 30336 4310 30388
rect 11698 30336 11704 30388
rect 11756 30376 11762 30388
rect 11885 30379 11943 30385
rect 11885 30376 11897 30379
rect 11756 30348 11897 30376
rect 11756 30336 11762 30348
rect 11885 30345 11897 30348
rect 11931 30345 11943 30379
rect 11885 30339 11943 30345
rect 3418 30240 3424 30252
rect 3379 30212 3424 30240
rect 3418 30200 3424 30212
rect 3476 30200 3482 30252
rect 3605 30243 3663 30249
rect 3605 30209 3617 30243
rect 3651 30240 3663 30243
rect 4065 30243 4123 30249
rect 4065 30240 4077 30243
rect 3651 30212 4077 30240
rect 3651 30209 3663 30212
rect 3605 30203 3663 30209
rect 4065 30209 4077 30212
rect 4111 30209 4123 30243
rect 4065 30203 4123 30209
rect 11701 30243 11759 30249
rect 11701 30209 11713 30243
rect 11747 30240 11759 30243
rect 12434 30240 12440 30252
rect 11747 30212 12440 30240
rect 11747 30209 11759 30212
rect 11701 30203 11759 30209
rect 12434 30200 12440 30212
rect 12492 30200 12498 30252
rect 24394 30200 24400 30252
rect 24452 30240 24458 30252
rect 24765 30243 24823 30249
rect 24765 30240 24777 30243
rect 24452 30212 24777 30240
rect 24452 30200 24458 30212
rect 24765 30209 24777 30212
rect 24811 30209 24823 30243
rect 24765 30203 24823 30209
rect 3237 30175 3295 30181
rect 3237 30141 3249 30175
rect 3283 30172 3295 30175
rect 4154 30172 4160 30184
rect 3283 30144 4160 30172
rect 3283 30141 3295 30144
rect 3237 30135 3295 30141
rect 4154 30132 4160 30144
rect 4212 30132 4218 30184
rect 11517 30175 11575 30181
rect 11517 30141 11529 30175
rect 11563 30172 11575 30175
rect 13814 30172 13820 30184
rect 11563 30144 13820 30172
rect 11563 30141 11575 30144
rect 11517 30135 11575 30141
rect 13814 30132 13820 30144
rect 13872 30132 13878 30184
rect 24486 30172 24492 30184
rect 24447 30144 24492 30172
rect 24486 30132 24492 30144
rect 24544 30132 24550 30184
rect 12434 29996 12440 30048
rect 12492 30036 12498 30048
rect 12492 30008 12537 30036
rect 12492 29996 12498 30008
rect 25406 29996 25412 30048
rect 25464 30036 25470 30048
rect 25501 30039 25559 30045
rect 25501 30036 25513 30039
rect 25464 30008 25513 30036
rect 25464 29996 25470 30008
rect 25501 30005 25513 30008
rect 25547 30005 25559 30039
rect 25501 29999 25559 30005
rect 1104 29946 38824 29968
rect 1104 29894 5674 29946
rect 5726 29894 5738 29946
rect 5790 29894 5802 29946
rect 5854 29894 5866 29946
rect 5918 29894 5930 29946
rect 5982 29894 15122 29946
rect 15174 29894 15186 29946
rect 15238 29894 15250 29946
rect 15302 29894 15314 29946
rect 15366 29894 15378 29946
rect 15430 29894 24570 29946
rect 24622 29894 24634 29946
rect 24686 29894 24698 29946
rect 24750 29894 24762 29946
rect 24814 29894 24826 29946
rect 24878 29894 34018 29946
rect 34070 29894 34082 29946
rect 34134 29894 34146 29946
rect 34198 29894 34210 29946
rect 34262 29894 34274 29946
rect 34326 29894 38824 29946
rect 1104 29872 38824 29894
rect 1670 29792 1676 29844
rect 1728 29832 1734 29844
rect 2593 29835 2651 29841
rect 2593 29832 2605 29835
rect 1728 29804 2605 29832
rect 1728 29792 1734 29804
rect 2593 29801 2605 29804
rect 2639 29801 2651 29835
rect 2593 29795 2651 29801
rect 11514 29792 11520 29844
rect 11572 29832 11578 29844
rect 11793 29835 11851 29841
rect 11793 29832 11805 29835
rect 11572 29804 11805 29832
rect 11572 29792 11578 29804
rect 11793 29801 11805 29804
rect 11839 29801 11851 29835
rect 11793 29795 11851 29801
rect 25133 29835 25191 29841
rect 25133 29801 25145 29835
rect 25179 29832 25191 29835
rect 25222 29832 25228 29844
rect 25179 29804 25228 29832
rect 25179 29801 25191 29804
rect 25133 29795 25191 29801
rect 25222 29792 25228 29804
rect 25280 29792 25286 29844
rect 28721 29835 28779 29841
rect 28721 29801 28733 29835
rect 28767 29832 28779 29835
rect 28810 29832 28816 29844
rect 28767 29804 28816 29832
rect 28767 29801 28779 29804
rect 28721 29795 28779 29801
rect 28810 29792 28816 29804
rect 28868 29792 28874 29844
rect 24964 29736 26188 29764
rect 23934 29656 23940 29708
rect 23992 29696 23998 29708
rect 24762 29696 24768 29708
rect 23992 29668 24768 29696
rect 23992 29656 23998 29668
rect 24762 29656 24768 29668
rect 24820 29656 24826 29708
rect 2777 29631 2835 29637
rect 2777 29597 2789 29631
rect 2823 29628 2835 29631
rect 2958 29628 2964 29640
rect 2823 29600 2964 29628
rect 2823 29597 2835 29600
rect 2777 29591 2835 29597
rect 2958 29588 2964 29600
rect 3016 29588 3022 29640
rect 12526 29628 12532 29640
rect 12487 29600 12532 29628
rect 12526 29588 12532 29600
rect 12584 29588 12590 29640
rect 12618 29588 12624 29640
rect 12676 29628 12682 29640
rect 12805 29631 12863 29637
rect 12805 29628 12817 29631
rect 12676 29600 12817 29628
rect 12676 29588 12682 29600
rect 12805 29597 12817 29600
rect 12851 29597 12863 29631
rect 12805 29591 12863 29597
rect 24118 29588 24124 29640
rect 24176 29628 24182 29640
rect 24964 29637 24992 29736
rect 24949 29631 25007 29637
rect 24949 29628 24961 29631
rect 24176 29600 24961 29628
rect 24176 29588 24182 29600
rect 24949 29597 24961 29600
rect 24995 29597 25007 29631
rect 26160 29628 26188 29736
rect 28368 29668 28580 29696
rect 28368 29628 28396 29668
rect 28552 29637 28580 29668
rect 26160 29600 28396 29628
rect 28445 29631 28503 29637
rect 24949 29591 25007 29597
rect 28445 29597 28457 29631
rect 28491 29597 28503 29631
rect 28445 29591 28503 29597
rect 28537 29631 28595 29637
rect 28537 29597 28549 29631
rect 28583 29628 28595 29631
rect 28902 29628 28908 29640
rect 28583 29600 28908 29628
rect 28583 29597 28595 29600
rect 28537 29591 28595 29597
rect 24762 29520 24768 29572
rect 24820 29560 24826 29572
rect 25593 29563 25651 29569
rect 25593 29560 25605 29563
rect 24820 29532 25605 29560
rect 24820 29520 24826 29532
rect 25593 29529 25605 29532
rect 25639 29560 25651 29563
rect 28460 29560 28488 29591
rect 28902 29588 28908 29600
rect 28960 29588 28966 29640
rect 29549 29563 29607 29569
rect 29549 29560 29561 29563
rect 25639 29532 26234 29560
rect 28460 29532 29561 29560
rect 25639 29529 25651 29532
rect 25593 29523 25651 29529
rect 3881 29495 3939 29501
rect 3881 29461 3893 29495
rect 3927 29492 3939 29495
rect 4154 29492 4160 29504
rect 3927 29464 4160 29492
rect 3927 29461 3939 29464
rect 3881 29455 3939 29461
rect 4154 29452 4160 29464
rect 4212 29492 4218 29504
rect 4614 29492 4620 29504
rect 4212 29464 4620 29492
rect 4212 29452 4218 29464
rect 4614 29452 4620 29464
rect 4672 29452 4678 29504
rect 26206 29492 26234 29532
rect 29549 29529 29561 29532
rect 29595 29560 29607 29563
rect 31386 29560 31392 29572
rect 29595 29532 31392 29560
rect 29595 29529 29607 29532
rect 29549 29523 29607 29529
rect 31386 29520 31392 29532
rect 31444 29520 31450 29572
rect 32674 29492 32680 29504
rect 26206 29464 32680 29492
rect 32674 29452 32680 29464
rect 32732 29452 32738 29504
rect 1104 29402 38824 29424
rect 1104 29350 10398 29402
rect 10450 29350 10462 29402
rect 10514 29350 10526 29402
rect 10578 29350 10590 29402
rect 10642 29350 10654 29402
rect 10706 29350 19846 29402
rect 19898 29350 19910 29402
rect 19962 29350 19974 29402
rect 20026 29350 20038 29402
rect 20090 29350 20102 29402
rect 20154 29350 29294 29402
rect 29346 29350 29358 29402
rect 29410 29350 29422 29402
rect 29474 29350 29486 29402
rect 29538 29350 29550 29402
rect 29602 29350 38824 29402
rect 1104 29328 38824 29350
rect 12526 29248 12532 29300
rect 12584 29288 12590 29300
rect 12805 29291 12863 29297
rect 12805 29288 12817 29291
rect 12584 29260 12817 29288
rect 12584 29248 12590 29260
rect 12805 29257 12817 29260
rect 12851 29257 12863 29291
rect 12805 29251 12863 29257
rect 24394 29248 24400 29300
rect 24452 29288 24458 29300
rect 24765 29291 24823 29297
rect 24765 29288 24777 29291
rect 24452 29260 24777 29288
rect 24452 29248 24458 29260
rect 24765 29257 24777 29260
rect 24811 29257 24823 29291
rect 24765 29251 24823 29257
rect 29089 29291 29147 29297
rect 29089 29257 29101 29291
rect 29135 29288 29147 29291
rect 29730 29288 29736 29300
rect 29135 29260 29736 29288
rect 29135 29257 29147 29260
rect 29089 29251 29147 29257
rect 29730 29248 29736 29260
rect 29788 29248 29794 29300
rect 31386 29288 31392 29300
rect 31347 29260 31392 29288
rect 31386 29248 31392 29260
rect 31444 29248 31450 29300
rect 32674 29288 32680 29300
rect 32635 29260 32680 29288
rect 32674 29248 32680 29260
rect 32732 29288 32738 29300
rect 34790 29288 34796 29300
rect 32732 29260 34796 29288
rect 32732 29248 32738 29260
rect 34790 29248 34796 29260
rect 34848 29248 34854 29300
rect 1673 29155 1731 29161
rect 1673 29121 1685 29155
rect 1719 29152 1731 29155
rect 11790 29152 11796 29164
rect 1719 29124 2084 29152
rect 11751 29124 11796 29152
rect 1719 29121 1731 29124
rect 1673 29115 1731 29121
rect 2056 29028 2084 29124
rect 11790 29112 11796 29124
rect 11848 29112 11854 29164
rect 12986 29152 12992 29164
rect 12947 29124 12992 29152
rect 12986 29112 12992 29124
rect 13044 29112 13050 29164
rect 15838 29152 15844 29164
rect 15799 29124 15844 29152
rect 15838 29112 15844 29124
rect 15896 29112 15902 29164
rect 17494 29152 17500 29164
rect 17455 29124 17500 29152
rect 17494 29112 17500 29124
rect 17552 29112 17558 29164
rect 24946 29152 24952 29164
rect 24907 29124 24952 29152
rect 24946 29112 24952 29124
rect 25004 29112 25010 29164
rect 28902 29152 28908 29164
rect 28863 29124 28908 29152
rect 28902 29112 28908 29124
rect 28960 29112 28966 29164
rect 31294 29152 31300 29164
rect 31255 29124 31300 29152
rect 31294 29112 31300 29124
rect 31352 29112 31358 29164
rect 32306 29112 32312 29164
rect 32364 29152 32370 29164
rect 32585 29155 32643 29161
rect 32585 29152 32597 29155
rect 32364 29124 32597 29152
rect 32364 29112 32370 29124
rect 32585 29121 32597 29124
rect 32631 29121 32643 29155
rect 32585 29115 32643 29121
rect 11517 29087 11575 29093
rect 11517 29053 11529 29087
rect 11563 29084 11575 29087
rect 12434 29084 12440 29096
rect 11563 29056 12440 29084
rect 11563 29053 11575 29056
rect 11517 29047 11575 29053
rect 12434 29044 12440 29056
rect 12492 29044 12498 29096
rect 13814 29044 13820 29096
rect 13872 29084 13878 29096
rect 15657 29087 15715 29093
rect 15657 29084 15669 29087
rect 13872 29056 15669 29084
rect 13872 29044 13878 29056
rect 15657 29053 15669 29056
rect 15703 29053 15715 29087
rect 17218 29084 17224 29096
rect 17179 29056 17224 29084
rect 15657 29047 15715 29053
rect 17218 29044 17224 29056
rect 17276 29044 17282 29096
rect 28721 29087 28779 29093
rect 28721 29053 28733 29087
rect 28767 29084 28779 29087
rect 31202 29084 31208 29096
rect 28767 29056 31208 29084
rect 28767 29053 28779 29056
rect 28721 29047 28779 29053
rect 31202 29044 31208 29056
rect 31260 29044 31266 29096
rect 1486 29016 1492 29028
rect 1447 28988 1492 29016
rect 1486 28976 1492 28988
rect 1544 28976 1550 29028
rect 2038 28976 2044 29028
rect 2096 29016 2102 29028
rect 2133 29019 2191 29025
rect 2133 29016 2145 29019
rect 2096 28988 2145 29016
rect 2096 28976 2102 28988
rect 2133 28985 2145 28988
rect 2179 28985 2191 29019
rect 2958 29016 2964 29028
rect 2919 28988 2964 29016
rect 2133 28979 2191 28985
rect 2958 28976 2964 28988
rect 3016 28976 3022 29028
rect 16025 29019 16083 29025
rect 16025 28985 16037 29019
rect 16071 29016 16083 29019
rect 16666 29016 16672 29028
rect 16071 28988 16672 29016
rect 16071 28985 16083 28988
rect 16025 28979 16083 28985
rect 16666 28976 16672 28988
rect 16724 28976 16730 29028
rect 18233 29019 18291 29025
rect 18233 28985 18245 29019
rect 18279 29016 18291 29019
rect 18322 29016 18328 29028
rect 18279 28988 18328 29016
rect 18279 28985 18291 28988
rect 18233 28979 18291 28985
rect 18322 28976 18328 28988
rect 18380 29016 18386 29028
rect 19426 29016 19432 29028
rect 18380 28988 19432 29016
rect 18380 28976 18386 28988
rect 19426 28976 19432 28988
rect 19484 28976 19490 29028
rect 13446 28948 13452 28960
rect 13407 28920 13452 28948
rect 13446 28908 13452 28920
rect 13504 28908 13510 28960
rect 1104 28858 38824 28880
rect 1104 28806 5674 28858
rect 5726 28806 5738 28858
rect 5790 28806 5802 28858
rect 5854 28806 5866 28858
rect 5918 28806 5930 28858
rect 5982 28806 15122 28858
rect 15174 28806 15186 28858
rect 15238 28806 15250 28858
rect 15302 28806 15314 28858
rect 15366 28806 15378 28858
rect 15430 28806 24570 28858
rect 24622 28806 24634 28858
rect 24686 28806 24698 28858
rect 24750 28806 24762 28858
rect 24814 28806 24826 28858
rect 24878 28806 34018 28858
rect 34070 28806 34082 28858
rect 34134 28806 34146 28858
rect 34198 28806 34210 28858
rect 34262 28806 34274 28858
rect 34326 28806 38824 28858
rect 1104 28784 38824 28806
rect 12529 28747 12587 28753
rect 12529 28713 12541 28747
rect 12575 28744 12587 28747
rect 12986 28744 12992 28756
rect 12575 28716 12992 28744
rect 12575 28713 12587 28716
rect 12529 28707 12587 28713
rect 12986 28704 12992 28716
rect 13044 28704 13050 28756
rect 16853 28747 16911 28753
rect 16853 28713 16865 28747
rect 16899 28744 16911 28747
rect 17494 28744 17500 28756
rect 16899 28716 17500 28744
rect 16899 28713 16911 28716
rect 16853 28707 16911 28713
rect 17494 28704 17500 28716
rect 17552 28704 17558 28756
rect 34790 28744 34796 28756
rect 34751 28716 34796 28744
rect 34790 28704 34796 28716
rect 34848 28704 34854 28756
rect 17218 28636 17224 28688
rect 17276 28676 17282 28688
rect 20073 28679 20131 28685
rect 20073 28676 20085 28679
rect 17276 28648 20085 28676
rect 17276 28636 17282 28648
rect 20073 28645 20085 28648
rect 20119 28645 20131 28679
rect 20073 28639 20131 28645
rect 12434 28608 12440 28620
rect 12360 28580 12440 28608
rect 9122 28540 9128 28552
rect 9083 28512 9128 28540
rect 9122 28500 9128 28512
rect 9180 28500 9186 28552
rect 12250 28540 12256 28552
rect 12211 28512 12256 28540
rect 12250 28500 12256 28512
rect 12308 28500 12314 28552
rect 12360 28549 12388 28580
rect 12434 28568 12440 28580
rect 12492 28608 12498 28620
rect 13446 28608 13452 28620
rect 12492 28580 13452 28608
rect 12492 28568 12498 28580
rect 13446 28568 13452 28580
rect 13504 28568 13510 28620
rect 13814 28568 13820 28620
rect 13872 28608 13878 28620
rect 14369 28611 14427 28617
rect 14369 28608 14381 28611
rect 13872 28580 14381 28608
rect 13872 28568 13878 28580
rect 14369 28577 14381 28580
rect 14415 28577 14427 28611
rect 14369 28571 14427 28577
rect 20993 28611 21051 28617
rect 20993 28577 21005 28611
rect 21039 28608 21051 28611
rect 21174 28608 21180 28620
rect 21039 28580 21180 28608
rect 21039 28577 21051 28580
rect 20993 28571 21051 28577
rect 21174 28568 21180 28580
rect 21232 28568 21238 28620
rect 12345 28543 12403 28549
rect 12345 28509 12357 28543
rect 12391 28509 12403 28543
rect 12345 28503 12403 28509
rect 13173 28543 13231 28549
rect 13173 28509 13185 28543
rect 13219 28540 13231 28543
rect 13998 28540 14004 28552
rect 13219 28512 14004 28540
rect 13219 28509 13231 28512
rect 13173 28503 13231 28509
rect 13998 28500 14004 28512
rect 14056 28500 14062 28552
rect 14090 28500 14096 28552
rect 14148 28540 14154 28552
rect 16666 28540 16672 28552
rect 14148 28512 14241 28540
rect 16627 28512 16672 28540
rect 14148 28500 14154 28512
rect 16666 28500 16672 28512
rect 16724 28500 16730 28552
rect 20257 28543 20315 28549
rect 20257 28509 20269 28543
rect 20303 28509 20315 28543
rect 20714 28540 20720 28552
rect 20675 28512 20720 28540
rect 20257 28503 20315 28509
rect 8386 28364 8392 28416
rect 8444 28404 8450 28416
rect 8941 28407 8999 28413
rect 8941 28404 8953 28407
rect 8444 28376 8953 28404
rect 8444 28364 8450 28376
rect 8941 28373 8953 28376
rect 8987 28373 8999 28407
rect 8941 28367 8999 28373
rect 12618 28364 12624 28416
rect 12676 28404 12682 28416
rect 12989 28407 13047 28413
rect 12989 28404 13001 28407
rect 12676 28376 13001 28404
rect 12676 28364 12682 28376
rect 12989 28373 13001 28376
rect 13035 28373 13047 28407
rect 14108 28404 14136 28500
rect 20272 28472 20300 28503
rect 20714 28500 20720 28512
rect 20772 28540 20778 28552
rect 22005 28543 22063 28549
rect 22005 28540 22017 28543
rect 20772 28512 22017 28540
rect 20772 28500 20778 28512
rect 22005 28509 22017 28512
rect 22051 28509 22063 28543
rect 22005 28503 22063 28509
rect 21266 28472 21272 28484
rect 20272 28444 21272 28472
rect 21266 28432 21272 28444
rect 21324 28432 21330 28484
rect 31294 28472 31300 28484
rect 22066 28444 31300 28472
rect 15473 28407 15531 28413
rect 15473 28404 15485 28407
rect 14108 28376 15485 28404
rect 12989 28367 13047 28373
rect 15473 28373 15485 28376
rect 15519 28404 15531 28407
rect 22066 28404 22094 28444
rect 31294 28432 31300 28444
rect 31352 28472 31358 28484
rect 31570 28472 31576 28484
rect 31352 28444 31576 28472
rect 31352 28432 31358 28444
rect 31570 28432 31576 28444
rect 31628 28432 31634 28484
rect 32306 28404 32312 28416
rect 15519 28376 22094 28404
rect 32267 28376 32312 28404
rect 15519 28373 15531 28376
rect 15473 28367 15531 28373
rect 32306 28364 32312 28376
rect 32364 28364 32370 28416
rect 1104 28314 38824 28336
rect 1104 28262 10398 28314
rect 10450 28262 10462 28314
rect 10514 28262 10526 28314
rect 10578 28262 10590 28314
rect 10642 28262 10654 28314
rect 10706 28262 19846 28314
rect 19898 28262 19910 28314
rect 19962 28262 19974 28314
rect 20026 28262 20038 28314
rect 20090 28262 20102 28314
rect 20154 28262 29294 28314
rect 29346 28262 29358 28314
rect 29410 28262 29422 28314
rect 29474 28262 29486 28314
rect 29538 28262 29550 28314
rect 29602 28262 38824 28314
rect 1104 28240 38824 28262
rect 24946 28200 24952 28212
rect 24907 28172 24952 28200
rect 24946 28160 24952 28172
rect 25004 28160 25010 28212
rect 28994 28160 29000 28212
rect 29052 28200 29058 28212
rect 29181 28203 29239 28209
rect 29181 28200 29193 28203
rect 29052 28172 29193 28200
rect 29052 28160 29058 28172
rect 29181 28169 29193 28172
rect 29227 28169 29239 28203
rect 29181 28163 29239 28169
rect 19061 28135 19119 28141
rect 19061 28101 19073 28135
rect 19107 28132 19119 28135
rect 19613 28135 19671 28141
rect 19613 28132 19625 28135
rect 19107 28104 19625 28132
rect 19107 28101 19119 28104
rect 19061 28095 19119 28101
rect 19613 28101 19625 28104
rect 19659 28132 19671 28135
rect 32306 28132 32312 28144
rect 19659 28104 32312 28132
rect 19659 28101 19671 28104
rect 19613 28095 19671 28101
rect 32306 28092 32312 28104
rect 32364 28092 32370 28144
rect 1673 28067 1731 28073
rect 1673 28033 1685 28067
rect 1719 28064 1731 28067
rect 8386 28064 8392 28076
rect 1719 28036 2268 28064
rect 8347 28036 8392 28064
rect 1719 28033 1731 28036
rect 1673 28027 1731 28033
rect 1486 27860 1492 27872
rect 1447 27832 1492 27860
rect 1486 27820 1492 27832
rect 1544 27820 1550 27872
rect 2240 27869 2268 28036
rect 8386 28024 8392 28036
rect 8444 28024 8450 28076
rect 20990 28064 20996 28076
rect 20951 28036 20996 28064
rect 20990 28024 20996 28036
rect 21048 28024 21054 28076
rect 21266 28064 21272 28076
rect 21227 28036 21272 28064
rect 21266 28024 21272 28036
rect 21324 28064 21330 28076
rect 21324 28036 22094 28064
rect 21324 28024 21330 28036
rect 8110 27996 8116 28008
rect 8071 27968 8116 27996
rect 8110 27956 8116 27968
rect 8168 27956 8174 28008
rect 22066 27996 22094 28036
rect 24118 28024 24124 28076
rect 24176 28064 24182 28076
rect 24765 28067 24823 28073
rect 24765 28064 24777 28067
rect 24176 28036 24777 28064
rect 24176 28024 24182 28036
rect 24765 28033 24777 28036
rect 24811 28033 24823 28067
rect 28166 28064 28172 28076
rect 28127 28036 28172 28064
rect 24765 28027 24823 28033
rect 28166 28024 28172 28036
rect 28224 28024 28230 28076
rect 28442 28064 28448 28076
rect 28403 28036 28448 28064
rect 28442 28024 28448 28036
rect 28500 28024 28506 28076
rect 31846 28024 31852 28076
rect 31904 28064 31910 28076
rect 34333 28067 34391 28073
rect 34333 28064 34345 28067
rect 31904 28036 34345 28064
rect 31904 28024 31910 28036
rect 34333 28033 34345 28036
rect 34379 28064 34391 28067
rect 35161 28067 35219 28073
rect 35161 28064 35173 28067
rect 34379 28036 35173 28064
rect 34379 28033 34391 28036
rect 34333 28027 34391 28033
rect 35161 28033 35173 28036
rect 35207 28033 35219 28067
rect 35161 28027 35219 28033
rect 35345 28067 35403 28073
rect 35345 28033 35357 28067
rect 35391 28064 35403 28067
rect 35805 28067 35863 28073
rect 35805 28064 35817 28067
rect 35391 28036 35817 28064
rect 35391 28033 35403 28036
rect 35345 28027 35403 28033
rect 35805 28033 35817 28036
rect 35851 28033 35863 28067
rect 35805 28027 35863 28033
rect 23474 27996 23480 28008
rect 22066 27968 23480 27996
rect 23474 27956 23480 27968
rect 23532 27956 23538 28008
rect 24581 27999 24639 28005
rect 24581 27996 24593 27999
rect 24320 27968 24593 27996
rect 12250 27888 12256 27940
rect 12308 27928 12314 27940
rect 12897 27931 12955 27937
rect 12897 27928 12909 27931
rect 12308 27900 12909 27928
rect 12308 27888 12314 27900
rect 12897 27897 12909 27900
rect 12943 27928 12955 27931
rect 19334 27928 19340 27940
rect 12943 27900 19340 27928
rect 12943 27897 12955 27900
rect 12897 27891 12955 27897
rect 19334 27888 19340 27900
rect 19392 27888 19398 27940
rect 19426 27888 19432 27940
rect 19484 27928 19490 27940
rect 20257 27931 20315 27937
rect 20257 27928 20269 27931
rect 19484 27900 20269 27928
rect 19484 27888 19490 27900
rect 20257 27897 20269 27900
rect 20303 27897 20315 27931
rect 20257 27891 20315 27897
rect 24320 27872 24348 27968
rect 24581 27965 24593 27968
rect 24627 27965 24639 27999
rect 24581 27959 24639 27965
rect 31202 27956 31208 28008
rect 31260 27996 31266 28008
rect 34149 27999 34207 28005
rect 34149 27996 34161 27999
rect 31260 27968 34161 27996
rect 31260 27956 31266 27968
rect 34149 27965 34161 27968
rect 34195 27965 34207 27999
rect 34149 27959 34207 27965
rect 34514 27956 34520 28008
rect 34572 27996 34578 28008
rect 34790 27996 34796 28008
rect 34572 27968 34796 27996
rect 34572 27956 34578 27968
rect 34790 27956 34796 27968
rect 34848 27996 34854 28008
rect 34977 27999 35035 28005
rect 34977 27996 34989 27999
rect 34848 27968 34989 27996
rect 34848 27956 34854 27968
rect 34977 27965 34989 27968
rect 35023 27965 35035 27999
rect 34977 27959 35035 27965
rect 2225 27863 2283 27869
rect 2225 27829 2237 27863
rect 2271 27860 2283 27863
rect 2314 27860 2320 27872
rect 2271 27832 2320 27860
rect 2271 27829 2283 27832
rect 2225 27823 2283 27829
rect 2314 27820 2320 27832
rect 2372 27820 2378 27872
rect 8386 27820 8392 27872
rect 8444 27860 8450 27872
rect 9125 27863 9183 27869
rect 9125 27860 9137 27863
rect 8444 27832 9137 27860
rect 8444 27820 8450 27832
rect 9125 27829 9137 27832
rect 9171 27829 9183 27863
rect 13446 27860 13452 27872
rect 13407 27832 13452 27860
rect 9125 27823 9183 27829
rect 13446 27820 13452 27832
rect 13504 27820 13510 27872
rect 19702 27860 19708 27872
rect 19663 27832 19708 27860
rect 19702 27820 19708 27832
rect 19760 27820 19766 27872
rect 24121 27863 24179 27869
rect 24121 27829 24133 27863
rect 24167 27860 24179 27863
rect 24302 27860 24308 27872
rect 24167 27832 24308 27860
rect 24167 27829 24179 27832
rect 24121 27823 24179 27829
rect 24302 27820 24308 27832
rect 24360 27820 24366 27872
rect 34517 27863 34575 27869
rect 34517 27829 34529 27863
rect 34563 27860 34575 27863
rect 34974 27860 34980 27872
rect 34563 27832 34980 27860
rect 34563 27829 34575 27832
rect 34517 27823 34575 27829
rect 34974 27820 34980 27832
rect 35032 27820 35038 27872
rect 35894 27820 35900 27872
rect 35952 27860 35958 27872
rect 35989 27863 36047 27869
rect 35989 27860 36001 27863
rect 35952 27832 36001 27860
rect 35952 27820 35958 27832
rect 35989 27829 36001 27832
rect 36035 27829 36047 27863
rect 35989 27823 36047 27829
rect 1104 27770 38824 27792
rect 1104 27718 5674 27770
rect 5726 27718 5738 27770
rect 5790 27718 5802 27770
rect 5854 27718 5866 27770
rect 5918 27718 5930 27770
rect 5982 27718 15122 27770
rect 15174 27718 15186 27770
rect 15238 27718 15250 27770
rect 15302 27718 15314 27770
rect 15366 27718 15378 27770
rect 15430 27718 24570 27770
rect 24622 27718 24634 27770
rect 24686 27718 24698 27770
rect 24750 27718 24762 27770
rect 24814 27718 24826 27770
rect 24878 27718 34018 27770
rect 34070 27718 34082 27770
rect 34134 27718 34146 27770
rect 34198 27718 34210 27770
rect 34262 27718 34274 27770
rect 34326 27718 38824 27770
rect 1104 27696 38824 27718
rect 8941 27659 8999 27665
rect 4172 27628 5672 27656
rect 3050 27548 3056 27600
rect 3108 27588 3114 27600
rect 4172 27588 4200 27628
rect 3108 27560 4200 27588
rect 5644 27588 5672 27628
rect 8941 27625 8953 27659
rect 8987 27656 8999 27659
rect 9122 27656 9128 27668
rect 8987 27628 9128 27656
rect 8987 27625 8999 27628
rect 8941 27619 8999 27625
rect 9122 27616 9128 27628
rect 9180 27616 9186 27668
rect 20990 27656 20996 27668
rect 20951 27628 20996 27656
rect 20990 27616 20996 27628
rect 21048 27616 21054 27668
rect 6089 27591 6147 27597
rect 6089 27588 6101 27591
rect 5644 27560 6101 27588
rect 3108 27548 3114 27560
rect 6089 27557 6101 27560
rect 6135 27588 6147 27591
rect 8386 27588 8392 27600
rect 6135 27560 8392 27588
rect 6135 27557 6147 27560
rect 6089 27551 6147 27557
rect 8386 27548 8392 27560
rect 8444 27548 8450 27600
rect 23474 27548 23480 27600
rect 23532 27588 23538 27600
rect 24765 27591 24823 27597
rect 24765 27588 24777 27591
rect 23532 27560 24777 27588
rect 23532 27548 23538 27560
rect 24765 27557 24777 27560
rect 24811 27557 24823 27591
rect 24765 27551 24823 27557
rect 31386 27548 31392 27600
rect 31444 27588 31450 27600
rect 31665 27591 31723 27597
rect 31665 27588 31677 27591
rect 31444 27560 31677 27588
rect 31444 27548 31450 27560
rect 31665 27557 31677 27560
rect 31711 27557 31723 27591
rect 31665 27551 31723 27557
rect 6748 27492 9168 27520
rect 6748 27464 6776 27492
rect 2685 27455 2743 27461
rect 2685 27421 2697 27455
rect 2731 27452 2743 27455
rect 2866 27452 2872 27464
rect 2731 27424 2872 27452
rect 2731 27421 2743 27424
rect 2685 27415 2743 27421
rect 2866 27412 2872 27424
rect 2924 27412 2930 27464
rect 5074 27452 5080 27464
rect 5035 27424 5080 27452
rect 5074 27412 5080 27424
rect 5132 27412 5138 27464
rect 5353 27455 5411 27461
rect 5353 27421 5365 27455
rect 5399 27452 5411 27455
rect 5534 27452 5540 27464
rect 5399 27424 5540 27452
rect 5399 27421 5411 27424
rect 5353 27415 5411 27421
rect 5534 27412 5540 27424
rect 5592 27412 5598 27464
rect 6730 27452 6736 27464
rect 6691 27424 6736 27452
rect 6730 27412 6736 27424
rect 6788 27412 6794 27464
rect 6914 27412 6920 27464
rect 6972 27452 6978 27464
rect 9140 27461 9168 27492
rect 24118 27480 24124 27532
rect 24176 27520 24182 27532
rect 24176 27492 28672 27520
rect 24176 27480 24182 27492
rect 9125 27455 9183 27461
rect 6972 27424 7017 27452
rect 6972 27412 6978 27424
rect 9125 27421 9137 27455
rect 9171 27452 9183 27455
rect 9214 27452 9220 27464
rect 9171 27424 9220 27452
rect 9171 27421 9183 27424
rect 9125 27415 9183 27421
rect 9214 27412 9220 27424
rect 9272 27412 9278 27464
rect 9309 27455 9367 27461
rect 9309 27421 9321 27455
rect 9355 27452 9367 27455
rect 19981 27455 20039 27461
rect 19981 27452 19993 27455
rect 9355 27424 9904 27452
rect 9355 27421 9367 27424
rect 9309 27415 9367 27421
rect 5718 27344 5724 27396
rect 5776 27384 5782 27396
rect 7374 27384 7380 27396
rect 5776 27356 7380 27384
rect 5776 27344 5782 27356
rect 7374 27344 7380 27356
rect 7432 27384 7438 27396
rect 8110 27384 8116 27396
rect 7432 27356 8116 27384
rect 7432 27344 7438 27356
rect 8110 27344 8116 27356
rect 8168 27344 8174 27396
rect 9876 27328 9904 27424
rect 19444 27424 19993 27452
rect 2869 27319 2927 27325
rect 2869 27285 2881 27319
rect 2915 27316 2927 27319
rect 3234 27316 3240 27328
rect 2915 27288 3240 27316
rect 2915 27285 2927 27288
rect 2869 27279 2927 27285
rect 3234 27276 3240 27288
rect 3292 27276 3298 27328
rect 6546 27316 6552 27328
rect 6507 27288 6552 27316
rect 6546 27276 6552 27288
rect 6604 27276 6610 27328
rect 9858 27316 9864 27328
rect 9819 27288 9864 27316
rect 9858 27276 9864 27288
rect 9916 27276 9922 27328
rect 19334 27276 19340 27328
rect 19392 27316 19398 27328
rect 19444 27325 19472 27424
rect 19981 27421 19993 27424
rect 20027 27421 20039 27455
rect 19981 27415 20039 27421
rect 20165 27455 20223 27461
rect 20165 27421 20177 27455
rect 20211 27421 20223 27455
rect 20165 27415 20223 27421
rect 20349 27455 20407 27461
rect 20349 27421 20361 27455
rect 20395 27452 20407 27455
rect 20809 27455 20867 27461
rect 20809 27452 20821 27455
rect 20395 27424 20821 27452
rect 20395 27421 20407 27424
rect 20349 27415 20407 27421
rect 20809 27421 20821 27424
rect 20855 27421 20867 27455
rect 28534 27452 28540 27464
rect 28495 27424 28540 27452
rect 20809 27415 20867 27421
rect 20180 27384 20208 27415
rect 28534 27412 28540 27424
rect 28592 27412 28598 27464
rect 28644 27461 28672 27492
rect 28629 27455 28687 27461
rect 28629 27421 28641 27455
rect 28675 27421 28687 27455
rect 34974 27452 34980 27464
rect 34935 27424 34980 27452
rect 28629 27415 28687 27421
rect 34974 27412 34980 27424
rect 35032 27412 35038 27464
rect 35618 27452 35624 27464
rect 35579 27424 35624 27452
rect 35618 27412 35624 27424
rect 35676 27412 35682 27464
rect 35897 27455 35955 27461
rect 35897 27421 35909 27455
rect 35943 27421 35955 27455
rect 36722 27452 36728 27464
rect 36683 27424 36728 27452
rect 35897 27415 35955 27421
rect 20714 27384 20720 27396
rect 20180 27356 20720 27384
rect 20714 27344 20720 27356
rect 20772 27344 20778 27396
rect 24946 27384 24952 27396
rect 24907 27356 24952 27384
rect 24946 27344 24952 27356
rect 25004 27344 25010 27396
rect 35912 27384 35940 27415
rect 36722 27412 36728 27424
rect 36780 27412 36786 27464
rect 35866 27356 35940 27384
rect 19429 27319 19487 27325
rect 19429 27316 19441 27319
rect 19392 27288 19441 27316
rect 19392 27276 19398 27288
rect 19429 27285 19441 27288
rect 19475 27285 19487 27319
rect 19429 27279 19487 27285
rect 28718 27276 28724 27328
rect 28776 27316 28782 27328
rect 28813 27319 28871 27325
rect 28813 27316 28825 27319
rect 28776 27288 28825 27316
rect 28776 27276 28782 27288
rect 28813 27285 28825 27288
rect 28859 27285 28871 27319
rect 28813 27279 28871 27285
rect 35161 27319 35219 27325
rect 35161 27285 35173 27319
rect 35207 27316 35219 27319
rect 35866 27316 35894 27356
rect 35207 27288 35894 27316
rect 35207 27285 35219 27288
rect 35161 27279 35219 27285
rect 1104 27226 38824 27248
rect 1104 27174 10398 27226
rect 10450 27174 10462 27226
rect 10514 27174 10526 27226
rect 10578 27174 10590 27226
rect 10642 27174 10654 27226
rect 10706 27174 19846 27226
rect 19898 27174 19910 27226
rect 19962 27174 19974 27226
rect 20026 27174 20038 27226
rect 20090 27174 20102 27226
rect 20154 27174 29294 27226
rect 29346 27174 29358 27226
rect 29410 27174 29422 27226
rect 29474 27174 29486 27226
rect 29538 27174 29550 27226
rect 29602 27174 38824 27226
rect 1104 27152 38824 27174
rect 2501 27115 2559 27121
rect 2501 27081 2513 27115
rect 2547 27112 2559 27115
rect 3050 27112 3056 27124
rect 2547 27084 3056 27112
rect 2547 27081 2559 27084
rect 2501 27075 2559 27081
rect 3050 27072 3056 27084
rect 3108 27072 3114 27124
rect 5534 27112 5540 27124
rect 5495 27084 5540 27112
rect 5534 27072 5540 27084
rect 5592 27072 5598 27124
rect 24118 27112 24124 27124
rect 24079 27084 24124 27112
rect 24118 27072 24124 27084
rect 24176 27072 24182 27124
rect 28442 27072 28448 27124
rect 28500 27112 28506 27124
rect 28537 27115 28595 27121
rect 28537 27112 28549 27115
rect 28500 27084 28549 27112
rect 28500 27072 28506 27084
rect 28537 27081 28549 27084
rect 28583 27081 28595 27115
rect 28537 27075 28595 27081
rect 3970 27004 3976 27056
rect 4028 27044 4034 27056
rect 6730 27044 6736 27056
rect 4028 27016 6736 27044
rect 4028 27004 4034 27016
rect 6730 27004 6736 27016
rect 6788 27004 6794 27056
rect 3234 26976 3240 26988
rect 3195 26948 3240 26976
rect 3234 26936 3240 26948
rect 3292 26936 3298 26988
rect 3513 26979 3571 26985
rect 3513 26945 3525 26979
rect 3559 26976 3571 26979
rect 5074 26976 5080 26988
rect 3559 26948 5080 26976
rect 3559 26945 3571 26948
rect 3513 26939 3571 26945
rect 5074 26936 5080 26948
rect 5132 26976 5138 26988
rect 5626 26976 5632 26988
rect 5132 26948 5632 26976
rect 5132 26936 5138 26948
rect 5626 26936 5632 26948
rect 5684 26936 5690 26988
rect 5721 26979 5779 26985
rect 5721 26945 5733 26979
rect 5767 26976 5779 26979
rect 6546 26976 6552 26988
rect 5767 26948 6552 26976
rect 5767 26945 5779 26948
rect 5721 26939 5779 26945
rect 6546 26936 6552 26948
rect 6604 26936 6610 26988
rect 7834 26976 7840 26988
rect 7795 26948 7840 26976
rect 7834 26936 7840 26948
rect 7892 26936 7898 26988
rect 23566 26936 23572 26988
rect 23624 26976 23630 26988
rect 23937 26979 23995 26985
rect 23937 26976 23949 26979
rect 23624 26948 23949 26976
rect 23624 26936 23630 26948
rect 23937 26945 23949 26948
rect 23983 26945 23995 26979
rect 28718 26976 28724 26988
rect 28679 26948 28724 26976
rect 23937 26939 23995 26945
rect 28718 26936 28724 26948
rect 28776 26936 28782 26988
rect 30650 26936 30656 26988
rect 30708 26976 30714 26988
rect 31294 26976 31300 26988
rect 30708 26948 31300 26976
rect 30708 26936 30714 26948
rect 31294 26936 31300 26948
rect 31352 26936 31358 26988
rect 31389 26979 31447 26985
rect 31389 26945 31401 26979
rect 31435 26976 31447 26979
rect 31846 26976 31852 26988
rect 31435 26948 31852 26976
rect 31435 26945 31447 26948
rect 31389 26939 31447 26945
rect 31846 26936 31852 26948
rect 31904 26936 31910 26988
rect 32950 26976 32956 26988
rect 32911 26948 32956 26976
rect 32950 26936 32956 26948
rect 33008 26936 33014 26988
rect 35894 26936 35900 26988
rect 35952 26976 35958 26988
rect 36722 26976 36728 26988
rect 35952 26948 35997 26976
rect 36683 26948 36728 26976
rect 35952 26936 35958 26948
rect 36722 26936 36728 26948
rect 36780 26936 36786 26988
rect 33229 26911 33287 26917
rect 33229 26877 33241 26911
rect 33275 26908 33287 26911
rect 33778 26908 33784 26920
rect 33275 26880 33784 26908
rect 33275 26877 33287 26880
rect 33229 26871 33287 26877
rect 33778 26868 33784 26880
rect 33836 26908 33842 26920
rect 35618 26908 35624 26920
rect 33836 26880 35624 26908
rect 33836 26868 33842 26880
rect 35618 26868 35624 26880
rect 35676 26868 35682 26920
rect 7650 26772 7656 26784
rect 7611 26744 7656 26772
rect 7650 26732 7656 26744
rect 7708 26732 7714 26784
rect 9858 26732 9864 26784
rect 9916 26772 9922 26784
rect 14918 26772 14924 26784
rect 9916 26744 14924 26772
rect 9916 26732 9922 26744
rect 14918 26732 14924 26744
rect 14976 26772 14982 26784
rect 15473 26775 15531 26781
rect 15473 26772 15485 26775
rect 14976 26744 15485 26772
rect 14976 26732 14982 26744
rect 15473 26741 15485 26744
rect 15519 26772 15531 26775
rect 19518 26772 19524 26784
rect 15519 26744 19524 26772
rect 15519 26741 15531 26744
rect 15473 26735 15531 26741
rect 19518 26732 19524 26744
rect 19576 26732 19582 26784
rect 20533 26775 20591 26781
rect 20533 26741 20545 26775
rect 20579 26772 20591 26775
rect 20714 26772 20720 26784
rect 20579 26744 20720 26772
rect 20579 26741 20591 26744
rect 20533 26735 20591 26741
rect 20714 26732 20720 26744
rect 20772 26772 20778 26784
rect 21266 26772 21272 26784
rect 20772 26744 21272 26772
rect 20772 26732 20778 26744
rect 21266 26732 21272 26744
rect 21324 26732 21330 26784
rect 31573 26775 31631 26781
rect 31573 26741 31585 26775
rect 31619 26772 31631 26775
rect 31662 26772 31668 26784
rect 31619 26744 31668 26772
rect 31619 26741 31631 26744
rect 31573 26735 31631 26741
rect 31662 26732 31668 26744
rect 31720 26732 31726 26784
rect 32207 26775 32265 26781
rect 32207 26741 32219 26775
rect 32253 26772 32265 26775
rect 33870 26772 33876 26784
rect 32253 26744 33876 26772
rect 32253 26741 32265 26744
rect 32207 26735 32265 26741
rect 33870 26732 33876 26744
rect 33928 26732 33934 26784
rect 1104 26682 38824 26704
rect 1104 26630 5674 26682
rect 5726 26630 5738 26682
rect 5790 26630 5802 26682
rect 5854 26630 5866 26682
rect 5918 26630 5930 26682
rect 5982 26630 15122 26682
rect 15174 26630 15186 26682
rect 15238 26630 15250 26682
rect 15302 26630 15314 26682
rect 15366 26630 15378 26682
rect 15430 26630 24570 26682
rect 24622 26630 24634 26682
rect 24686 26630 24698 26682
rect 24750 26630 24762 26682
rect 24814 26630 24826 26682
rect 24878 26630 34018 26682
rect 34070 26630 34082 26682
rect 34134 26630 34146 26682
rect 34198 26630 34210 26682
rect 34262 26630 34274 26682
rect 34326 26630 38824 26682
rect 1104 26608 38824 26630
rect 2866 26568 2872 26580
rect 2827 26540 2872 26568
rect 2866 26528 2872 26540
rect 2924 26528 2930 26580
rect 8386 26568 8392 26580
rect 8347 26540 8392 26568
rect 8386 26528 8392 26540
rect 8444 26528 8450 26580
rect 13998 26528 14004 26580
rect 14056 26568 14062 26580
rect 19245 26571 19303 26577
rect 19245 26568 19257 26571
rect 14056 26540 19257 26568
rect 14056 26528 14062 26540
rect 19245 26537 19257 26540
rect 19291 26537 19303 26571
rect 19245 26531 19303 26537
rect 31849 26571 31907 26577
rect 31849 26537 31861 26571
rect 31895 26568 31907 26571
rect 32950 26568 32956 26580
rect 31895 26540 32956 26568
rect 31895 26537 31907 26540
rect 31849 26531 31907 26537
rect 32950 26528 32956 26540
rect 33008 26528 33014 26580
rect 2225 26503 2283 26509
rect 2225 26469 2237 26503
rect 2271 26469 2283 26503
rect 2225 26463 2283 26469
rect 1673 26367 1731 26373
rect 1673 26333 1685 26367
rect 1719 26364 1731 26367
rect 2240 26364 2268 26463
rect 7374 26432 7380 26444
rect 7335 26404 7380 26432
rect 7374 26392 7380 26404
rect 7432 26392 7438 26444
rect 14918 26432 14924 26444
rect 14879 26404 14924 26432
rect 14918 26392 14924 26404
rect 14976 26392 14982 26444
rect 2406 26364 2412 26376
rect 1719 26336 2268 26364
rect 2367 26336 2412 26364
rect 1719 26333 1731 26336
rect 1673 26327 1731 26333
rect 2406 26324 2412 26336
rect 2464 26364 2470 26376
rect 2958 26364 2964 26376
rect 2464 26336 2964 26364
rect 2464 26324 2470 26336
rect 2958 26324 2964 26336
rect 3016 26324 3022 26376
rect 3053 26367 3111 26373
rect 3053 26333 3065 26367
rect 3099 26333 3111 26367
rect 3053 26327 3111 26333
rect 3068 26296 3096 26327
rect 3142 26324 3148 26376
rect 3200 26364 3206 26376
rect 3789 26367 3847 26373
rect 3789 26364 3801 26367
rect 3200 26336 3801 26364
rect 3200 26324 3206 26336
rect 3789 26333 3801 26336
rect 3835 26364 3847 26367
rect 3878 26364 3884 26376
rect 3835 26336 3884 26364
rect 3835 26333 3847 26336
rect 3789 26327 3847 26333
rect 3878 26324 3884 26336
rect 3936 26324 3942 26376
rect 7650 26364 7656 26376
rect 7611 26336 7656 26364
rect 7650 26324 7656 26336
rect 7708 26324 7714 26376
rect 12342 26364 12348 26376
rect 12303 26336 12348 26364
rect 12342 26324 12348 26336
rect 12400 26324 12406 26376
rect 15010 26324 15016 26376
rect 15068 26364 15074 26376
rect 15105 26367 15163 26373
rect 15105 26364 15117 26367
rect 15068 26336 15117 26364
rect 15068 26324 15074 26336
rect 15105 26333 15117 26336
rect 15151 26333 15163 26367
rect 15105 26327 15163 26333
rect 15562 26324 15568 26376
rect 15620 26364 15626 26376
rect 15749 26367 15807 26373
rect 15749 26364 15761 26367
rect 15620 26336 15761 26364
rect 15620 26324 15626 26336
rect 15749 26333 15761 26336
rect 15795 26333 15807 26367
rect 16022 26364 16028 26376
rect 15983 26336 16028 26364
rect 15749 26327 15807 26333
rect 16022 26324 16028 26336
rect 16080 26324 16086 26376
rect 19429 26367 19487 26373
rect 19429 26333 19441 26367
rect 19475 26364 19487 26367
rect 21818 26364 21824 26376
rect 19475 26336 21824 26364
rect 19475 26333 19487 26336
rect 19429 26327 19487 26333
rect 21818 26324 21824 26336
rect 21876 26324 21882 26376
rect 24854 26364 24860 26376
rect 24815 26336 24860 26364
rect 24854 26324 24860 26336
rect 24912 26324 24918 26376
rect 31662 26364 31668 26376
rect 31623 26336 31668 26364
rect 31662 26324 31668 26336
rect 31720 26324 31726 26376
rect 3970 26296 3976 26308
rect 3068 26268 3976 26296
rect 3970 26256 3976 26268
rect 4028 26256 4034 26308
rect 19610 26296 19616 26308
rect 19571 26268 19616 26296
rect 19610 26256 19616 26268
rect 19668 26256 19674 26308
rect 1486 26228 1492 26240
rect 1447 26200 1492 26228
rect 1486 26188 1492 26200
rect 1544 26188 1550 26240
rect 12158 26228 12164 26240
rect 12119 26200 12164 26228
rect 12158 26188 12164 26200
rect 12216 26188 12222 26240
rect 15289 26231 15347 26237
rect 15289 26197 15301 26231
rect 15335 26228 15347 26231
rect 15746 26228 15752 26240
rect 15335 26200 15752 26228
rect 15335 26197 15347 26200
rect 15289 26191 15347 26197
rect 15746 26188 15752 26200
rect 15804 26188 15810 26240
rect 16761 26231 16819 26237
rect 16761 26197 16773 26231
rect 16807 26228 16819 26231
rect 17034 26228 17040 26240
rect 16807 26200 17040 26228
rect 16807 26197 16819 26200
rect 16761 26191 16819 26197
rect 17034 26188 17040 26200
rect 17092 26188 17098 26240
rect 25038 26228 25044 26240
rect 24999 26200 25044 26228
rect 25038 26188 25044 26200
rect 25096 26188 25102 26240
rect 1104 26138 38824 26160
rect 1104 26086 10398 26138
rect 10450 26086 10462 26138
rect 10514 26086 10526 26138
rect 10578 26086 10590 26138
rect 10642 26086 10654 26138
rect 10706 26086 19846 26138
rect 19898 26086 19910 26138
rect 19962 26086 19974 26138
rect 20026 26086 20038 26138
rect 20090 26086 20102 26138
rect 20154 26086 29294 26138
rect 29346 26086 29358 26138
rect 29410 26086 29422 26138
rect 29474 26086 29486 26138
rect 29538 26086 29550 26138
rect 29602 26086 38824 26138
rect 1104 26064 38824 26086
rect 7745 26027 7803 26033
rect 7745 25993 7757 26027
rect 7791 26024 7803 26027
rect 7834 26024 7840 26036
rect 7791 25996 7840 26024
rect 7791 25993 7803 25996
rect 7745 25987 7803 25993
rect 7834 25984 7840 25996
rect 7892 25984 7898 26036
rect 15933 26027 15991 26033
rect 15933 25993 15945 26027
rect 15979 26024 15991 26027
rect 16022 26024 16028 26036
rect 15979 25996 16028 26024
rect 15979 25993 15991 25996
rect 15933 25987 15991 25993
rect 16022 25984 16028 25996
rect 16080 25984 16086 26036
rect 24854 25984 24860 26036
rect 24912 26024 24918 26036
rect 25777 26027 25835 26033
rect 25777 26024 25789 26027
rect 24912 25996 25789 26024
rect 24912 25984 24918 25996
rect 25777 25993 25789 25996
rect 25823 25993 25835 26027
rect 25777 25987 25835 25993
rect 7561 25891 7619 25897
rect 7561 25857 7573 25891
rect 7607 25888 7619 25891
rect 9214 25888 9220 25900
rect 7607 25860 9220 25888
rect 7607 25857 7619 25860
rect 7561 25851 7619 25857
rect 9214 25848 9220 25860
rect 9272 25848 9278 25900
rect 11977 25891 12035 25897
rect 11977 25857 11989 25891
rect 12023 25888 12035 25891
rect 12158 25888 12164 25900
rect 12023 25860 12164 25888
rect 12023 25857 12035 25860
rect 11977 25851 12035 25857
rect 12158 25848 12164 25860
rect 12216 25848 12222 25900
rect 15746 25888 15752 25900
rect 15707 25860 15752 25888
rect 15746 25848 15752 25860
rect 15804 25848 15810 25900
rect 25038 25888 25044 25900
rect 24999 25860 25044 25888
rect 25038 25848 25044 25860
rect 25096 25848 25102 25900
rect 25958 25888 25964 25900
rect 25919 25860 25964 25888
rect 25958 25848 25964 25860
rect 26016 25848 26022 25900
rect 28442 25888 28448 25900
rect 28403 25860 28448 25888
rect 28442 25848 28448 25860
rect 28500 25848 28506 25900
rect 7374 25820 7380 25832
rect 7335 25792 7380 25820
rect 7374 25780 7380 25792
rect 7432 25780 7438 25832
rect 11698 25820 11704 25832
rect 11659 25792 11704 25820
rect 11698 25780 11704 25792
rect 11756 25780 11762 25832
rect 25314 25780 25320 25832
rect 25372 25820 25378 25832
rect 26145 25823 26203 25829
rect 25372 25792 26096 25820
rect 25372 25780 25378 25792
rect 2406 25644 2412 25696
rect 2464 25684 2470 25696
rect 2593 25687 2651 25693
rect 2593 25684 2605 25687
rect 2464 25656 2605 25684
rect 2464 25644 2470 25656
rect 2593 25653 2605 25656
rect 2639 25684 2651 25687
rect 4338 25684 4344 25696
rect 2639 25656 4344 25684
rect 2639 25653 2651 25656
rect 2593 25647 2651 25653
rect 4338 25644 4344 25656
rect 4396 25644 4402 25696
rect 12434 25644 12440 25696
rect 12492 25684 12498 25696
rect 12713 25687 12771 25693
rect 12713 25684 12725 25687
rect 12492 25656 12725 25684
rect 12492 25644 12498 25656
rect 12713 25653 12725 25656
rect 12759 25684 12771 25687
rect 17034 25684 17040 25696
rect 12759 25656 17040 25684
rect 12759 25653 12771 25656
rect 12713 25647 12771 25653
rect 17034 25644 17040 25656
rect 17092 25644 17098 25696
rect 22830 25644 22836 25696
rect 22888 25684 22894 25696
rect 24305 25687 24363 25693
rect 24305 25684 24317 25687
rect 22888 25656 24317 25684
rect 22888 25644 22894 25656
rect 24305 25653 24317 25656
rect 24351 25653 24363 25687
rect 26068 25684 26096 25792
rect 26145 25789 26157 25823
rect 26191 25789 26203 25823
rect 27065 25823 27123 25829
rect 27065 25820 27077 25823
rect 26145 25783 26203 25789
rect 26804 25792 27077 25820
rect 26160 25752 26188 25783
rect 26804 25752 26832 25792
rect 27065 25789 27077 25792
rect 27111 25820 27123 25823
rect 30650 25820 30656 25832
rect 27111 25792 30656 25820
rect 27111 25789 27123 25792
rect 27065 25783 27123 25789
rect 30650 25780 30656 25792
rect 30708 25780 30714 25832
rect 27706 25752 27712 25764
rect 26160 25724 26832 25752
rect 26896 25724 27712 25752
rect 26896 25684 26924 25724
rect 27706 25712 27712 25724
rect 27764 25712 27770 25764
rect 26068 25656 26924 25684
rect 24305 25647 24363 25653
rect 27798 25644 27804 25696
rect 27856 25684 27862 25696
rect 28261 25687 28319 25693
rect 28261 25684 28273 25687
rect 27856 25656 28273 25684
rect 27856 25644 27862 25656
rect 28261 25653 28273 25656
rect 28307 25653 28319 25687
rect 28261 25647 28319 25653
rect 1104 25594 38824 25616
rect 1104 25542 5674 25594
rect 5726 25542 5738 25594
rect 5790 25542 5802 25594
rect 5854 25542 5866 25594
rect 5918 25542 5930 25594
rect 5982 25542 15122 25594
rect 15174 25542 15186 25594
rect 15238 25542 15250 25594
rect 15302 25542 15314 25594
rect 15366 25542 15378 25594
rect 15430 25542 24570 25594
rect 24622 25542 24634 25594
rect 24686 25542 24698 25594
rect 24750 25542 24762 25594
rect 24814 25542 24826 25594
rect 24878 25542 34018 25594
rect 34070 25542 34082 25594
rect 34134 25542 34146 25594
rect 34198 25542 34210 25594
rect 34262 25542 34274 25594
rect 34326 25542 38824 25594
rect 1104 25520 38824 25542
rect 12253 25483 12311 25489
rect 12253 25449 12265 25483
rect 12299 25480 12311 25483
rect 12342 25480 12348 25492
rect 12299 25452 12348 25480
rect 12299 25449 12311 25452
rect 12253 25443 12311 25449
rect 12342 25440 12348 25452
rect 12400 25440 12406 25492
rect 21818 25440 21824 25492
rect 21876 25480 21882 25492
rect 24397 25483 24455 25489
rect 24397 25480 24409 25483
rect 21876 25452 24409 25480
rect 21876 25440 21882 25452
rect 24397 25449 24409 25452
rect 24443 25449 24455 25483
rect 24397 25443 24455 25449
rect 12621 25347 12679 25353
rect 12621 25313 12633 25347
rect 12667 25344 12679 25347
rect 12710 25344 12716 25356
rect 12667 25316 12716 25344
rect 12667 25313 12679 25316
rect 12621 25307 12679 25313
rect 12710 25304 12716 25316
rect 12768 25304 12774 25356
rect 15562 25344 15568 25356
rect 15523 25316 15568 25344
rect 15562 25304 15568 25316
rect 15620 25304 15626 25356
rect 21818 25344 21824 25356
rect 21779 25316 21824 25344
rect 21818 25304 21824 25316
rect 21876 25304 21882 25356
rect 1673 25279 1731 25285
rect 1673 25245 1685 25279
rect 1719 25276 1731 25279
rect 12437 25279 12495 25285
rect 1719 25248 2268 25276
rect 1719 25245 1731 25248
rect 1673 25239 1731 25245
rect 2240 25152 2268 25248
rect 12437 25245 12449 25279
rect 12483 25276 12495 25279
rect 15010 25276 15016 25288
rect 12483 25248 15016 25276
rect 12483 25245 12495 25248
rect 12437 25239 12495 25245
rect 15010 25236 15016 25248
rect 15068 25236 15074 25288
rect 15838 25276 15844 25288
rect 15799 25248 15844 25276
rect 15838 25236 15844 25248
rect 15896 25236 15902 25288
rect 20530 25276 20536 25288
rect 20272 25248 20536 25276
rect 1486 25140 1492 25152
rect 1447 25112 1492 25140
rect 1486 25100 1492 25112
rect 1544 25100 1550 25152
rect 2222 25140 2228 25152
rect 2183 25112 2228 25140
rect 2222 25100 2228 25112
rect 2280 25100 2286 25152
rect 16577 25143 16635 25149
rect 16577 25109 16589 25143
rect 16623 25140 16635 25143
rect 17034 25140 17040 25152
rect 16623 25112 17040 25140
rect 16623 25109 16635 25112
rect 16577 25103 16635 25109
rect 17034 25100 17040 25112
rect 17092 25100 17098 25152
rect 19702 25100 19708 25152
rect 19760 25140 19766 25152
rect 20272 25149 20300 25248
rect 20530 25236 20536 25248
rect 20588 25276 20594 25288
rect 20809 25279 20867 25285
rect 20809 25276 20821 25279
rect 20588 25248 20821 25276
rect 20588 25236 20594 25248
rect 20809 25245 20821 25248
rect 20855 25245 20867 25279
rect 20809 25239 20867 25245
rect 20990 25236 20996 25288
rect 21048 25276 21054 25288
rect 22094 25276 22100 25288
rect 21048 25248 21141 25276
rect 22055 25248 22100 25276
rect 21048 25236 21054 25248
rect 21100 25208 21128 25248
rect 22094 25236 22100 25248
rect 22152 25236 22158 25288
rect 24581 25279 24639 25285
rect 24581 25245 24593 25279
rect 24627 25276 24639 25279
rect 25314 25276 25320 25288
rect 24627 25248 25320 25276
rect 24627 25245 24639 25248
rect 24581 25239 24639 25245
rect 25314 25236 25320 25248
rect 25372 25236 25378 25288
rect 27525 25279 27583 25285
rect 27525 25245 27537 25279
rect 27571 25245 27583 25279
rect 27798 25276 27804 25288
rect 27759 25248 27804 25276
rect 27525 25239 27583 25245
rect 25958 25208 25964 25220
rect 21100 25180 25964 25208
rect 25958 25168 25964 25180
rect 26016 25168 26022 25220
rect 27540 25208 27568 25239
rect 27798 25236 27804 25248
rect 27856 25236 27862 25288
rect 27706 25208 27712 25220
rect 27540 25180 27712 25208
rect 27706 25168 27712 25180
rect 27764 25168 27770 25220
rect 20257 25143 20315 25149
rect 20257 25140 20269 25143
rect 19760 25112 20269 25140
rect 19760 25100 19766 25112
rect 20257 25109 20269 25112
rect 20303 25109 20315 25143
rect 20257 25103 20315 25109
rect 21177 25143 21235 25149
rect 21177 25109 21189 25143
rect 21223 25140 21235 25143
rect 21818 25140 21824 25152
rect 21223 25112 21824 25140
rect 21223 25109 21235 25112
rect 21177 25103 21235 25109
rect 21818 25100 21824 25112
rect 21876 25100 21882 25152
rect 22830 25140 22836 25152
rect 22791 25112 22836 25140
rect 22830 25100 22836 25112
rect 22888 25140 22894 25152
rect 28537 25143 28595 25149
rect 28537 25140 28549 25143
rect 22888 25112 28549 25140
rect 22888 25100 22894 25112
rect 28537 25109 28549 25112
rect 28583 25140 28595 25143
rect 28718 25140 28724 25152
rect 28583 25112 28724 25140
rect 28583 25109 28595 25112
rect 28537 25103 28595 25109
rect 28718 25100 28724 25112
rect 28776 25100 28782 25152
rect 1104 25050 38824 25072
rect 1104 24998 10398 25050
rect 10450 24998 10462 25050
rect 10514 24998 10526 25050
rect 10578 24998 10590 25050
rect 10642 24998 10654 25050
rect 10706 24998 19846 25050
rect 19898 24998 19910 25050
rect 19962 24998 19974 25050
rect 20026 24998 20038 25050
rect 20090 24998 20102 25050
rect 20154 24998 29294 25050
rect 29346 24998 29358 25050
rect 29410 24998 29422 25050
rect 29474 24998 29486 25050
rect 29538 24998 29550 25050
rect 29602 24998 38824 25050
rect 1104 24976 38824 24998
rect 2222 24896 2228 24948
rect 2280 24936 2286 24948
rect 13262 24936 13268 24948
rect 2280 24908 13268 24936
rect 2280 24896 2286 24908
rect 13262 24896 13268 24908
rect 13320 24896 13326 24948
rect 15838 24896 15844 24948
rect 15896 24936 15902 24948
rect 15933 24939 15991 24945
rect 15933 24936 15945 24939
rect 15896 24908 15945 24936
rect 15896 24896 15902 24908
rect 15933 24905 15945 24908
rect 15979 24905 15991 24939
rect 15933 24899 15991 24905
rect 28353 24939 28411 24945
rect 28353 24905 28365 24939
rect 28399 24936 28411 24939
rect 28442 24936 28448 24948
rect 28399 24908 28448 24936
rect 28399 24905 28411 24908
rect 28353 24899 28411 24905
rect 28442 24896 28448 24908
rect 28500 24896 28506 24948
rect 14660 24840 15240 24868
rect 2314 24760 2320 24812
rect 2372 24800 2378 24812
rect 12713 24803 12771 24809
rect 12713 24800 12725 24803
rect 2372 24772 12725 24800
rect 2372 24760 2378 24772
rect 12713 24769 12725 24772
rect 12759 24800 12771 24803
rect 13449 24803 13507 24809
rect 13449 24800 13461 24803
rect 12759 24772 13461 24800
rect 12759 24769 12771 24772
rect 12713 24763 12771 24769
rect 13449 24769 13461 24772
rect 13495 24800 13507 24803
rect 14660 24800 14688 24840
rect 14921 24803 14979 24809
rect 14921 24800 14933 24803
rect 13495 24772 14688 24800
rect 14844 24772 14933 24800
rect 13495 24769 13507 24772
rect 13449 24763 13507 24769
rect 12710 24556 12716 24608
rect 12768 24596 12774 24608
rect 12805 24599 12863 24605
rect 12805 24596 12817 24599
rect 12768 24568 12817 24596
rect 12768 24556 12774 24568
rect 12805 24565 12817 24568
rect 12851 24565 12863 24599
rect 12805 24559 12863 24565
rect 13538 24556 13544 24608
rect 13596 24596 13602 24608
rect 14461 24599 14519 24605
rect 14461 24596 14473 24599
rect 13596 24568 14473 24596
rect 13596 24556 13602 24568
rect 14461 24565 14473 24568
rect 14507 24596 14519 24599
rect 14844 24596 14872 24772
rect 14921 24769 14933 24772
rect 14967 24769 14979 24803
rect 14921 24763 14979 24769
rect 15010 24760 15016 24812
rect 15068 24800 15074 24812
rect 15105 24803 15163 24809
rect 15105 24800 15117 24803
rect 15068 24772 15117 24800
rect 15068 24760 15074 24772
rect 15105 24769 15117 24772
rect 15151 24769 15163 24803
rect 15105 24763 15163 24769
rect 15212 24732 15240 24840
rect 15289 24803 15347 24809
rect 15289 24769 15301 24803
rect 15335 24800 15347 24803
rect 15749 24803 15807 24809
rect 15749 24800 15761 24803
rect 15335 24772 15761 24800
rect 15335 24769 15347 24772
rect 15289 24763 15347 24769
rect 15749 24769 15761 24772
rect 15795 24769 15807 24803
rect 15749 24763 15807 24769
rect 19610 24760 19616 24812
rect 19668 24800 19674 24812
rect 19981 24803 20039 24809
rect 19981 24800 19993 24803
rect 19668 24772 19993 24800
rect 19668 24760 19674 24772
rect 19981 24769 19993 24772
rect 20027 24769 20039 24803
rect 21818 24800 21824 24812
rect 21779 24772 21824 24800
rect 19981 24763 20039 24769
rect 21818 24760 21824 24772
rect 21876 24760 21882 24812
rect 25958 24760 25964 24812
rect 26016 24800 26022 24812
rect 28537 24803 28595 24809
rect 28537 24800 28549 24803
rect 26016 24772 28549 24800
rect 26016 24760 26022 24772
rect 28537 24769 28549 24772
rect 28583 24800 28595 24803
rect 28626 24800 28632 24812
rect 28583 24772 28632 24800
rect 28583 24769 28595 24772
rect 28537 24763 28595 24769
rect 28626 24760 28632 24772
rect 28684 24760 28690 24812
rect 32950 24800 32956 24812
rect 32911 24772 32956 24800
rect 32950 24760 32956 24772
rect 33008 24760 33014 24812
rect 33597 24803 33655 24809
rect 33597 24769 33609 24803
rect 33643 24769 33655 24803
rect 33597 24763 33655 24769
rect 28721 24735 28779 24741
rect 15212 24704 22094 24732
rect 20165 24667 20223 24673
rect 20165 24633 20177 24667
rect 20211 24664 20223 24667
rect 20990 24664 20996 24676
rect 20211 24636 20996 24664
rect 20211 24633 20223 24636
rect 20165 24627 20223 24633
rect 20990 24624 20996 24636
rect 21048 24624 21054 24676
rect 22066 24664 22094 24704
rect 28721 24701 28733 24735
rect 28767 24732 28779 24735
rect 31202 24732 31208 24744
rect 28767 24704 31208 24732
rect 28767 24701 28779 24704
rect 28721 24695 28779 24701
rect 31202 24692 31208 24704
rect 31260 24692 31266 24744
rect 32858 24692 32864 24744
rect 32916 24732 32922 24744
rect 33612 24732 33640 24763
rect 32916 24704 33640 24732
rect 32916 24692 32922 24704
rect 30558 24664 30564 24676
rect 22066 24636 30564 24664
rect 30558 24624 30564 24636
rect 30616 24624 30622 24676
rect 15654 24596 15660 24608
rect 14507 24568 15660 24596
rect 14507 24565 14519 24568
rect 14461 24559 14519 24565
rect 15654 24556 15660 24568
rect 15712 24556 15718 24608
rect 22005 24599 22063 24605
rect 22005 24565 22017 24599
rect 22051 24596 22063 24599
rect 22094 24596 22100 24608
rect 22051 24568 22100 24596
rect 22051 24565 22063 24568
rect 22005 24559 22063 24565
rect 22094 24556 22100 24568
rect 22152 24556 22158 24608
rect 33134 24596 33140 24608
rect 33095 24568 33140 24596
rect 33134 24556 33140 24568
rect 33192 24556 33198 24608
rect 33778 24596 33784 24608
rect 33739 24568 33784 24596
rect 33778 24556 33784 24568
rect 33836 24556 33842 24608
rect 1104 24506 38824 24528
rect 1104 24454 5674 24506
rect 5726 24454 5738 24506
rect 5790 24454 5802 24506
rect 5854 24454 5866 24506
rect 5918 24454 5930 24506
rect 5982 24454 15122 24506
rect 15174 24454 15186 24506
rect 15238 24454 15250 24506
rect 15302 24454 15314 24506
rect 15366 24454 15378 24506
rect 15430 24454 24570 24506
rect 24622 24454 24634 24506
rect 24686 24454 24698 24506
rect 24750 24454 24762 24506
rect 24814 24454 24826 24506
rect 24878 24454 34018 24506
rect 34070 24454 34082 24506
rect 34134 24454 34146 24506
rect 34198 24454 34210 24506
rect 34262 24454 34274 24506
rect 34326 24454 38824 24506
rect 1104 24432 38824 24454
rect 19702 24256 19708 24268
rect 6886 24228 19708 24256
rect 3053 24191 3111 24197
rect 3053 24157 3065 24191
rect 3099 24188 3111 24191
rect 3789 24191 3847 24197
rect 3789 24188 3801 24191
rect 3099 24160 3801 24188
rect 3099 24157 3111 24160
rect 3053 24151 3111 24157
rect 3789 24157 3801 24160
rect 3835 24157 3847 24191
rect 3970 24188 3976 24200
rect 3931 24160 3976 24188
rect 3789 24151 3847 24157
rect 3970 24148 3976 24160
rect 4028 24148 4034 24200
rect 4154 24188 4160 24200
rect 4115 24160 4160 24188
rect 4154 24148 4160 24160
rect 4212 24188 4218 24200
rect 4614 24188 4620 24200
rect 4212 24160 4620 24188
rect 4212 24148 4218 24160
rect 4614 24148 4620 24160
rect 4672 24148 4678 24200
rect 4632 24120 4660 24148
rect 6886 24120 6914 24228
rect 19702 24216 19708 24228
rect 19760 24216 19766 24268
rect 20990 24256 20996 24268
rect 20088 24228 20996 24256
rect 8938 24188 8944 24200
rect 8899 24160 8944 24188
rect 8938 24148 8944 24160
rect 8996 24148 9002 24200
rect 9214 24188 9220 24200
rect 9175 24160 9220 24188
rect 9214 24148 9220 24160
rect 9272 24148 9278 24200
rect 19429 24191 19487 24197
rect 19429 24157 19441 24191
rect 19475 24188 19487 24191
rect 19518 24188 19524 24200
rect 19475 24160 19524 24188
rect 19475 24157 19487 24160
rect 19429 24151 19487 24157
rect 19518 24148 19524 24160
rect 19576 24188 19582 24200
rect 20088 24197 20116 24228
rect 20990 24216 20996 24228
rect 21048 24216 21054 24268
rect 28445 24259 28503 24265
rect 28445 24225 28457 24259
rect 28491 24256 28503 24259
rect 28534 24256 28540 24268
rect 28491 24228 28540 24256
rect 28491 24225 28503 24228
rect 28445 24219 28503 24225
rect 28534 24216 28540 24228
rect 28592 24256 28598 24268
rect 31294 24256 31300 24268
rect 28592 24228 31300 24256
rect 28592 24216 28598 24228
rect 31294 24216 31300 24228
rect 31352 24216 31358 24268
rect 19889 24191 19947 24197
rect 19889 24188 19901 24191
rect 19576 24160 19901 24188
rect 19576 24148 19582 24160
rect 19889 24157 19901 24160
rect 19935 24157 19947 24191
rect 19889 24151 19947 24157
rect 20073 24191 20131 24197
rect 20073 24157 20085 24191
rect 20119 24157 20131 24191
rect 20073 24151 20131 24157
rect 20257 24191 20315 24197
rect 20257 24157 20269 24191
rect 20303 24188 20315 24191
rect 20901 24191 20959 24197
rect 20901 24188 20913 24191
rect 20303 24160 20913 24188
rect 20303 24157 20315 24160
rect 20257 24151 20315 24157
rect 20901 24157 20913 24160
rect 20947 24157 20959 24191
rect 28626 24188 28632 24200
rect 28587 24160 28632 24188
rect 20901 24151 20959 24157
rect 28626 24148 28632 24160
rect 28684 24148 28690 24200
rect 32858 24188 32864 24200
rect 30944 24160 32864 24188
rect 4632 24092 6914 24120
rect 28534 24080 28540 24132
rect 28592 24120 28598 24132
rect 30944 24120 30972 24160
rect 32858 24148 32864 24160
rect 32916 24148 32922 24200
rect 33134 24188 33140 24200
rect 33095 24160 33140 24188
rect 33134 24148 33140 24160
rect 33192 24148 33198 24200
rect 33870 24148 33876 24200
rect 33928 24188 33934 24200
rect 33965 24191 34023 24197
rect 33965 24188 33977 24191
rect 33928 24160 33977 24188
rect 33928 24148 33934 24160
rect 33965 24157 33977 24160
rect 34011 24157 34023 24191
rect 33965 24151 34023 24157
rect 31113 24123 31171 24129
rect 31113 24120 31125 24123
rect 28592 24092 30972 24120
rect 31036 24092 31125 24120
rect 28592 24080 28598 24092
rect 3237 24055 3295 24061
rect 3237 24021 3249 24055
rect 3283 24052 3295 24055
rect 3602 24052 3608 24064
rect 3283 24024 3608 24052
rect 3283 24021 3295 24024
rect 3237 24015 3295 24021
rect 3602 24012 3608 24024
rect 3660 24012 3666 24064
rect 20622 24012 20628 24064
rect 20680 24052 20686 24064
rect 20717 24055 20775 24061
rect 20717 24052 20729 24055
rect 20680 24024 20729 24052
rect 20680 24012 20686 24024
rect 20717 24021 20729 24024
rect 20763 24021 20775 24055
rect 28810 24052 28816 24064
rect 28771 24024 28816 24052
rect 20717 24015 20775 24021
rect 28810 24012 28816 24024
rect 28868 24012 28874 24064
rect 30558 24012 30564 24064
rect 30616 24052 30622 24064
rect 31036 24052 31064 24092
rect 31113 24089 31125 24092
rect 31159 24120 31171 24123
rect 31757 24123 31815 24129
rect 31757 24120 31769 24123
rect 31159 24092 31769 24120
rect 31159 24089 31171 24092
rect 31113 24083 31171 24089
rect 31757 24089 31769 24092
rect 31803 24089 31815 24123
rect 31757 24083 31815 24089
rect 31202 24052 31208 24064
rect 30616 24024 31064 24052
rect 31163 24024 31208 24052
rect 30616 24012 30622 24024
rect 31202 24012 31208 24024
rect 31260 24012 31266 24064
rect 1104 23962 38824 23984
rect 1104 23910 10398 23962
rect 10450 23910 10462 23962
rect 10514 23910 10526 23962
rect 10578 23910 10590 23962
rect 10642 23910 10654 23962
rect 10706 23910 19846 23962
rect 19898 23910 19910 23962
rect 19962 23910 19974 23962
rect 20026 23910 20038 23962
rect 20090 23910 20102 23962
rect 20154 23910 29294 23962
rect 29346 23910 29358 23962
rect 29410 23910 29422 23962
rect 29474 23910 29486 23962
rect 29538 23910 29550 23962
rect 29602 23910 38824 23962
rect 1104 23888 38824 23910
rect 8018 23848 8024 23860
rect 7979 23820 8024 23848
rect 8018 23808 8024 23820
rect 8076 23808 8082 23860
rect 8386 23808 8392 23860
rect 8444 23848 8450 23860
rect 8481 23851 8539 23857
rect 8481 23848 8493 23851
rect 8444 23820 8493 23848
rect 8444 23808 8450 23820
rect 8481 23817 8493 23820
rect 8527 23817 8539 23851
rect 8481 23811 8539 23817
rect 25866 23808 25872 23860
rect 25924 23848 25930 23860
rect 28534 23848 28540 23860
rect 25924 23820 28540 23848
rect 25924 23808 25930 23820
rect 28534 23808 28540 23820
rect 28592 23808 28598 23860
rect 28718 23848 28724 23860
rect 28679 23820 28724 23848
rect 28718 23808 28724 23820
rect 28776 23808 28782 23860
rect 29181 23851 29239 23857
rect 29181 23817 29193 23851
rect 29227 23817 29239 23851
rect 32950 23848 32956 23860
rect 32911 23820 32956 23848
rect 29181 23811 29239 23817
rect 9490 23780 9496 23792
rect 7852 23752 9496 23780
rect 1673 23715 1731 23721
rect 1673 23681 1685 23715
rect 1719 23712 1731 23715
rect 1854 23712 1860 23724
rect 1719 23684 1860 23712
rect 1719 23681 1731 23684
rect 1673 23675 1731 23681
rect 1854 23672 1860 23684
rect 1912 23672 1918 23724
rect 3602 23712 3608 23724
rect 3563 23684 3608 23712
rect 3602 23672 3608 23684
rect 3660 23672 3666 23724
rect 7852 23721 7880 23752
rect 9490 23740 9496 23752
rect 9548 23740 9554 23792
rect 13449 23783 13507 23789
rect 13449 23749 13461 23783
rect 13495 23780 13507 23783
rect 13538 23780 13544 23792
rect 13495 23752 13544 23780
rect 13495 23749 13507 23752
rect 13449 23743 13507 23749
rect 13538 23740 13544 23752
rect 13596 23740 13602 23792
rect 29196 23780 29224 23811
rect 32950 23808 32956 23820
rect 33008 23808 33014 23860
rect 33870 23808 33876 23860
rect 33928 23848 33934 23860
rect 36722 23848 36728 23860
rect 33928 23820 36728 23848
rect 33928 23808 33934 23820
rect 36722 23808 36728 23820
rect 36780 23808 36786 23860
rect 28000 23752 29224 23780
rect 3881 23715 3939 23721
rect 3881 23681 3893 23715
rect 3927 23712 3939 23715
rect 7837 23715 7895 23721
rect 7837 23712 7849 23715
rect 3927 23684 7849 23712
rect 3927 23681 3939 23684
rect 3881 23675 3939 23681
rect 7837 23681 7849 23684
rect 7883 23681 7895 23715
rect 7837 23675 7895 23681
rect 9217 23715 9275 23721
rect 9217 23681 9229 23715
rect 9263 23712 9275 23715
rect 9858 23712 9864 23724
rect 9263 23684 9864 23712
rect 9263 23681 9275 23684
rect 9217 23675 9275 23681
rect 9858 23672 9864 23684
rect 9916 23672 9922 23724
rect 13262 23712 13268 23724
rect 13175 23684 13268 23712
rect 13262 23672 13268 23684
rect 13320 23712 13326 23724
rect 13906 23712 13912 23724
rect 13320 23684 13912 23712
rect 13320 23672 13326 23684
rect 13906 23672 13912 23684
rect 13964 23672 13970 23724
rect 16850 23712 16856 23724
rect 16811 23684 16856 23712
rect 16850 23672 16856 23684
rect 16908 23672 16914 23724
rect 20622 23712 20628 23724
rect 20583 23684 20628 23712
rect 20622 23672 20628 23684
rect 20680 23672 20686 23724
rect 20898 23712 20904 23724
rect 20811 23684 20904 23712
rect 20898 23672 20904 23684
rect 20956 23712 20962 23724
rect 21726 23712 21732 23724
rect 20956 23684 21732 23712
rect 20956 23672 20962 23684
rect 21726 23672 21732 23684
rect 21784 23672 21790 23724
rect 28000 23721 28028 23752
rect 33778 23740 33784 23792
rect 33836 23780 33842 23792
rect 33836 23752 35664 23780
rect 33836 23740 33842 23752
rect 27985 23715 28043 23721
rect 27985 23681 27997 23715
rect 28031 23681 28043 23715
rect 27985 23675 28043 23681
rect 28810 23672 28816 23724
rect 28868 23712 28874 23724
rect 29365 23715 29423 23721
rect 29365 23712 29377 23715
rect 28868 23684 29377 23712
rect 28868 23672 28874 23684
rect 29365 23681 29377 23684
rect 29411 23681 29423 23715
rect 31294 23712 31300 23724
rect 31255 23684 31300 23712
rect 29365 23675 29423 23681
rect 31294 23672 31300 23684
rect 31352 23672 31358 23724
rect 31846 23672 31852 23724
rect 31904 23712 31910 23724
rect 35636 23721 35664 23752
rect 32769 23715 32827 23721
rect 32769 23712 32781 23715
rect 31904 23684 32781 23712
rect 31904 23672 31910 23684
rect 32769 23681 32781 23684
rect 32815 23712 32827 23715
rect 34793 23715 34851 23721
rect 34793 23712 34805 23715
rect 32815 23684 34805 23712
rect 32815 23681 32827 23684
rect 32769 23675 32827 23681
rect 34793 23681 34805 23684
rect 34839 23681 34851 23715
rect 34793 23675 34851 23681
rect 35621 23715 35679 23721
rect 35621 23681 35633 23715
rect 35667 23681 35679 23715
rect 35621 23675 35679 23681
rect 35894 23672 35900 23724
rect 35952 23712 35958 23724
rect 36722 23712 36728 23724
rect 35952 23684 35997 23712
rect 36683 23684 36728 23712
rect 35952 23672 35958 23684
rect 36722 23672 36728 23684
rect 36780 23672 36786 23724
rect 9490 23604 9496 23656
rect 9548 23644 9554 23656
rect 27706 23644 27712 23656
rect 9548 23616 9593 23644
rect 27667 23616 27712 23644
rect 9548 23604 9554 23616
rect 27706 23604 27712 23616
rect 27764 23604 27770 23656
rect 31573 23647 31631 23653
rect 31573 23613 31585 23647
rect 31619 23644 31631 23647
rect 32030 23644 32036 23656
rect 31619 23616 32036 23644
rect 31619 23613 31631 23616
rect 31573 23607 31631 23613
rect 30285 23579 30343 23585
rect 30285 23545 30297 23579
rect 30331 23576 30343 23579
rect 31588 23576 31616 23607
rect 32030 23604 32036 23616
rect 32088 23604 32094 23656
rect 32585 23647 32643 23653
rect 32585 23644 32597 23647
rect 32140 23616 32597 23644
rect 30331 23548 31616 23576
rect 30331 23545 30343 23548
rect 30285 23539 30343 23545
rect 1486 23508 1492 23520
rect 1447 23480 1492 23508
rect 1486 23468 1492 23480
rect 1544 23468 1550 23520
rect 2866 23508 2872 23520
rect 2827 23480 2872 23508
rect 2866 23468 2872 23480
rect 2924 23468 2930 23520
rect 9950 23508 9956 23520
rect 9911 23480 9956 23508
rect 9950 23468 9956 23480
rect 10008 23508 10014 23520
rect 12250 23508 12256 23520
rect 10008 23480 12256 23508
rect 10008 23468 10014 23480
rect 12250 23468 12256 23480
rect 12308 23468 12314 23520
rect 13906 23508 13912 23520
rect 13867 23480 13912 23508
rect 13906 23468 13912 23480
rect 13964 23468 13970 23520
rect 16666 23508 16672 23520
rect 16627 23480 16672 23508
rect 16666 23468 16672 23480
rect 16724 23468 16730 23520
rect 19889 23511 19947 23517
rect 19889 23477 19901 23511
rect 19935 23508 19947 23511
rect 20990 23508 20996 23520
rect 19935 23480 20996 23508
rect 19935 23477 19947 23480
rect 19889 23471 19947 23477
rect 20990 23468 20996 23480
rect 21048 23508 21054 23520
rect 22830 23508 22836 23520
rect 21048 23480 22836 23508
rect 21048 23468 21054 23480
rect 22830 23468 22836 23480
rect 22888 23468 22894 23520
rect 31294 23468 31300 23520
rect 31352 23508 31358 23520
rect 32140 23508 32168 23616
rect 32585 23613 32597 23616
rect 32631 23613 32643 23647
rect 32585 23607 32643 23613
rect 34149 23647 34207 23653
rect 34149 23613 34161 23647
rect 34195 23644 34207 23647
rect 34606 23644 34612 23656
rect 34195 23616 34612 23644
rect 34195 23613 34207 23616
rect 34149 23607 34207 23613
rect 34606 23604 34612 23616
rect 34664 23604 34670 23656
rect 31352 23480 32168 23508
rect 34977 23511 35035 23517
rect 31352 23468 31358 23480
rect 34977 23477 34989 23511
rect 35023 23508 35035 23511
rect 35526 23508 35532 23520
rect 35023 23480 35532 23508
rect 35023 23477 35035 23480
rect 34977 23471 35035 23477
rect 35526 23468 35532 23480
rect 35584 23468 35590 23520
rect 1104 23418 38824 23440
rect 1104 23366 5674 23418
rect 5726 23366 5738 23418
rect 5790 23366 5802 23418
rect 5854 23366 5866 23418
rect 5918 23366 5930 23418
rect 5982 23366 15122 23418
rect 15174 23366 15186 23418
rect 15238 23366 15250 23418
rect 15302 23366 15314 23418
rect 15366 23366 15378 23418
rect 15430 23366 24570 23418
rect 24622 23366 24634 23418
rect 24686 23366 24698 23418
rect 24750 23366 24762 23418
rect 24814 23366 24826 23418
rect 24878 23366 34018 23418
rect 34070 23366 34082 23418
rect 34134 23366 34146 23418
rect 34198 23366 34210 23418
rect 34262 23366 34274 23418
rect 34326 23366 38824 23418
rect 1104 23344 38824 23366
rect 9858 23304 9864 23316
rect 9819 23276 9864 23304
rect 9858 23264 9864 23276
rect 9916 23264 9922 23316
rect 15381 23307 15439 23313
rect 15381 23273 15393 23307
rect 15427 23304 15439 23307
rect 15562 23304 15568 23316
rect 15427 23276 15568 23304
rect 15427 23273 15439 23276
rect 15381 23267 15439 23273
rect 15562 23264 15568 23276
rect 15620 23264 15626 23316
rect 35713 23307 35771 23313
rect 35713 23273 35725 23307
rect 35759 23304 35771 23307
rect 35894 23304 35900 23316
rect 35759 23276 35900 23304
rect 35759 23273 35771 23276
rect 35713 23267 35771 23273
rect 35894 23264 35900 23276
rect 35952 23264 35958 23316
rect 5537 23171 5595 23177
rect 5537 23137 5549 23171
rect 5583 23168 5595 23171
rect 6914 23168 6920 23180
rect 5583 23140 6920 23168
rect 5583 23137 5595 23140
rect 5537 23131 5595 23137
rect 6914 23128 6920 23140
rect 6972 23128 6978 23180
rect 8938 23128 8944 23180
rect 8996 23168 9002 23180
rect 9582 23168 9588 23180
rect 8996 23140 9588 23168
rect 8996 23128 9002 23140
rect 5442 23060 5448 23112
rect 5500 23100 5506 23112
rect 5721 23103 5779 23109
rect 5721 23100 5733 23103
rect 5500 23072 5733 23100
rect 5500 23060 5506 23072
rect 5721 23069 5733 23072
rect 5767 23069 5779 23103
rect 9030 23100 9036 23112
rect 8991 23072 9036 23100
rect 5721 23063 5779 23069
rect 9030 23060 9036 23072
rect 9088 23060 9094 23112
rect 9232 23109 9260 23140
rect 9582 23128 9588 23140
rect 9640 23128 9646 23180
rect 31205 23171 31263 23177
rect 31205 23137 31217 23171
rect 31251 23168 31263 23171
rect 31846 23168 31852 23180
rect 31251 23140 31852 23168
rect 31251 23137 31263 23140
rect 31205 23131 31263 23137
rect 31846 23128 31852 23140
rect 31904 23128 31910 23180
rect 9217 23103 9275 23109
rect 9217 23069 9229 23103
rect 9263 23069 9275 23103
rect 9217 23063 9275 23069
rect 9401 23103 9459 23109
rect 9401 23069 9413 23103
rect 9447 23100 9459 23103
rect 10045 23103 10103 23109
rect 10045 23100 10057 23103
rect 9447 23072 10057 23100
rect 9447 23069 9459 23072
rect 9401 23063 9459 23069
rect 10045 23069 10057 23072
rect 10091 23069 10103 23103
rect 10045 23063 10103 23069
rect 11698 23060 11704 23112
rect 11756 23100 11762 23112
rect 15565 23103 15623 23109
rect 15565 23100 15577 23103
rect 11756 23072 15577 23100
rect 11756 23060 11762 23072
rect 15565 23069 15577 23072
rect 15611 23100 15623 23103
rect 16025 23103 16083 23109
rect 16025 23100 16037 23103
rect 15611 23072 16037 23100
rect 15611 23069 15623 23072
rect 15565 23063 15623 23069
rect 16025 23069 16037 23072
rect 16071 23069 16083 23103
rect 16025 23063 16083 23069
rect 16301 23103 16359 23109
rect 16301 23069 16313 23103
rect 16347 23100 16359 23103
rect 16666 23100 16672 23112
rect 16347 23072 16672 23100
rect 16347 23069 16359 23072
rect 16301 23063 16359 23069
rect 16666 23060 16672 23072
rect 16724 23060 16730 23112
rect 30926 23100 30932 23112
rect 30887 23072 30932 23100
rect 30926 23060 30932 23072
rect 30984 23060 30990 23112
rect 35526 23100 35532 23112
rect 35487 23072 35532 23100
rect 35526 23060 35532 23072
rect 35584 23060 35590 23112
rect 9048 23032 9076 23060
rect 9950 23032 9956 23044
rect 9048 23004 9956 23032
rect 9950 22992 9956 23004
rect 10008 22992 10014 23044
rect 5905 22967 5963 22973
rect 5905 22933 5917 22967
rect 5951 22964 5963 22967
rect 5994 22964 6000 22976
rect 5951 22936 6000 22964
rect 5951 22933 5963 22936
rect 5905 22927 5963 22933
rect 5994 22924 6000 22936
rect 6052 22924 6058 22976
rect 17034 22964 17040 22976
rect 16995 22936 17040 22964
rect 17034 22924 17040 22936
rect 17092 22924 17098 22976
rect 1104 22874 38824 22896
rect 1104 22822 10398 22874
rect 10450 22822 10462 22874
rect 10514 22822 10526 22874
rect 10578 22822 10590 22874
rect 10642 22822 10654 22874
rect 10706 22822 19846 22874
rect 19898 22822 19910 22874
rect 19962 22822 19974 22874
rect 20026 22822 20038 22874
rect 20090 22822 20102 22874
rect 20154 22822 29294 22874
rect 29346 22822 29358 22874
rect 29410 22822 29422 22874
rect 29474 22822 29486 22874
rect 29538 22822 29550 22874
rect 29602 22822 38824 22874
rect 1104 22800 38824 22822
rect 3878 22760 3884 22772
rect 3344 22732 3884 22760
rect 3344 22633 3372 22732
rect 3878 22720 3884 22732
rect 3936 22720 3942 22772
rect 9490 22720 9496 22772
rect 9548 22760 9554 22772
rect 9953 22763 10011 22769
rect 9953 22760 9965 22763
rect 9548 22732 9965 22760
rect 9548 22720 9554 22732
rect 9953 22729 9965 22732
rect 9999 22729 10011 22763
rect 9953 22723 10011 22729
rect 16669 22763 16727 22769
rect 16669 22729 16681 22763
rect 16715 22760 16727 22763
rect 16850 22760 16856 22772
rect 16715 22732 16856 22760
rect 16715 22729 16727 22732
rect 16669 22723 16727 22729
rect 16850 22720 16856 22732
rect 16908 22720 16914 22772
rect 12636 22664 14780 22692
rect 3145 22627 3203 22633
rect 3145 22593 3157 22627
rect 3191 22593 3203 22627
rect 3145 22587 3203 22593
rect 3329 22627 3387 22633
rect 3329 22593 3341 22627
rect 3375 22593 3387 22627
rect 3329 22587 3387 22593
rect 3160 22556 3188 22587
rect 4614 22584 4620 22636
rect 4672 22624 4678 22636
rect 5442 22624 5448 22636
rect 4672 22596 5448 22624
rect 4672 22584 4678 22596
rect 5442 22584 5448 22596
rect 5500 22624 5506 22636
rect 7009 22627 7067 22633
rect 7009 22624 7021 22627
rect 5500 22596 7021 22624
rect 5500 22584 5506 22596
rect 7009 22593 7021 22596
rect 7055 22593 7067 22627
rect 10134 22624 10140 22636
rect 10095 22596 10140 22624
rect 7009 22587 7067 22593
rect 10134 22584 10140 22596
rect 10192 22584 10198 22636
rect 12636 22633 12664 22664
rect 14752 22636 14780 22664
rect 12621 22627 12679 22633
rect 12621 22593 12633 22627
rect 12667 22593 12679 22627
rect 12621 22587 12679 22593
rect 12805 22627 12863 22633
rect 12805 22593 12817 22627
rect 12851 22624 12863 22627
rect 13449 22627 13507 22633
rect 13449 22624 13461 22627
rect 12851 22596 13461 22624
rect 12851 22593 12863 22596
rect 12805 22587 12863 22593
rect 13449 22593 13461 22596
rect 13495 22593 13507 22627
rect 13449 22587 13507 22593
rect 14734 22584 14740 22636
rect 14792 22624 14798 22636
rect 15010 22624 15016 22636
rect 14792 22596 15016 22624
rect 14792 22584 14798 22596
rect 15010 22584 15016 22596
rect 15068 22624 15074 22636
rect 16853 22627 16911 22633
rect 16853 22624 16865 22627
rect 15068 22596 16865 22624
rect 15068 22584 15074 22596
rect 16853 22593 16865 22596
rect 16899 22593 16911 22627
rect 16853 22587 16911 22593
rect 17037 22627 17095 22633
rect 17037 22593 17049 22627
rect 17083 22624 17095 22627
rect 17497 22627 17555 22633
rect 17497 22624 17509 22627
rect 17083 22596 17509 22624
rect 17083 22593 17095 22596
rect 17037 22587 17095 22593
rect 17497 22593 17509 22596
rect 17543 22624 17555 22627
rect 20806 22624 20812 22636
rect 17543 22596 20812 22624
rect 17543 22593 17555 22596
rect 17497 22587 17555 22593
rect 20806 22584 20812 22596
rect 20864 22584 20870 22636
rect 25682 22624 25688 22636
rect 25643 22596 25688 22624
rect 25682 22584 25688 22596
rect 25740 22584 25746 22636
rect 4632 22556 4660 22584
rect 3160 22528 4660 22556
rect 7193 22559 7251 22565
rect 7193 22525 7205 22559
rect 7239 22556 7251 22559
rect 7374 22556 7380 22568
rect 7239 22528 7380 22556
rect 7239 22525 7251 22528
rect 7193 22519 7251 22525
rect 7374 22516 7380 22528
rect 7432 22556 7438 22568
rect 12437 22559 12495 22565
rect 12437 22556 12449 22559
rect 7432 22528 12449 22556
rect 7432 22516 7438 22528
rect 12437 22525 12449 22528
rect 12483 22556 12495 22559
rect 13814 22556 13820 22568
rect 12483 22528 13820 22556
rect 12483 22525 12495 22528
rect 12437 22519 12495 22525
rect 13814 22516 13820 22528
rect 13872 22516 13878 22568
rect 3878 22448 3884 22500
rect 3936 22488 3942 22500
rect 13538 22488 13544 22500
rect 3936 22460 13544 22488
rect 3936 22448 3942 22460
rect 13538 22448 13544 22460
rect 13596 22448 13602 22500
rect 1394 22420 1400 22432
rect 1355 22392 1400 22420
rect 1394 22380 1400 22392
rect 1452 22380 1458 22432
rect 2961 22423 3019 22429
rect 2961 22389 2973 22423
rect 3007 22420 3019 22423
rect 3050 22420 3056 22432
rect 3007 22392 3056 22420
rect 3007 22389 3019 22392
rect 2961 22383 3019 22389
rect 3050 22380 3056 22392
rect 3108 22380 3114 22432
rect 6825 22423 6883 22429
rect 6825 22389 6837 22423
rect 6871 22420 6883 22423
rect 6914 22420 6920 22432
rect 6871 22392 6920 22420
rect 6871 22389 6883 22392
rect 6825 22383 6883 22389
rect 6914 22380 6920 22392
rect 6972 22380 6978 22432
rect 12986 22380 12992 22432
rect 13044 22420 13050 22432
rect 13265 22423 13323 22429
rect 13265 22420 13277 22423
rect 13044 22392 13277 22420
rect 13044 22380 13050 22392
rect 13265 22389 13277 22392
rect 13311 22389 13323 22423
rect 13265 22383 13323 22389
rect 25869 22423 25927 22429
rect 25869 22389 25881 22423
rect 25915 22420 25927 22423
rect 26234 22420 26240 22432
rect 25915 22392 26240 22420
rect 25915 22389 25927 22392
rect 25869 22383 25927 22389
rect 26234 22380 26240 22392
rect 26292 22380 26298 22432
rect 1104 22330 38824 22352
rect 1104 22278 5674 22330
rect 5726 22278 5738 22330
rect 5790 22278 5802 22330
rect 5854 22278 5866 22330
rect 5918 22278 5930 22330
rect 5982 22278 15122 22330
rect 15174 22278 15186 22330
rect 15238 22278 15250 22330
rect 15302 22278 15314 22330
rect 15366 22278 15378 22330
rect 15430 22278 24570 22330
rect 24622 22278 24634 22330
rect 24686 22278 24698 22330
rect 24750 22278 24762 22330
rect 24814 22278 24826 22330
rect 24878 22278 34018 22330
rect 34070 22278 34082 22330
rect 34134 22278 34146 22330
rect 34198 22278 34210 22330
rect 34262 22278 34274 22330
rect 34326 22278 38824 22330
rect 1104 22256 38824 22278
rect 10134 22176 10140 22228
rect 10192 22216 10198 22228
rect 10781 22219 10839 22225
rect 10781 22216 10793 22219
rect 10192 22188 10793 22216
rect 10192 22176 10198 22188
rect 10781 22185 10793 22188
rect 10827 22185 10839 22219
rect 10781 22179 10839 22185
rect 11698 22176 11704 22228
rect 11756 22216 11762 22228
rect 11793 22219 11851 22225
rect 11793 22216 11805 22219
rect 11756 22188 11805 22216
rect 11756 22176 11762 22188
rect 11793 22185 11805 22188
rect 11839 22216 11851 22219
rect 11839 22188 13308 22216
rect 11839 22185 11851 22188
rect 11793 22179 11851 22185
rect 13280 22089 13308 22188
rect 13265 22083 13323 22089
rect 13265 22049 13277 22083
rect 13311 22049 13323 22083
rect 14734 22080 14740 22092
rect 14695 22052 14740 22080
rect 13265 22043 13323 22049
rect 14734 22040 14740 22052
rect 14792 22040 14798 22092
rect 23474 22040 23480 22092
rect 23532 22080 23538 22092
rect 24394 22080 24400 22092
rect 23532 22052 24400 22080
rect 23532 22040 23538 22052
rect 24394 22040 24400 22052
rect 24452 22040 24458 22092
rect 5813 22015 5871 22021
rect 5813 21981 5825 22015
rect 5859 22012 5871 22015
rect 5994 22012 6000 22024
rect 5859 21984 6000 22012
rect 5859 21981 5871 21984
rect 5813 21975 5871 21981
rect 5994 21972 6000 21984
rect 6052 21972 6058 22024
rect 6914 21972 6920 22024
rect 6972 22012 6978 22024
rect 6972 21984 7017 22012
rect 6972 21972 6978 21984
rect 10042 21972 10048 22024
rect 10100 22012 10106 22024
rect 11149 22015 11207 22021
rect 11149 22012 11161 22015
rect 10100 21984 11161 22012
rect 10100 21972 10106 21984
rect 11149 21981 11161 21984
rect 11195 22012 11207 22015
rect 11609 22015 11667 22021
rect 11609 22012 11621 22015
rect 11195 21984 11621 22012
rect 11195 21981 11207 21984
rect 11149 21975 11207 21981
rect 11609 21981 11621 21984
rect 11655 21981 11667 22015
rect 12986 22012 12992 22024
rect 12947 21984 12992 22012
rect 11609 21975 11667 21981
rect 12986 21972 12992 21984
rect 13044 21972 13050 22024
rect 15013 22015 15071 22021
rect 15013 21981 15025 22015
rect 15059 21981 15071 22015
rect 23658 22012 23664 22024
rect 23619 21984 23664 22012
rect 15013 21975 15071 21981
rect 10965 21947 11023 21953
rect 10965 21913 10977 21947
rect 11011 21944 11023 21947
rect 12066 21944 12072 21956
rect 11011 21916 12072 21944
rect 11011 21913 11023 21916
rect 10965 21907 11023 21913
rect 12066 21904 12072 21916
rect 12124 21944 12130 21956
rect 14826 21944 14832 21956
rect 12124 21916 14832 21944
rect 12124 21904 12130 21916
rect 14826 21904 14832 21916
rect 14884 21944 14890 21956
rect 15028 21944 15056 21975
rect 23658 21972 23664 21984
rect 23716 21972 23722 22024
rect 24673 22015 24731 22021
rect 24673 21981 24685 22015
rect 24719 21981 24731 22015
rect 24673 21975 24731 21981
rect 14884 21916 15056 21944
rect 14884 21904 14890 21916
rect 5994 21876 6000 21888
rect 5955 21848 6000 21876
rect 5994 21836 6000 21848
rect 6052 21836 6058 21888
rect 7006 21836 7012 21888
rect 7064 21876 7070 21888
rect 7101 21879 7159 21885
rect 7101 21876 7113 21879
rect 7064 21848 7113 21876
rect 7064 21836 7070 21848
rect 7101 21845 7113 21848
rect 7147 21845 7159 21879
rect 7101 21839 7159 21845
rect 12158 21836 12164 21888
rect 12216 21876 12222 21888
rect 12253 21879 12311 21885
rect 12253 21876 12265 21879
rect 12216 21848 12265 21876
rect 12216 21836 12222 21848
rect 12253 21845 12265 21848
rect 12299 21876 12311 21879
rect 12342 21876 12348 21888
rect 12299 21848 12348 21876
rect 12299 21845 12311 21848
rect 12253 21839 12311 21845
rect 12342 21836 12348 21848
rect 12400 21836 12406 21888
rect 23845 21879 23903 21885
rect 23845 21845 23857 21879
rect 23891 21876 23903 21879
rect 24688 21876 24716 21975
rect 25866 21972 25872 22024
rect 25924 22012 25930 22024
rect 25961 22015 26019 22021
rect 25961 22012 25973 22015
rect 25924 21984 25973 22012
rect 25924 21972 25930 21984
rect 25961 21981 25973 21984
rect 26007 21981 26019 22015
rect 26234 22012 26240 22024
rect 26195 21984 26240 22012
rect 25961 21975 26019 21981
rect 26234 21972 26240 21984
rect 26292 21972 26298 22024
rect 27062 22012 27068 22024
rect 27023 21984 27068 22012
rect 27062 21972 27068 21984
rect 27120 22012 27126 22024
rect 33870 22012 33876 22024
rect 27120 21984 33876 22012
rect 27120 21972 27126 21984
rect 33870 21972 33876 21984
rect 33928 21972 33934 22024
rect 25406 21876 25412 21888
rect 23891 21848 24716 21876
rect 25367 21848 25412 21876
rect 23891 21845 23903 21848
rect 23845 21839 23903 21845
rect 25406 21836 25412 21848
rect 25464 21836 25470 21888
rect 1104 21786 38824 21808
rect 1104 21734 10398 21786
rect 10450 21734 10462 21786
rect 10514 21734 10526 21786
rect 10578 21734 10590 21786
rect 10642 21734 10654 21786
rect 10706 21734 19846 21786
rect 19898 21734 19910 21786
rect 19962 21734 19974 21786
rect 20026 21734 20038 21786
rect 20090 21734 20102 21786
rect 20154 21734 29294 21786
rect 29346 21734 29358 21786
rect 29410 21734 29422 21786
rect 29474 21734 29486 21786
rect 29538 21734 29550 21786
rect 29602 21734 38824 21786
rect 1104 21712 38824 21734
rect 18969 21675 19027 21681
rect 18969 21641 18981 21675
rect 19015 21672 19027 21675
rect 19334 21672 19340 21684
rect 19015 21644 19340 21672
rect 19015 21641 19027 21644
rect 18969 21635 19027 21641
rect 19334 21632 19340 21644
rect 19392 21632 19398 21684
rect 22373 21675 22431 21681
rect 22373 21641 22385 21675
rect 22419 21672 22431 21675
rect 23474 21672 23480 21684
rect 22419 21644 23480 21672
rect 22419 21641 22431 21644
rect 22373 21635 22431 21641
rect 23474 21632 23480 21644
rect 23532 21632 23538 21684
rect 23658 21672 23664 21684
rect 23619 21644 23664 21672
rect 23658 21632 23664 21644
rect 23716 21632 23722 21684
rect 25317 21675 25375 21681
rect 25317 21641 25329 21675
rect 25363 21672 25375 21675
rect 25682 21672 25688 21684
rect 25363 21644 25688 21672
rect 25363 21641 25375 21644
rect 25317 21635 25375 21641
rect 25682 21632 25688 21644
rect 25740 21632 25746 21684
rect 3050 21536 3056 21548
rect 3011 21508 3056 21536
rect 3050 21496 3056 21508
rect 3108 21496 3114 21548
rect 18782 21536 18788 21548
rect 18695 21508 18788 21536
rect 18782 21496 18788 21508
rect 18840 21536 18846 21548
rect 19242 21536 19248 21548
rect 18840 21508 19248 21536
rect 18840 21496 18846 21508
rect 19242 21496 19248 21508
rect 19300 21496 19306 21548
rect 19702 21496 19708 21548
rect 19760 21536 19766 21548
rect 19889 21539 19947 21545
rect 19889 21536 19901 21539
rect 19760 21508 19901 21536
rect 19760 21496 19766 21508
rect 19889 21505 19901 21508
rect 19935 21505 19947 21539
rect 19889 21499 19947 21505
rect 20346 21496 20352 21548
rect 20404 21536 20410 21548
rect 22189 21539 22247 21545
rect 22189 21536 22201 21539
rect 20404 21508 22201 21536
rect 20404 21496 20410 21508
rect 22189 21505 22201 21508
rect 22235 21505 22247 21539
rect 23474 21536 23480 21548
rect 23435 21508 23480 21536
rect 22189 21499 22247 21505
rect 23474 21496 23480 21508
rect 23532 21496 23538 21548
rect 25130 21536 25136 21548
rect 25091 21508 25136 21536
rect 25130 21496 25136 21508
rect 25188 21536 25194 21548
rect 30926 21536 30932 21548
rect 25188 21508 30932 21536
rect 25188 21496 25194 21508
rect 30926 21496 30932 21508
rect 30984 21496 30990 21548
rect 34057 21539 34115 21545
rect 34057 21505 34069 21539
rect 34103 21536 34115 21539
rect 34514 21536 34520 21548
rect 34103 21508 34520 21536
rect 34103 21505 34115 21508
rect 34057 21499 34115 21505
rect 34514 21496 34520 21508
rect 34572 21496 34578 21548
rect 34701 21539 34759 21545
rect 34701 21505 34713 21539
rect 34747 21505 34759 21539
rect 34701 21499 34759 21505
rect 23293 21471 23351 21477
rect 23293 21437 23305 21471
rect 23339 21468 23351 21471
rect 23382 21468 23388 21480
rect 23339 21440 23388 21468
rect 23339 21437 23351 21440
rect 23293 21431 23351 21437
rect 23382 21428 23388 21440
rect 23440 21468 23446 21480
rect 24949 21471 25007 21477
rect 24949 21468 24961 21471
rect 23440 21440 24961 21468
rect 23440 21428 23446 21440
rect 24949 21437 24961 21440
rect 24995 21437 25007 21471
rect 24949 21431 25007 21437
rect 34422 21428 34428 21480
rect 34480 21468 34486 21480
rect 34716 21468 34744 21499
rect 34480 21440 34744 21468
rect 34480 21428 34486 21440
rect 2869 21335 2927 21341
rect 2869 21301 2881 21335
rect 2915 21332 2927 21335
rect 2958 21332 2964 21344
rect 2915 21304 2964 21332
rect 2915 21301 2927 21304
rect 2869 21295 2927 21301
rect 2958 21292 2964 21304
rect 3016 21292 3022 21344
rect 20073 21335 20131 21341
rect 20073 21301 20085 21335
rect 20119 21332 20131 21335
rect 20254 21332 20260 21344
rect 20119 21304 20260 21332
rect 20119 21301 20131 21304
rect 20073 21295 20131 21301
rect 20254 21292 20260 21304
rect 20312 21292 20318 21344
rect 34885 21335 34943 21341
rect 34885 21301 34897 21335
rect 34931 21332 34943 21335
rect 35986 21332 35992 21344
rect 34931 21304 35992 21332
rect 34931 21301 34943 21304
rect 34885 21295 34943 21301
rect 35986 21292 35992 21304
rect 36044 21292 36050 21344
rect 1104 21242 38824 21264
rect 1104 21190 5674 21242
rect 5726 21190 5738 21242
rect 5790 21190 5802 21242
rect 5854 21190 5866 21242
rect 5918 21190 5930 21242
rect 5982 21190 15122 21242
rect 15174 21190 15186 21242
rect 15238 21190 15250 21242
rect 15302 21190 15314 21242
rect 15366 21190 15378 21242
rect 15430 21190 24570 21242
rect 24622 21190 24634 21242
rect 24686 21190 24698 21242
rect 24750 21190 24762 21242
rect 24814 21190 24826 21242
rect 24878 21190 34018 21242
rect 34070 21190 34082 21242
rect 34134 21190 34146 21242
rect 34198 21190 34210 21242
rect 34262 21190 34274 21242
rect 34326 21190 38824 21242
rect 1104 21168 38824 21190
rect 20898 21128 20904 21140
rect 1688 21100 16574 21128
rect 1688 20933 1716 21100
rect 1673 20927 1731 20933
rect 1673 20893 1685 20927
rect 1719 20924 1731 20927
rect 1762 20924 1768 20936
rect 1719 20896 1768 20924
rect 1719 20893 1731 20896
rect 1673 20887 1731 20893
rect 1762 20884 1768 20896
rect 1820 20884 1826 20936
rect 2958 20924 2964 20936
rect 2919 20896 2964 20924
rect 2958 20884 2964 20896
rect 3016 20884 3022 20936
rect 3237 20927 3295 20933
rect 3237 20893 3249 20927
rect 3283 20924 3295 20927
rect 3878 20924 3884 20936
rect 3283 20896 3884 20924
rect 3283 20893 3295 20896
rect 3237 20887 3295 20893
rect 3878 20884 3884 20896
rect 3936 20884 3942 20936
rect 5994 20924 6000 20936
rect 5955 20896 6000 20924
rect 5994 20884 6000 20896
rect 6052 20884 6058 20936
rect 6273 20927 6331 20933
rect 6273 20893 6285 20927
rect 6319 20924 6331 20927
rect 6638 20924 6644 20936
rect 6319 20896 6644 20924
rect 6319 20893 6331 20896
rect 6273 20887 6331 20893
rect 3896 20856 3924 20884
rect 6288 20856 6316 20887
rect 6638 20884 6644 20896
rect 6696 20924 6702 20936
rect 6733 20927 6791 20933
rect 6733 20924 6745 20927
rect 6696 20896 6745 20924
rect 6696 20884 6702 20896
rect 6733 20893 6745 20896
rect 6779 20893 6791 20927
rect 7006 20924 7012 20936
rect 6967 20896 7012 20924
rect 6733 20887 6791 20893
rect 7006 20884 7012 20896
rect 7064 20884 7070 20936
rect 3896 20828 6316 20856
rect 16546 20856 16574 21100
rect 19996 21100 20904 21128
rect 19996 21001 20024 21100
rect 20898 21088 20904 21100
rect 20956 21088 20962 21140
rect 19981 20995 20039 21001
rect 19981 20961 19993 20995
rect 20027 20961 20039 20995
rect 19981 20955 20039 20961
rect 20254 20924 20260 20936
rect 20215 20896 20260 20924
rect 20254 20884 20260 20896
rect 20312 20884 20318 20936
rect 29730 20924 29736 20936
rect 29691 20896 29736 20924
rect 29730 20884 29736 20896
rect 29788 20884 29794 20936
rect 30466 20884 30472 20936
rect 30524 20924 30530 20936
rect 30561 20927 30619 20933
rect 30561 20924 30573 20927
rect 30524 20896 30573 20924
rect 30524 20884 30530 20896
rect 30561 20893 30573 20896
rect 30607 20893 30619 20927
rect 35986 20924 35992 20936
rect 35947 20896 35992 20924
rect 30561 20887 30619 20893
rect 35986 20884 35992 20896
rect 36044 20884 36050 20936
rect 25406 20856 25412 20868
rect 16546 20828 25412 20856
rect 25406 20816 25412 20828
rect 25464 20816 25470 20868
rect 1486 20788 1492 20800
rect 1447 20760 1492 20788
rect 1486 20748 1492 20760
rect 1544 20748 1550 20800
rect 2222 20788 2228 20800
rect 2183 20760 2228 20788
rect 2222 20748 2228 20760
rect 2280 20788 2286 20800
rect 5261 20791 5319 20797
rect 5261 20788 5273 20791
rect 2280 20760 5273 20788
rect 2280 20748 2286 20760
rect 5261 20757 5273 20760
rect 5307 20788 5319 20791
rect 6730 20788 6736 20800
rect 5307 20760 6736 20788
rect 5307 20757 5319 20760
rect 5261 20751 5319 20757
rect 6730 20748 6736 20760
rect 6788 20788 6794 20800
rect 7745 20791 7803 20797
rect 7745 20788 7757 20791
rect 6788 20760 7757 20788
rect 6788 20748 6794 20760
rect 7745 20757 7757 20760
rect 7791 20757 7803 20791
rect 19242 20788 19248 20800
rect 19203 20760 19248 20788
rect 7745 20751 7803 20757
rect 19242 20748 19248 20760
rect 19300 20748 19306 20800
rect 20990 20788 20996 20800
rect 20951 20760 20996 20788
rect 20990 20748 20996 20760
rect 21048 20748 21054 20800
rect 29914 20788 29920 20800
rect 29875 20760 29920 20788
rect 29914 20748 29920 20760
rect 29972 20748 29978 20800
rect 30374 20788 30380 20800
rect 30335 20760 30380 20788
rect 30374 20748 30380 20760
rect 30432 20748 30438 20800
rect 36173 20791 36231 20797
rect 36173 20757 36185 20791
rect 36219 20788 36231 20791
rect 36906 20788 36912 20800
rect 36219 20760 36912 20788
rect 36219 20757 36231 20760
rect 36173 20751 36231 20757
rect 36906 20748 36912 20760
rect 36964 20748 36970 20800
rect 1104 20698 38824 20720
rect 1104 20646 10398 20698
rect 10450 20646 10462 20698
rect 10514 20646 10526 20698
rect 10578 20646 10590 20698
rect 10642 20646 10654 20698
rect 10706 20646 19846 20698
rect 19898 20646 19910 20698
rect 19962 20646 19974 20698
rect 20026 20646 20038 20698
rect 20090 20646 20102 20698
rect 20154 20646 29294 20698
rect 29346 20646 29358 20698
rect 29410 20646 29422 20698
rect 29474 20646 29486 20698
rect 29538 20646 29550 20698
rect 29602 20646 38824 20698
rect 1104 20624 38824 20646
rect 1762 20584 1768 20596
rect 1723 20556 1768 20584
rect 1762 20544 1768 20556
rect 1820 20544 1826 20596
rect 2774 20544 2780 20596
rect 2832 20584 2838 20596
rect 7745 20587 7803 20593
rect 7745 20584 7757 20587
rect 2832 20556 7757 20584
rect 2832 20544 2838 20556
rect 7745 20553 7757 20556
rect 7791 20584 7803 20587
rect 7791 20556 8340 20584
rect 7791 20553 7803 20556
rect 7745 20547 7803 20553
rect 8312 20525 8340 20556
rect 19702 20544 19708 20596
rect 19760 20584 19766 20596
rect 19797 20587 19855 20593
rect 19797 20584 19809 20587
rect 19760 20556 19809 20584
rect 19760 20544 19766 20556
rect 19797 20553 19809 20556
rect 19843 20553 19855 20587
rect 19797 20547 19855 20553
rect 29730 20544 29736 20596
rect 29788 20584 29794 20596
rect 30193 20587 30251 20593
rect 30193 20584 30205 20587
rect 29788 20556 30205 20584
rect 29788 20544 29794 20556
rect 30193 20553 30205 20556
rect 30239 20553 30251 20587
rect 30193 20547 30251 20553
rect 8297 20519 8355 20525
rect 8297 20485 8309 20519
rect 8343 20485 8355 20519
rect 8297 20479 8355 20485
rect 18325 20519 18383 20525
rect 18325 20485 18337 20519
rect 18371 20516 18383 20519
rect 19242 20516 19248 20528
rect 18371 20488 19248 20516
rect 18371 20485 18383 20488
rect 18325 20479 18383 20485
rect 16945 20451 17003 20457
rect 16945 20417 16957 20451
rect 16991 20448 17003 20451
rect 18340 20448 18368 20479
rect 19242 20476 19248 20488
rect 19300 20516 19306 20528
rect 22922 20516 22928 20528
rect 19300 20488 22928 20516
rect 19300 20476 19306 20488
rect 22922 20476 22928 20488
rect 22980 20476 22986 20528
rect 19610 20448 19616 20460
rect 16991 20420 18368 20448
rect 19571 20420 19616 20448
rect 16991 20417 17003 20420
rect 16945 20411 17003 20417
rect 19610 20408 19616 20420
rect 19668 20408 19674 20460
rect 27522 20408 27528 20460
rect 27580 20448 27586 20460
rect 29549 20451 29607 20457
rect 29549 20448 29561 20451
rect 27580 20420 29561 20448
rect 27580 20408 27586 20420
rect 29549 20417 29561 20420
rect 29595 20448 29607 20451
rect 30377 20451 30435 20457
rect 30377 20448 30389 20451
rect 29595 20420 30389 20448
rect 29595 20417 29607 20420
rect 29549 20411 29607 20417
rect 30377 20417 30389 20420
rect 30423 20417 30435 20451
rect 30377 20411 30435 20417
rect 30561 20451 30619 20457
rect 30561 20417 30573 20451
rect 30607 20448 30619 20451
rect 31294 20448 31300 20460
rect 30607 20420 31300 20448
rect 30607 20417 30619 20420
rect 30561 20411 30619 20417
rect 31294 20408 31300 20420
rect 31352 20448 31358 20460
rect 33137 20451 33195 20457
rect 33137 20448 33149 20451
rect 31352 20420 33149 20448
rect 31352 20408 31358 20420
rect 33137 20417 33149 20420
rect 33183 20417 33195 20451
rect 33137 20411 33195 20417
rect 33226 20408 33232 20460
rect 33284 20448 33290 20460
rect 33321 20451 33379 20457
rect 33321 20448 33333 20451
rect 33284 20420 33333 20448
rect 33284 20408 33290 20420
rect 33321 20417 33333 20420
rect 33367 20448 33379 20451
rect 34241 20451 34299 20457
rect 34241 20448 34253 20451
rect 33367 20420 34253 20448
rect 33367 20417 33379 20420
rect 33321 20411 33379 20417
rect 34241 20417 34253 20420
rect 34287 20448 34299 20451
rect 34330 20448 34336 20460
rect 34287 20420 34336 20448
rect 34287 20417 34299 20420
rect 34241 20411 34299 20417
rect 34330 20408 34336 20420
rect 34388 20408 34394 20460
rect 34425 20451 34483 20457
rect 34425 20417 34437 20451
rect 34471 20448 34483 20451
rect 35069 20451 35127 20457
rect 35069 20448 35081 20451
rect 34471 20420 35081 20448
rect 34471 20417 34483 20420
rect 34425 20411 34483 20417
rect 35069 20417 35081 20420
rect 35115 20417 35127 20451
rect 35069 20411 35127 20417
rect 17218 20380 17224 20392
rect 17179 20352 17224 20380
rect 17218 20340 17224 20352
rect 17276 20380 17282 20392
rect 19429 20383 19487 20389
rect 19429 20380 19441 20383
rect 17276 20352 19441 20380
rect 17276 20340 17282 20352
rect 19429 20349 19441 20352
rect 19475 20380 19487 20383
rect 23382 20380 23388 20392
rect 19475 20352 23388 20380
rect 19475 20349 19487 20352
rect 19429 20343 19487 20349
rect 23382 20340 23388 20352
rect 23440 20340 23446 20392
rect 29365 20383 29423 20389
rect 29365 20349 29377 20383
rect 29411 20349 29423 20383
rect 29365 20343 29423 20349
rect 29733 20383 29791 20389
rect 29733 20349 29745 20383
rect 29779 20380 29791 20383
rect 30466 20380 30472 20392
rect 29779 20352 30472 20380
rect 29779 20349 29791 20352
rect 29733 20343 29791 20349
rect 29380 20312 29408 20343
rect 30466 20340 30472 20352
rect 30524 20340 30530 20392
rect 34057 20383 34115 20389
rect 34057 20349 34069 20383
rect 34103 20349 34115 20383
rect 34057 20343 34115 20349
rect 31202 20312 31208 20324
rect 29380 20284 31208 20312
rect 31202 20272 31208 20284
rect 31260 20312 31266 20324
rect 34072 20312 34100 20343
rect 31260 20284 34100 20312
rect 31260 20272 31266 20284
rect 9582 20244 9588 20256
rect 9543 20216 9588 20244
rect 9582 20204 9588 20216
rect 9640 20204 9646 20256
rect 33505 20247 33563 20253
rect 33505 20213 33517 20247
rect 33551 20244 33563 20247
rect 33870 20244 33876 20256
rect 33551 20216 33876 20244
rect 33551 20213 33563 20216
rect 33505 20207 33563 20213
rect 33870 20204 33876 20216
rect 33928 20204 33934 20256
rect 35253 20247 35311 20253
rect 35253 20213 35265 20247
rect 35299 20244 35311 20247
rect 35986 20244 35992 20256
rect 35299 20216 35992 20244
rect 35299 20213 35311 20216
rect 35253 20207 35311 20213
rect 35986 20204 35992 20216
rect 36044 20204 36050 20256
rect 1104 20154 38824 20176
rect 1104 20102 5674 20154
rect 5726 20102 5738 20154
rect 5790 20102 5802 20154
rect 5854 20102 5866 20154
rect 5918 20102 5930 20154
rect 5982 20102 15122 20154
rect 15174 20102 15186 20154
rect 15238 20102 15250 20154
rect 15302 20102 15314 20154
rect 15366 20102 15378 20154
rect 15430 20102 24570 20154
rect 24622 20102 24634 20154
rect 24686 20102 24698 20154
rect 24750 20102 24762 20154
rect 24814 20102 24826 20154
rect 24878 20102 34018 20154
rect 34070 20102 34082 20154
rect 34134 20102 34146 20154
rect 34198 20102 34210 20154
rect 34262 20102 34274 20154
rect 34326 20102 38824 20154
rect 1104 20080 38824 20102
rect 6638 20040 6644 20052
rect 6599 20012 6644 20040
rect 6638 20000 6644 20012
rect 6696 20000 6702 20052
rect 14826 20040 14832 20052
rect 14787 20012 14832 20040
rect 14826 20000 14832 20012
rect 14884 20000 14890 20052
rect 16853 20043 16911 20049
rect 16853 20009 16865 20043
rect 16899 20040 16911 20043
rect 17034 20040 17040 20052
rect 16899 20012 17040 20040
rect 16899 20009 16911 20012
rect 16853 20003 16911 20009
rect 17034 20000 17040 20012
rect 17092 20000 17098 20052
rect 17313 19975 17371 19981
rect 17313 19972 17325 19975
rect 16546 19944 17325 19972
rect 15105 19907 15163 19913
rect 15105 19873 15117 19907
rect 15151 19904 15163 19907
rect 15562 19904 15568 19916
rect 15151 19876 15568 19904
rect 15151 19873 15163 19876
rect 15105 19867 15163 19873
rect 15562 19864 15568 19876
rect 15620 19904 15626 19916
rect 15841 19907 15899 19913
rect 15841 19904 15853 19907
rect 15620 19876 15853 19904
rect 15620 19864 15626 19876
rect 15841 19873 15853 19876
rect 15887 19873 15899 19907
rect 15841 19867 15899 19873
rect 1673 19839 1731 19845
rect 1673 19805 1685 19839
rect 1719 19836 1731 19839
rect 1719 19808 2268 19836
rect 1719 19805 1731 19808
rect 1673 19799 1731 19805
rect 2240 19777 2268 19808
rect 6270 19796 6276 19848
rect 6328 19836 6334 19848
rect 6457 19839 6515 19845
rect 6457 19836 6469 19839
rect 6328 19808 6469 19836
rect 6328 19796 6334 19808
rect 6457 19805 6469 19808
rect 6503 19805 6515 19839
rect 6457 19799 6515 19805
rect 9674 19796 9680 19848
rect 9732 19836 9738 19848
rect 15197 19839 15255 19845
rect 15197 19836 15209 19839
rect 9732 19808 15209 19836
rect 9732 19796 9738 19808
rect 15197 19805 15209 19808
rect 15243 19805 15255 19839
rect 15197 19799 15255 19805
rect 16117 19839 16175 19845
rect 16117 19805 16129 19839
rect 16163 19836 16175 19839
rect 16546 19836 16574 19944
rect 17313 19941 17325 19944
rect 17359 19941 17371 19975
rect 17313 19935 17371 19941
rect 20530 19864 20536 19916
rect 20588 19904 20594 19916
rect 20625 19907 20683 19913
rect 20625 19904 20637 19907
rect 20588 19876 20637 19904
rect 20588 19864 20594 19876
rect 20625 19873 20637 19876
rect 20671 19904 20683 19907
rect 21085 19907 21143 19913
rect 21085 19904 21097 19907
rect 20671 19876 21097 19904
rect 20671 19873 20683 19876
rect 20625 19867 20683 19873
rect 21085 19873 21097 19876
rect 21131 19873 21143 19907
rect 21085 19867 21143 19873
rect 16163 19808 16574 19836
rect 16163 19805 16175 19808
rect 16117 19799 16175 19805
rect 17034 19796 17040 19848
rect 17092 19836 17098 19848
rect 17497 19839 17555 19845
rect 17497 19836 17509 19839
rect 17092 19808 17509 19836
rect 17092 19796 17098 19808
rect 17497 19805 17509 19808
rect 17543 19805 17555 19839
rect 17497 19799 17555 19805
rect 21269 19839 21327 19845
rect 21269 19805 21281 19839
rect 21315 19805 21327 19839
rect 21269 19799 21327 19805
rect 2225 19771 2283 19777
rect 2225 19737 2237 19771
rect 2271 19768 2283 19771
rect 11698 19768 11704 19780
rect 2271 19740 11704 19768
rect 2271 19737 2283 19740
rect 2225 19731 2283 19737
rect 11698 19728 11704 19740
rect 11756 19728 11762 19780
rect 14550 19728 14556 19780
rect 14608 19768 14614 19780
rect 14737 19771 14795 19777
rect 14737 19768 14749 19771
rect 14608 19740 14749 19768
rect 14608 19728 14614 19740
rect 14737 19737 14749 19740
rect 14783 19737 14795 19771
rect 20346 19768 20352 19780
rect 14737 19731 14795 19737
rect 16546 19740 20352 19768
rect 1486 19700 1492 19712
rect 1447 19672 1492 19700
rect 1486 19660 1492 19672
rect 1544 19660 1550 19712
rect 15381 19703 15439 19709
rect 15381 19669 15393 19703
rect 15427 19700 15439 19703
rect 16546 19700 16574 19740
rect 20346 19728 20352 19740
rect 20404 19728 20410 19780
rect 21284 19768 21312 19799
rect 28902 19796 28908 19848
rect 28960 19836 28966 19848
rect 29641 19839 29699 19845
rect 29641 19836 29653 19839
rect 28960 19808 29653 19836
rect 28960 19796 28966 19808
rect 29641 19805 29653 19808
rect 29687 19805 29699 19839
rect 29914 19836 29920 19848
rect 29875 19808 29920 19836
rect 29641 19799 29699 19805
rect 29914 19796 29920 19808
rect 29972 19796 29978 19848
rect 33870 19836 33876 19848
rect 33831 19808 33876 19836
rect 33870 19796 33876 19808
rect 33928 19796 33934 19848
rect 35713 19839 35771 19845
rect 35713 19805 35725 19839
rect 35759 19836 35771 19839
rect 35986 19836 35992 19848
rect 35759 19808 35894 19836
rect 35947 19808 35992 19836
rect 35759 19805 35771 19808
rect 35713 19799 35771 19805
rect 35866 19780 35894 19808
rect 35986 19796 35992 19808
rect 36044 19796 36050 19848
rect 25038 19768 25044 19780
rect 21284 19740 25044 19768
rect 25038 19728 25044 19740
rect 25096 19768 25102 19780
rect 27522 19768 27528 19780
rect 25096 19740 27528 19768
rect 25096 19728 25102 19740
rect 27522 19728 27528 19740
rect 27580 19728 27586 19780
rect 35866 19740 35900 19780
rect 35894 19728 35900 19740
rect 35952 19728 35958 19780
rect 15427 19672 16574 19700
rect 21453 19703 21511 19709
rect 15427 19669 15439 19672
rect 15381 19663 15439 19669
rect 21453 19669 21465 19703
rect 21499 19700 21511 19703
rect 22002 19700 22008 19712
rect 21499 19672 22008 19700
rect 21499 19669 21511 19672
rect 21453 19663 21511 19669
rect 22002 19660 22008 19672
rect 22060 19660 22066 19712
rect 30466 19660 30472 19712
rect 30524 19700 30530 19712
rect 30653 19703 30711 19709
rect 30653 19700 30665 19703
rect 30524 19672 30665 19700
rect 30524 19660 30530 19672
rect 30653 19669 30665 19672
rect 30699 19669 30711 19703
rect 30653 19663 30711 19669
rect 34057 19703 34115 19709
rect 34057 19669 34069 19703
rect 34103 19700 34115 19703
rect 34698 19700 34704 19712
rect 34103 19672 34704 19700
rect 34103 19669 34115 19672
rect 34057 19663 34115 19669
rect 34698 19660 34704 19672
rect 34756 19660 34762 19712
rect 36725 19703 36783 19709
rect 36725 19669 36737 19703
rect 36771 19700 36783 19703
rect 37458 19700 37464 19712
rect 36771 19672 37464 19700
rect 36771 19669 36783 19672
rect 36725 19663 36783 19669
rect 37458 19660 37464 19672
rect 37516 19660 37522 19712
rect 1104 19610 38824 19632
rect 1104 19558 10398 19610
rect 10450 19558 10462 19610
rect 10514 19558 10526 19610
rect 10578 19558 10590 19610
rect 10642 19558 10654 19610
rect 10706 19558 19846 19610
rect 19898 19558 19910 19610
rect 19962 19558 19974 19610
rect 20026 19558 20038 19610
rect 20090 19558 20102 19610
rect 20154 19558 29294 19610
rect 29346 19558 29358 19610
rect 29410 19558 29422 19610
rect 29474 19558 29486 19610
rect 29538 19558 29550 19610
rect 29602 19558 38824 19610
rect 1104 19536 38824 19558
rect 11698 19456 11704 19508
rect 11756 19496 11762 19508
rect 17034 19496 17040 19508
rect 11756 19468 16896 19496
rect 16995 19468 17040 19496
rect 11756 19456 11762 19468
rect 10689 19431 10747 19437
rect 10689 19428 10701 19431
rect 10060 19400 10701 19428
rect 3421 19363 3479 19369
rect 3421 19329 3433 19363
rect 3467 19360 3479 19363
rect 4614 19360 4620 19372
rect 3467 19332 4620 19360
rect 3467 19329 3479 19332
rect 3421 19323 3479 19329
rect 4614 19320 4620 19332
rect 4672 19320 4678 19372
rect 7098 19360 7104 19372
rect 7059 19332 7104 19360
rect 7098 19320 7104 19332
rect 7156 19320 7162 19372
rect 9398 19320 9404 19372
rect 9456 19360 9462 19372
rect 10060 19369 10088 19400
rect 10689 19397 10701 19400
rect 10735 19397 10747 19431
rect 16868 19428 16896 19468
rect 17034 19456 17040 19468
rect 17092 19456 17098 19508
rect 25501 19499 25559 19505
rect 17144 19468 22094 19496
rect 17144 19428 17172 19468
rect 16868 19400 17172 19428
rect 22066 19428 22094 19468
rect 25501 19465 25513 19499
rect 25547 19496 25559 19499
rect 28902 19496 28908 19508
rect 25547 19468 28908 19496
rect 25547 19465 25559 19468
rect 25501 19459 25559 19465
rect 28902 19456 28908 19468
rect 28960 19456 28966 19508
rect 30466 19456 30472 19508
rect 30524 19496 30530 19508
rect 30653 19499 30711 19505
rect 30653 19496 30665 19499
rect 30524 19468 30665 19496
rect 30524 19456 30530 19468
rect 30653 19465 30665 19468
rect 30699 19465 30711 19499
rect 30653 19459 30711 19465
rect 33965 19499 34023 19505
rect 33965 19465 33977 19499
rect 34011 19496 34023 19499
rect 37458 19496 37464 19508
rect 34011 19468 37464 19496
rect 34011 19465 34023 19468
rect 33965 19459 34023 19465
rect 33980 19428 34008 19459
rect 37458 19456 37464 19468
rect 37516 19456 37522 19508
rect 22066 19400 34008 19428
rect 10689 19391 10747 19397
rect 10045 19363 10103 19369
rect 10045 19360 10057 19363
rect 9456 19332 10057 19360
rect 9456 19320 9462 19332
rect 10045 19329 10057 19332
rect 10091 19329 10103 19363
rect 10045 19323 10103 19329
rect 10137 19363 10195 19369
rect 10137 19329 10149 19363
rect 10183 19360 10195 19363
rect 11330 19360 11336 19372
rect 10183 19332 11336 19360
rect 10183 19329 10195 19332
rect 10137 19323 10195 19329
rect 11330 19320 11336 19332
rect 11388 19320 11394 19372
rect 14826 19320 14832 19372
rect 14884 19360 14890 19372
rect 16853 19363 16911 19369
rect 16853 19360 16865 19363
rect 14884 19332 16865 19360
rect 14884 19320 14890 19332
rect 16853 19329 16865 19332
rect 16899 19329 16911 19363
rect 22002 19360 22008 19372
rect 21963 19332 22008 19360
rect 16853 19323 16911 19329
rect 22002 19320 22008 19332
rect 22060 19320 22066 19372
rect 25317 19363 25375 19369
rect 25317 19329 25329 19363
rect 25363 19360 25375 19363
rect 25958 19360 25964 19372
rect 25363 19332 25820 19360
rect 25919 19332 25964 19360
rect 25363 19329 25375 19332
rect 25317 19323 25375 19329
rect 3237 19295 3295 19301
rect 3237 19261 3249 19295
rect 3283 19292 3295 19295
rect 4065 19295 4123 19301
rect 4065 19292 4077 19295
rect 3283 19264 4077 19292
rect 3283 19261 3295 19264
rect 3237 19255 3295 19261
rect 4065 19261 4077 19264
rect 4111 19292 4123 19295
rect 4154 19292 4160 19304
rect 4111 19264 4160 19292
rect 4111 19261 4123 19264
rect 4065 19255 4123 19261
rect 4154 19252 4160 19264
rect 4212 19252 4218 19304
rect 16669 19295 16727 19301
rect 16669 19261 16681 19295
rect 16715 19292 16727 19295
rect 17218 19292 17224 19304
rect 16715 19264 17224 19292
rect 16715 19261 16727 19264
rect 16669 19255 16727 19261
rect 17218 19252 17224 19264
rect 17276 19252 17282 19304
rect 25792 19224 25820 19332
rect 25958 19320 25964 19332
rect 26016 19320 26022 19372
rect 28902 19320 28908 19372
rect 28960 19360 28966 19372
rect 29641 19363 29699 19369
rect 29641 19360 29653 19363
rect 28960 19332 29653 19360
rect 28960 19320 28966 19332
rect 29641 19329 29653 19332
rect 29687 19329 29699 19363
rect 29641 19323 29699 19329
rect 29917 19363 29975 19369
rect 29917 19329 29929 19363
rect 29963 19360 29975 19363
rect 30374 19360 30380 19372
rect 29963 19332 30380 19360
rect 29963 19329 29975 19332
rect 29917 19323 29975 19329
rect 30374 19320 30380 19332
rect 30432 19320 30438 19372
rect 34698 19360 34704 19372
rect 34659 19332 34704 19360
rect 34698 19320 34704 19332
rect 34756 19320 34762 19372
rect 34977 19363 35035 19369
rect 34977 19329 34989 19363
rect 35023 19360 35035 19363
rect 35894 19360 35900 19372
rect 35023 19332 35900 19360
rect 35023 19329 35035 19332
rect 34977 19323 35035 19329
rect 35894 19320 35900 19332
rect 35952 19360 35958 19372
rect 36630 19360 36636 19372
rect 35952 19332 36636 19360
rect 35952 19320 35958 19332
rect 36630 19320 36636 19332
rect 36688 19320 36694 19372
rect 26145 19227 26203 19233
rect 26145 19224 26157 19227
rect 25792 19196 26157 19224
rect 26145 19193 26157 19196
rect 26191 19224 26203 19227
rect 26234 19224 26240 19236
rect 26191 19196 26240 19224
rect 26191 19193 26203 19196
rect 26145 19187 26203 19193
rect 26234 19184 26240 19196
rect 26292 19184 26298 19236
rect 3605 19159 3663 19165
rect 3605 19125 3617 19159
rect 3651 19156 3663 19159
rect 3970 19156 3976 19168
rect 3651 19128 3976 19156
rect 3651 19125 3663 19128
rect 3605 19119 3663 19125
rect 3970 19116 3976 19128
rect 4028 19116 4034 19168
rect 6917 19159 6975 19165
rect 6917 19125 6929 19159
rect 6963 19156 6975 19159
rect 7006 19156 7012 19168
rect 6963 19128 7012 19156
rect 6963 19125 6975 19128
rect 6917 19119 6975 19125
rect 7006 19116 7012 19128
rect 7064 19116 7070 19168
rect 21634 19116 21640 19168
rect 21692 19156 21698 19168
rect 21821 19159 21879 19165
rect 21821 19156 21833 19159
rect 21692 19128 21833 19156
rect 21692 19116 21698 19128
rect 21821 19125 21833 19128
rect 21867 19125 21879 19159
rect 21821 19119 21879 19125
rect 1104 19066 38824 19088
rect 1104 19014 5674 19066
rect 5726 19014 5738 19066
rect 5790 19014 5802 19066
rect 5854 19014 5866 19066
rect 5918 19014 5930 19066
rect 5982 19014 15122 19066
rect 15174 19014 15186 19066
rect 15238 19014 15250 19066
rect 15302 19014 15314 19066
rect 15366 19014 15378 19066
rect 15430 19014 24570 19066
rect 24622 19014 24634 19066
rect 24686 19014 24698 19066
rect 24750 19014 24762 19066
rect 24814 19014 24826 19066
rect 24878 19014 34018 19066
rect 34070 19014 34082 19066
rect 34134 19014 34146 19066
rect 34198 19014 34210 19066
rect 34262 19014 34274 19066
rect 34326 19014 38824 19066
rect 1104 18992 38824 19014
rect 6730 18912 6736 18964
rect 6788 18952 6794 18964
rect 7377 18955 7435 18961
rect 7377 18952 7389 18955
rect 6788 18924 7389 18952
rect 6788 18912 6794 18924
rect 7377 18921 7389 18924
rect 7423 18921 7435 18955
rect 10042 18952 10048 18964
rect 10003 18924 10048 18952
rect 7377 18915 7435 18921
rect 10042 18912 10048 18924
rect 10100 18912 10106 18964
rect 20898 18952 20904 18964
rect 20811 18924 20904 18952
rect 20898 18912 20904 18924
rect 20956 18952 20962 18964
rect 26237 18955 26295 18961
rect 26237 18952 26249 18955
rect 20956 18924 26249 18952
rect 20956 18912 20962 18924
rect 26237 18921 26249 18924
rect 26283 18952 26295 18955
rect 29822 18952 29828 18964
rect 26283 18924 29828 18952
rect 26283 18921 26295 18924
rect 26237 18915 26295 18921
rect 29822 18912 29828 18924
rect 29880 18952 29886 18964
rect 30466 18952 30472 18964
rect 29880 18924 30472 18952
rect 29880 18912 29886 18924
rect 30466 18912 30472 18924
rect 30524 18912 30530 18964
rect 9490 18776 9496 18828
rect 9548 18816 9554 18828
rect 10597 18819 10655 18825
rect 10597 18816 10609 18819
rect 9548 18788 10609 18816
rect 9548 18776 9554 18788
rect 10597 18785 10609 18788
rect 10643 18785 10655 18819
rect 10597 18779 10655 18785
rect 23382 18776 23388 18828
rect 23440 18816 23446 18828
rect 24397 18819 24455 18825
rect 24397 18816 24409 18819
rect 23440 18788 24409 18816
rect 23440 18776 23446 18788
rect 24397 18785 24409 18788
rect 24443 18785 24455 18819
rect 24397 18779 24455 18785
rect 3970 18748 3976 18760
rect 3931 18720 3976 18748
rect 3970 18708 3976 18720
rect 4028 18708 4034 18760
rect 6270 18708 6276 18760
rect 6328 18748 6334 18760
rect 6365 18751 6423 18757
rect 6365 18748 6377 18751
rect 6328 18720 6377 18748
rect 6328 18708 6334 18720
rect 6365 18717 6377 18720
rect 6411 18717 6423 18751
rect 6365 18711 6423 18717
rect 6641 18751 6699 18757
rect 6641 18717 6653 18751
rect 6687 18748 6699 18751
rect 7006 18748 7012 18760
rect 6687 18720 7012 18748
rect 6687 18717 6699 18720
rect 6641 18711 6699 18717
rect 7006 18708 7012 18720
rect 7064 18708 7070 18760
rect 9858 18748 9864 18760
rect 9819 18720 9864 18748
rect 9858 18708 9864 18720
rect 9916 18708 9922 18760
rect 21634 18748 21640 18760
rect 21595 18720 21640 18748
rect 21634 18708 21640 18720
rect 21692 18708 21698 18760
rect 21913 18751 21971 18757
rect 21913 18717 21925 18751
rect 21959 18717 21971 18751
rect 21913 18711 21971 18717
rect 10873 18683 10931 18689
rect 10873 18649 10885 18683
rect 10919 18680 10931 18683
rect 11146 18680 11152 18692
rect 10919 18652 11152 18680
rect 10919 18649 10931 18652
rect 10873 18643 10931 18649
rect 11146 18640 11152 18652
rect 11204 18640 11210 18692
rect 11330 18640 11336 18692
rect 11388 18640 11394 18692
rect 20622 18640 20628 18692
rect 20680 18680 20686 18692
rect 21928 18680 21956 18711
rect 24486 18708 24492 18760
rect 24544 18748 24550 18760
rect 24581 18751 24639 18757
rect 24581 18748 24593 18751
rect 24544 18720 24593 18748
rect 24544 18708 24550 18720
rect 24581 18717 24593 18720
rect 24627 18717 24639 18751
rect 24581 18711 24639 18717
rect 25225 18751 25283 18757
rect 25225 18717 25237 18751
rect 25271 18717 25283 18751
rect 25225 18711 25283 18717
rect 25240 18680 25268 18711
rect 25406 18708 25412 18760
rect 25464 18748 25470 18760
rect 25501 18751 25559 18757
rect 25501 18748 25513 18751
rect 25464 18720 25513 18748
rect 25464 18708 25470 18720
rect 25501 18717 25513 18720
rect 25547 18717 25559 18751
rect 36630 18748 36636 18760
rect 36591 18720 36636 18748
rect 25501 18711 25559 18717
rect 36630 18708 36636 18720
rect 36688 18708 36694 18760
rect 36906 18748 36912 18760
rect 36867 18720 36912 18748
rect 36906 18708 36912 18720
rect 36964 18708 36970 18760
rect 25958 18680 25964 18692
rect 20680 18652 25964 18680
rect 20680 18640 20686 18652
rect 25958 18640 25964 18652
rect 26016 18640 26022 18692
rect 3602 18572 3608 18624
rect 3660 18612 3666 18624
rect 3789 18615 3847 18621
rect 3789 18612 3801 18615
rect 3660 18584 3801 18612
rect 3660 18572 3666 18584
rect 3789 18581 3801 18584
rect 3835 18581 3847 18615
rect 3789 18575 3847 18581
rect 12250 18572 12256 18624
rect 12308 18612 12314 18624
rect 12345 18615 12403 18621
rect 12345 18612 12357 18615
rect 12308 18584 12357 18612
rect 12308 18572 12314 18584
rect 12345 18581 12357 18584
rect 12391 18581 12403 18615
rect 12345 18575 12403 18581
rect 24765 18615 24823 18621
rect 24765 18581 24777 18615
rect 24811 18612 24823 18615
rect 25222 18612 25228 18624
rect 24811 18584 25228 18612
rect 24811 18581 24823 18584
rect 24765 18575 24823 18581
rect 25222 18572 25228 18584
rect 25280 18572 25286 18624
rect 37458 18572 37464 18624
rect 37516 18612 37522 18624
rect 37645 18615 37703 18621
rect 37645 18612 37657 18615
rect 37516 18584 37657 18612
rect 37516 18572 37522 18584
rect 37645 18581 37657 18584
rect 37691 18581 37703 18615
rect 37645 18575 37703 18581
rect 1104 18522 38824 18544
rect 1104 18470 10398 18522
rect 10450 18470 10462 18522
rect 10514 18470 10526 18522
rect 10578 18470 10590 18522
rect 10642 18470 10654 18522
rect 10706 18470 19846 18522
rect 19898 18470 19910 18522
rect 19962 18470 19974 18522
rect 20026 18470 20038 18522
rect 20090 18470 20102 18522
rect 20154 18470 29294 18522
rect 29346 18470 29358 18522
rect 29410 18470 29422 18522
rect 29474 18470 29486 18522
rect 29538 18470 29550 18522
rect 29602 18470 38824 18522
rect 1104 18448 38824 18470
rect 6917 18411 6975 18417
rect 6917 18377 6929 18411
rect 6963 18408 6975 18411
rect 7098 18408 7104 18420
rect 6963 18380 7104 18408
rect 6963 18377 6975 18380
rect 6917 18371 6975 18377
rect 7098 18368 7104 18380
rect 7156 18368 7162 18420
rect 12894 18368 12900 18420
rect 12952 18408 12958 18420
rect 12989 18411 13047 18417
rect 12989 18408 13001 18411
rect 12952 18380 13001 18408
rect 12952 18368 12958 18380
rect 12989 18377 13001 18380
rect 13035 18377 13047 18411
rect 25406 18408 25412 18420
rect 25367 18380 25412 18408
rect 12989 18371 13047 18377
rect 25406 18368 25412 18380
rect 25464 18368 25470 18420
rect 7837 18343 7895 18349
rect 7837 18309 7849 18343
rect 7883 18340 7895 18343
rect 8294 18340 8300 18352
rect 7883 18312 8300 18340
rect 7883 18309 7895 18312
rect 7837 18303 7895 18309
rect 8294 18300 8300 18312
rect 8352 18340 8358 18352
rect 9582 18340 9588 18352
rect 8352 18312 9588 18340
rect 8352 18300 8358 18312
rect 9582 18300 9588 18312
rect 9640 18300 9646 18352
rect 11146 18300 11152 18352
rect 11204 18340 11210 18352
rect 14093 18343 14151 18349
rect 14093 18340 14105 18343
rect 11204 18312 14105 18340
rect 11204 18300 11210 18312
rect 14093 18309 14105 18312
rect 14139 18309 14151 18343
rect 14093 18303 14151 18309
rect 1673 18275 1731 18281
rect 1673 18241 1685 18275
rect 1719 18272 1731 18275
rect 1946 18272 1952 18284
rect 1719 18244 1952 18272
rect 1719 18241 1731 18244
rect 1673 18235 1731 18241
rect 1946 18232 1952 18244
rect 2004 18232 2010 18284
rect 3602 18272 3608 18284
rect 3563 18244 3608 18272
rect 3602 18232 3608 18244
rect 3660 18232 3666 18284
rect 3878 18272 3884 18284
rect 3839 18244 3884 18272
rect 3878 18232 3884 18244
rect 3936 18232 3942 18284
rect 7101 18275 7159 18281
rect 7101 18272 7113 18275
rect 6886 18244 7113 18272
rect 4614 18164 4620 18216
rect 4672 18204 4678 18216
rect 6886 18204 6914 18244
rect 7101 18241 7113 18244
rect 7147 18241 7159 18275
rect 7101 18235 7159 18241
rect 13633 18275 13691 18281
rect 13633 18241 13645 18275
rect 13679 18272 13691 18275
rect 14366 18272 14372 18284
rect 13679 18244 14372 18272
rect 13679 18241 13691 18244
rect 13633 18235 13691 18241
rect 14366 18232 14372 18244
rect 14424 18232 14430 18284
rect 14550 18232 14556 18284
rect 14608 18272 14614 18284
rect 25222 18272 25228 18284
rect 14608 18244 14653 18272
rect 25183 18244 25228 18272
rect 14608 18232 14614 18244
rect 25222 18232 25228 18244
rect 25280 18232 25286 18284
rect 7282 18204 7288 18216
rect 4672 18176 6914 18204
rect 7243 18176 7288 18204
rect 4672 18164 4678 18176
rect 7282 18164 7288 18176
rect 7340 18164 7346 18216
rect 9122 18164 9128 18216
rect 9180 18204 9186 18216
rect 9585 18207 9643 18213
rect 9585 18204 9597 18207
rect 9180 18176 9597 18204
rect 9180 18164 9186 18176
rect 9585 18173 9597 18176
rect 9631 18204 9643 18207
rect 10870 18204 10876 18216
rect 9631 18176 10876 18204
rect 9631 18173 9643 18176
rect 9585 18167 9643 18173
rect 10870 18164 10876 18176
rect 10928 18164 10934 18216
rect 12894 18164 12900 18216
rect 12952 18204 12958 18216
rect 13262 18204 13268 18216
rect 12952 18176 13268 18204
rect 12952 18164 12958 18176
rect 13262 18164 13268 18176
rect 13320 18204 13326 18216
rect 14185 18207 14243 18213
rect 14185 18204 14197 18207
rect 13320 18176 14197 18204
rect 13320 18164 13326 18176
rect 14185 18173 14197 18176
rect 14231 18173 14243 18207
rect 14185 18167 14243 18173
rect 1486 18068 1492 18080
rect 1447 18040 1492 18068
rect 1486 18028 1492 18040
rect 1544 18028 1550 18080
rect 1946 18028 1952 18080
rect 2004 18068 2010 18080
rect 2133 18071 2191 18077
rect 2133 18068 2145 18071
rect 2004 18040 2145 18068
rect 2004 18028 2010 18040
rect 2133 18037 2145 18040
rect 2179 18037 2191 18071
rect 2133 18031 2191 18037
rect 2222 18028 2228 18080
rect 2280 18068 2286 18080
rect 2869 18071 2927 18077
rect 2869 18068 2881 18071
rect 2280 18040 2881 18068
rect 2280 18028 2286 18040
rect 2869 18037 2881 18040
rect 2915 18037 2927 18071
rect 14274 18068 14280 18080
rect 14235 18040 14280 18068
rect 2869 18031 2927 18037
rect 14274 18028 14280 18040
rect 14332 18028 14338 18080
rect 1104 17978 38824 18000
rect 1104 17926 5674 17978
rect 5726 17926 5738 17978
rect 5790 17926 5802 17978
rect 5854 17926 5866 17978
rect 5918 17926 5930 17978
rect 5982 17926 15122 17978
rect 15174 17926 15186 17978
rect 15238 17926 15250 17978
rect 15302 17926 15314 17978
rect 15366 17926 15378 17978
rect 15430 17926 24570 17978
rect 24622 17926 24634 17978
rect 24686 17926 24698 17978
rect 24750 17926 24762 17978
rect 24814 17926 24826 17978
rect 24878 17926 34018 17978
rect 34070 17926 34082 17978
rect 34134 17926 34146 17978
rect 34198 17926 34210 17978
rect 34262 17926 34274 17978
rect 34326 17926 38824 17978
rect 1104 17904 38824 17926
rect 9309 17867 9367 17873
rect 9309 17833 9321 17867
rect 9355 17864 9367 17867
rect 9858 17864 9864 17876
rect 9355 17836 9864 17864
rect 9355 17833 9367 17836
rect 9309 17827 9367 17833
rect 9858 17824 9864 17836
rect 9916 17824 9922 17876
rect 14274 17824 14280 17876
rect 14332 17864 14338 17876
rect 14737 17867 14795 17873
rect 14737 17864 14749 17867
rect 14332 17836 14749 17864
rect 14332 17824 14338 17836
rect 14737 17833 14749 17836
rect 14783 17833 14795 17867
rect 14737 17827 14795 17833
rect 4614 17728 4620 17740
rect 4575 17700 4620 17728
rect 4614 17688 4620 17700
rect 4672 17688 4678 17740
rect 15381 17731 15439 17737
rect 15381 17728 15393 17731
rect 14752 17700 15393 17728
rect 14752 17672 14780 17700
rect 15381 17697 15393 17700
rect 15427 17697 15439 17731
rect 15381 17691 15439 17697
rect 24688 17700 27108 17728
rect 4893 17663 4951 17669
rect 4893 17629 4905 17663
rect 4939 17660 4951 17663
rect 4939 17632 6914 17660
rect 4939 17629 4951 17632
rect 4893 17623 4951 17629
rect 3970 17552 3976 17604
rect 4028 17592 4034 17604
rect 4908 17592 4936 17623
rect 4028 17564 4936 17592
rect 6886 17592 6914 17632
rect 8202 17620 8208 17672
rect 8260 17660 8266 17672
rect 9125 17663 9183 17669
rect 9125 17660 9137 17663
rect 8260 17632 9137 17660
rect 8260 17620 8266 17632
rect 9125 17629 9137 17632
rect 9171 17629 9183 17663
rect 9125 17623 9183 17629
rect 14366 17620 14372 17672
rect 14424 17660 14430 17672
rect 14734 17660 14740 17672
rect 14424 17632 14740 17660
rect 14424 17620 14430 17632
rect 14734 17620 14740 17632
rect 14792 17620 14798 17672
rect 14921 17663 14979 17669
rect 14921 17629 14933 17663
rect 14967 17660 14979 17663
rect 15470 17660 15476 17672
rect 14967 17632 15476 17660
rect 14967 17629 14979 17632
rect 14921 17623 14979 17629
rect 15470 17620 15476 17632
rect 15528 17620 15534 17672
rect 23566 17620 23572 17672
rect 23624 17660 23630 17672
rect 24486 17660 24492 17672
rect 23624 17632 24492 17660
rect 23624 17620 23630 17632
rect 24486 17620 24492 17632
rect 24544 17660 24550 17672
rect 24688 17669 24716 17700
rect 24673 17663 24731 17669
rect 24673 17660 24685 17663
rect 24544 17632 24685 17660
rect 24544 17620 24550 17632
rect 24673 17629 24685 17632
rect 24719 17629 24731 17663
rect 24673 17623 24731 17629
rect 24949 17663 25007 17669
rect 24949 17629 24961 17663
rect 24995 17660 25007 17663
rect 25038 17660 25044 17672
rect 24995 17632 25044 17660
rect 24995 17629 25007 17632
rect 24949 17623 25007 17629
rect 25038 17620 25044 17632
rect 25096 17660 25102 17672
rect 26326 17660 26332 17672
rect 25096 17632 26332 17660
rect 25096 17620 25102 17632
rect 26326 17620 26332 17632
rect 26384 17620 26390 17672
rect 26970 17660 26976 17672
rect 26931 17632 26976 17660
rect 26970 17620 26976 17632
rect 27028 17620 27034 17672
rect 27080 17669 27108 17700
rect 27065 17663 27123 17669
rect 27065 17629 27077 17663
rect 27111 17629 27123 17663
rect 27065 17623 27123 17629
rect 27249 17663 27307 17669
rect 27249 17629 27261 17663
rect 27295 17660 27307 17663
rect 28077 17663 28135 17669
rect 28077 17660 28089 17663
rect 27295 17632 28089 17660
rect 27295 17629 27307 17632
rect 27249 17623 27307 17629
rect 28077 17629 28089 17632
rect 28123 17629 28135 17663
rect 28077 17623 28135 17629
rect 8941 17595 8999 17601
rect 8941 17592 8953 17595
rect 6886 17564 8953 17592
rect 4028 17552 4034 17564
rect 8941 17561 8953 17564
rect 8987 17592 8999 17595
rect 10962 17592 10968 17604
rect 8987 17564 10968 17592
rect 8987 17561 8999 17564
rect 8941 17555 8999 17561
rect 10962 17552 10968 17564
rect 11020 17552 11026 17604
rect 17954 17552 17960 17604
rect 18012 17592 18018 17604
rect 19426 17592 19432 17604
rect 18012 17564 19432 17592
rect 18012 17552 18018 17564
rect 19426 17552 19432 17564
rect 19484 17552 19490 17604
rect 7282 17484 7288 17536
rect 7340 17524 7346 17536
rect 7469 17527 7527 17533
rect 7469 17524 7481 17527
rect 7340 17496 7481 17524
rect 7340 17484 7346 17496
rect 7469 17493 7481 17496
rect 7515 17524 7527 17527
rect 8846 17524 8852 17536
rect 7515 17496 8852 17524
rect 7515 17493 7527 17496
rect 7469 17487 7527 17493
rect 8846 17484 8852 17496
rect 8904 17484 8910 17536
rect 17770 17484 17776 17536
rect 17828 17524 17834 17536
rect 22094 17524 22100 17536
rect 17828 17496 22100 17524
rect 17828 17484 17834 17496
rect 22094 17484 22100 17496
rect 22152 17484 22158 17536
rect 28261 17527 28319 17533
rect 28261 17493 28273 17527
rect 28307 17524 28319 17527
rect 29086 17524 29092 17536
rect 28307 17496 29092 17524
rect 28307 17493 28319 17496
rect 28261 17487 28319 17493
rect 29086 17484 29092 17496
rect 29144 17484 29150 17536
rect 1104 17434 38824 17456
rect 1104 17382 10398 17434
rect 10450 17382 10462 17434
rect 10514 17382 10526 17434
rect 10578 17382 10590 17434
rect 10642 17382 10654 17434
rect 10706 17382 19846 17434
rect 19898 17382 19910 17434
rect 19962 17382 19974 17434
rect 20026 17382 20038 17434
rect 20090 17382 20102 17434
rect 20154 17382 29294 17434
rect 29346 17382 29358 17434
rect 29410 17382 29422 17434
rect 29474 17382 29486 17434
rect 29538 17382 29550 17434
rect 29602 17382 38824 17434
rect 1104 17360 38824 17382
rect 13446 17280 13452 17332
rect 13504 17320 13510 17332
rect 17589 17323 17647 17329
rect 17589 17320 17601 17323
rect 13504 17292 17601 17320
rect 13504 17280 13510 17292
rect 17589 17289 17601 17292
rect 17635 17289 17647 17323
rect 17770 17320 17776 17332
rect 17731 17292 17776 17320
rect 17589 17283 17647 17289
rect 17770 17280 17776 17292
rect 17828 17280 17834 17332
rect 18969 17323 19027 17329
rect 18969 17289 18981 17323
rect 19015 17320 19027 17323
rect 19610 17320 19616 17332
rect 19015 17292 19616 17320
rect 19015 17289 19027 17292
rect 18969 17283 19027 17289
rect 19610 17280 19616 17292
rect 19668 17280 19674 17332
rect 22465 17323 22523 17329
rect 22465 17289 22477 17323
rect 22511 17320 22523 17323
rect 25130 17320 25136 17332
rect 22511 17292 25136 17320
rect 22511 17289 22523 17292
rect 22465 17283 22523 17289
rect 25130 17280 25136 17292
rect 25188 17280 25194 17332
rect 26970 17280 26976 17332
rect 27028 17320 27034 17332
rect 27433 17323 27491 17329
rect 27433 17320 27445 17323
rect 27028 17292 27445 17320
rect 27028 17280 27034 17292
rect 27433 17289 27445 17292
rect 27479 17320 27491 17323
rect 30650 17320 30656 17332
rect 27479 17292 30656 17320
rect 27479 17289 27491 17292
rect 27433 17283 27491 17289
rect 30650 17280 30656 17292
rect 30708 17320 30714 17332
rect 30708 17292 32628 17320
rect 30708 17280 30714 17292
rect 18601 17255 18659 17261
rect 18601 17221 18613 17255
rect 18647 17221 18659 17255
rect 18601 17215 18659 17221
rect 18817 17255 18875 17261
rect 18817 17221 18829 17255
rect 18863 17252 18875 17255
rect 19794 17252 19800 17264
rect 18863 17224 19800 17252
rect 18863 17221 18875 17224
rect 18817 17215 18875 17221
rect 1673 17187 1731 17193
rect 1673 17153 1685 17187
rect 1719 17184 1731 17187
rect 2225 17187 2283 17193
rect 2225 17184 2237 17187
rect 1719 17156 2237 17184
rect 1719 17153 1731 17156
rect 1673 17147 1731 17153
rect 2225 17153 2237 17156
rect 2271 17184 2283 17187
rect 17954 17184 17960 17196
rect 2271 17156 17960 17184
rect 2271 17153 2283 17156
rect 2225 17147 2283 17153
rect 17954 17144 17960 17156
rect 18012 17144 18018 17196
rect 18616 17184 18644 17215
rect 19058 17184 19064 17196
rect 18616 17156 19064 17184
rect 19058 17144 19064 17156
rect 19116 17144 19122 17196
rect 19168 17116 19196 17224
rect 19794 17212 19800 17224
rect 19852 17212 19858 17264
rect 22094 17252 22100 17264
rect 22055 17224 22100 17252
rect 22094 17212 22100 17224
rect 22152 17212 22158 17264
rect 22278 17212 22284 17264
rect 22336 17261 22342 17264
rect 22336 17255 22355 17261
rect 22343 17221 22355 17255
rect 22336 17215 22355 17221
rect 22336 17212 22342 17215
rect 28902 17212 28908 17264
rect 28960 17212 28966 17264
rect 28813 17187 28871 17193
rect 28813 17153 28825 17187
rect 28859 17184 28871 17187
rect 28920 17184 28948 17212
rect 29086 17184 29092 17196
rect 28859 17156 28948 17184
rect 29047 17156 29092 17184
rect 28859 17153 28871 17156
rect 28813 17147 28871 17153
rect 29086 17144 29092 17156
rect 29144 17144 29150 17196
rect 32600 17193 32628 17292
rect 32585 17187 32643 17193
rect 32585 17153 32597 17187
rect 32631 17184 32643 17187
rect 33045 17187 33103 17193
rect 33045 17184 33057 17187
rect 32631 17156 33057 17184
rect 32631 17153 32643 17156
rect 32585 17147 32643 17153
rect 33045 17153 33057 17156
rect 33091 17153 33103 17187
rect 33226 17184 33232 17196
rect 33187 17156 33232 17184
rect 33045 17147 33103 17153
rect 33226 17144 33232 17156
rect 33284 17144 33290 17196
rect 35066 17144 35072 17196
rect 35124 17184 35130 17196
rect 35805 17187 35863 17193
rect 35805 17184 35817 17187
rect 35124 17156 35817 17184
rect 35124 17144 35130 17156
rect 35805 17153 35817 17156
rect 35851 17153 35863 17187
rect 35805 17147 35863 17153
rect 17788 17088 19196 17116
rect 17788 16992 17816 17088
rect 18141 17051 18199 17057
rect 18141 17017 18153 17051
rect 18187 17048 18199 17051
rect 29822 17048 29828 17060
rect 18187 17020 18828 17048
rect 29783 17020 29828 17048
rect 18187 17017 18199 17020
rect 18141 17011 18199 17017
rect 18800 16992 18828 17020
rect 29822 17008 29828 17020
rect 29880 17048 29886 17060
rect 30742 17048 30748 17060
rect 29880 17020 30748 17048
rect 29880 17008 29886 17020
rect 30742 17008 30748 17020
rect 30800 17008 30806 17060
rect 1486 16980 1492 16992
rect 1447 16952 1492 16980
rect 1486 16940 1492 16952
rect 1544 16940 1550 16992
rect 17770 16980 17776 16992
rect 17683 16952 17776 16980
rect 17770 16940 17776 16952
rect 17828 16940 17834 16992
rect 18782 16980 18788 16992
rect 18695 16952 18788 16980
rect 18782 16940 18788 16952
rect 18840 16980 18846 16992
rect 21450 16980 21456 16992
rect 18840 16952 21456 16980
rect 18840 16940 18846 16952
rect 21450 16940 21456 16952
rect 21508 16980 21514 16992
rect 22281 16983 22339 16989
rect 22281 16980 22293 16983
rect 21508 16952 22293 16980
rect 21508 16940 21514 16952
rect 22281 16949 22293 16952
rect 22327 16949 22339 16983
rect 33410 16980 33416 16992
rect 33371 16952 33416 16980
rect 22281 16943 22339 16949
rect 33410 16940 33416 16952
rect 33468 16940 33474 16992
rect 35989 16983 36047 16989
rect 35989 16949 36001 16983
rect 36035 16980 36047 16983
rect 36722 16980 36728 16992
rect 36035 16952 36728 16980
rect 36035 16949 36047 16952
rect 35989 16943 36047 16949
rect 36722 16940 36728 16952
rect 36780 16940 36786 16992
rect 1104 16890 38824 16912
rect 1104 16838 5674 16890
rect 5726 16838 5738 16890
rect 5790 16838 5802 16890
rect 5854 16838 5866 16890
rect 5918 16838 5930 16890
rect 5982 16838 15122 16890
rect 15174 16838 15186 16890
rect 15238 16838 15250 16890
rect 15302 16838 15314 16890
rect 15366 16838 15378 16890
rect 15430 16838 24570 16890
rect 24622 16838 24634 16890
rect 24686 16838 24698 16890
rect 24750 16838 24762 16890
rect 24814 16838 24826 16890
rect 24878 16838 34018 16890
rect 34070 16838 34082 16890
rect 34134 16838 34146 16890
rect 34198 16838 34210 16890
rect 34262 16838 34274 16890
rect 34326 16838 38824 16890
rect 1104 16816 38824 16838
rect 4154 16736 4160 16788
rect 4212 16776 4218 16788
rect 4709 16779 4767 16785
rect 4709 16776 4721 16779
rect 4212 16748 4721 16776
rect 4212 16736 4218 16748
rect 4709 16745 4721 16748
rect 4755 16776 4767 16779
rect 9030 16776 9036 16788
rect 4755 16748 9036 16776
rect 4755 16745 4767 16748
rect 4709 16739 4767 16745
rect 9030 16736 9036 16748
rect 9088 16736 9094 16788
rect 9674 16736 9680 16788
rect 9732 16776 9738 16788
rect 11885 16779 11943 16785
rect 11885 16776 11897 16779
rect 9732 16748 11897 16776
rect 9732 16736 9738 16748
rect 11885 16745 11897 16748
rect 11931 16745 11943 16779
rect 11885 16739 11943 16745
rect 21637 16779 21695 16785
rect 21637 16745 21649 16779
rect 21683 16776 21695 16779
rect 23474 16776 23480 16788
rect 21683 16748 23480 16776
rect 21683 16745 21695 16748
rect 21637 16739 21695 16745
rect 23474 16736 23480 16748
rect 23532 16736 23538 16788
rect 35066 16776 35072 16788
rect 35027 16748 35072 16776
rect 35066 16736 35072 16748
rect 35124 16736 35130 16788
rect 1578 16668 1584 16720
rect 1636 16708 1642 16720
rect 2222 16708 2228 16720
rect 1636 16680 2228 16708
rect 1636 16668 1642 16680
rect 2222 16668 2228 16680
rect 2280 16668 2286 16720
rect 6181 16711 6239 16717
rect 6181 16708 6193 16711
rect 3252 16680 6193 16708
rect 3252 16649 3280 16680
rect 6181 16677 6193 16680
rect 6227 16677 6239 16711
rect 6181 16671 6239 16677
rect 3237 16643 3295 16649
rect 3237 16609 3249 16643
rect 3283 16609 3295 16643
rect 3237 16603 3295 16609
rect 2958 16572 2964 16584
rect 2919 16544 2964 16572
rect 2958 16532 2964 16544
rect 3016 16532 3022 16584
rect 3970 16572 3976 16584
rect 3931 16544 3976 16572
rect 3970 16532 3976 16544
rect 4028 16532 4034 16584
rect 4154 16572 4160 16584
rect 4115 16544 4160 16572
rect 4154 16532 4160 16544
rect 4212 16532 4218 16584
rect 6196 16572 6224 16671
rect 9398 16668 9404 16720
rect 9456 16708 9462 16720
rect 9950 16708 9956 16720
rect 9456 16680 9956 16708
rect 9456 16668 9462 16680
rect 9950 16668 9956 16680
rect 10008 16668 10014 16720
rect 16114 16708 16120 16720
rect 16075 16680 16120 16708
rect 16114 16668 16120 16680
rect 16172 16668 16178 16720
rect 22278 16708 22284 16720
rect 20088 16680 22284 16708
rect 6914 16600 6920 16652
rect 6972 16640 6978 16652
rect 8202 16640 8208 16652
rect 6972 16612 8208 16640
rect 6972 16600 6978 16612
rect 8202 16600 8208 16612
rect 8260 16640 8266 16652
rect 9769 16643 9827 16649
rect 9769 16640 9781 16643
rect 8260 16612 9781 16640
rect 8260 16600 8266 16612
rect 9769 16609 9781 16612
rect 9815 16609 9827 16643
rect 9769 16603 9827 16609
rect 11698 16600 11704 16652
rect 11756 16640 11762 16652
rect 12066 16640 12072 16652
rect 11756 16612 12072 16640
rect 11756 16600 11762 16612
rect 12066 16600 12072 16612
rect 12124 16600 12130 16652
rect 19794 16640 19800 16652
rect 19755 16612 19800 16640
rect 19794 16600 19800 16612
rect 19852 16600 19858 16652
rect 20088 16649 20116 16680
rect 22278 16668 22284 16680
rect 22336 16708 22342 16720
rect 36725 16711 36783 16717
rect 22336 16680 22968 16708
rect 22336 16668 22342 16680
rect 20073 16643 20131 16649
rect 20073 16609 20085 16643
rect 20119 16609 20131 16643
rect 21082 16640 21088 16652
rect 21043 16612 21088 16640
rect 20073 16603 20131 16609
rect 21082 16600 21088 16612
rect 21140 16600 21146 16652
rect 22830 16640 22836 16652
rect 22791 16612 22836 16640
rect 22830 16600 22836 16612
rect 22888 16600 22894 16652
rect 22940 16649 22968 16680
rect 36725 16677 36737 16711
rect 36771 16708 36783 16711
rect 37458 16708 37464 16720
rect 36771 16680 37464 16708
rect 36771 16677 36783 16680
rect 36725 16671 36783 16677
rect 37458 16668 37464 16680
rect 37516 16668 37522 16720
rect 22925 16643 22983 16649
rect 22925 16609 22937 16643
rect 22971 16640 22983 16643
rect 23474 16640 23480 16652
rect 22971 16612 23480 16640
rect 22971 16609 22983 16612
rect 22925 16603 22983 16609
rect 23474 16600 23480 16612
rect 23532 16600 23538 16652
rect 33226 16600 33232 16652
rect 33284 16640 33290 16652
rect 33284 16612 34928 16640
rect 33284 16600 33290 16612
rect 6270 16572 6276 16584
rect 6183 16544 6276 16572
rect 6270 16532 6276 16544
rect 6328 16572 6334 16584
rect 7009 16575 7067 16581
rect 7009 16572 7021 16575
rect 6328 16544 7021 16572
rect 6328 16532 6334 16544
rect 7009 16541 7021 16544
rect 7055 16541 7067 16575
rect 7009 16535 7067 16541
rect 9582 16532 9588 16584
rect 9640 16572 9646 16584
rect 9950 16572 9956 16584
rect 9640 16544 9956 16572
rect 9640 16532 9646 16544
rect 9950 16532 9956 16544
rect 10008 16532 10014 16584
rect 10045 16575 10103 16581
rect 10045 16541 10057 16575
rect 10091 16572 10103 16575
rect 10778 16572 10784 16584
rect 10091 16544 10784 16572
rect 10091 16541 10103 16544
rect 10045 16535 10103 16541
rect 10778 16532 10784 16544
rect 10836 16572 10842 16584
rect 12161 16575 12219 16581
rect 12161 16572 12173 16575
rect 10836 16544 12173 16572
rect 10836 16532 10842 16544
rect 12161 16541 12173 16544
rect 12207 16541 12219 16575
rect 12161 16535 12219 16541
rect 14550 16532 14556 16584
rect 14608 16572 14614 16584
rect 22649 16575 22707 16581
rect 14608 16544 22416 16572
rect 14608 16532 14614 16544
rect 6365 16507 6423 16513
rect 6365 16473 6377 16507
rect 6411 16504 6423 16507
rect 6914 16504 6920 16516
rect 6411 16476 6920 16504
rect 6411 16473 6423 16476
rect 6365 16467 6423 16473
rect 6914 16464 6920 16476
rect 6972 16464 6978 16516
rect 10962 16464 10968 16516
rect 11020 16504 11026 16516
rect 11885 16507 11943 16513
rect 11885 16504 11897 16507
rect 11020 16476 11897 16504
rect 11020 16464 11026 16476
rect 11885 16473 11897 16476
rect 11931 16504 11943 16507
rect 14366 16504 14372 16516
rect 11931 16476 14372 16504
rect 11931 16473 11943 16476
rect 11885 16467 11943 16473
rect 14366 16464 14372 16476
rect 14424 16464 14430 16516
rect 15838 16504 15844 16516
rect 15799 16476 15844 16504
rect 15838 16464 15844 16476
rect 15896 16464 15902 16516
rect 21174 16464 21180 16516
rect 21232 16504 21238 16516
rect 21269 16507 21327 16513
rect 21269 16504 21281 16507
rect 21232 16476 21281 16504
rect 21232 16464 21238 16476
rect 21269 16473 21281 16476
rect 21315 16473 21327 16507
rect 21269 16467 21327 16473
rect 21361 16507 21419 16513
rect 21361 16473 21373 16507
rect 21407 16504 21419 16507
rect 22094 16504 22100 16516
rect 21407 16476 22100 16504
rect 21407 16473 21419 16476
rect 21361 16467 21419 16473
rect 22094 16464 22100 16476
rect 22152 16504 22158 16516
rect 22278 16504 22284 16516
rect 22152 16476 22284 16504
rect 22152 16464 22158 16476
rect 22278 16464 22284 16476
rect 22336 16464 22342 16516
rect 2774 16396 2780 16448
rect 2832 16436 2838 16448
rect 3789 16439 3847 16445
rect 3789 16436 3801 16439
rect 2832 16408 3801 16436
rect 2832 16396 2838 16408
rect 3789 16405 3801 16408
rect 3835 16405 3847 16439
rect 7098 16436 7104 16448
rect 7059 16408 7104 16436
rect 3789 16399 3847 16405
rect 7098 16396 7104 16408
rect 7156 16396 7162 16448
rect 11330 16436 11336 16448
rect 11291 16408 11336 16436
rect 11330 16396 11336 16408
rect 11388 16396 11394 16448
rect 12342 16436 12348 16448
rect 12303 16408 12348 16436
rect 12342 16396 12348 16408
rect 12400 16396 12406 16448
rect 16301 16439 16359 16445
rect 16301 16405 16313 16439
rect 16347 16436 16359 16439
rect 17770 16436 17776 16448
rect 16347 16408 17776 16436
rect 16347 16405 16359 16408
rect 16301 16399 16359 16405
rect 17770 16396 17776 16408
rect 17828 16396 17834 16448
rect 21450 16396 21456 16448
rect 21508 16436 21514 16448
rect 21818 16436 21824 16448
rect 21508 16408 21824 16436
rect 21508 16396 21514 16408
rect 21818 16396 21824 16408
rect 21876 16396 21882 16448
rect 22388 16436 22416 16544
rect 22649 16541 22661 16575
rect 22695 16572 22707 16575
rect 23566 16572 23572 16584
rect 22695 16544 23572 16572
rect 22695 16541 22707 16544
rect 22649 16535 22707 16541
rect 23566 16532 23572 16544
rect 23624 16532 23630 16584
rect 32122 16532 32128 16584
rect 32180 16572 32186 16584
rect 32493 16575 32551 16581
rect 32493 16572 32505 16575
rect 32180 16544 32505 16572
rect 32180 16532 32186 16544
rect 32493 16541 32505 16544
rect 32539 16541 32551 16575
rect 32493 16535 32551 16541
rect 33410 16532 33416 16584
rect 33468 16572 33474 16584
rect 33965 16575 34023 16581
rect 33965 16572 33977 16575
rect 33468 16544 33977 16572
rect 33468 16532 33474 16544
rect 33965 16541 33977 16544
rect 34011 16541 34023 16575
rect 33965 16535 34023 16541
rect 34606 16532 34612 16584
rect 34664 16572 34670 16584
rect 34900 16581 34928 16612
rect 34701 16575 34759 16581
rect 34701 16572 34713 16575
rect 34664 16544 34713 16572
rect 34664 16532 34670 16544
rect 34701 16541 34713 16544
rect 34747 16541 34759 16575
rect 34701 16535 34759 16541
rect 34885 16575 34943 16581
rect 34885 16541 34897 16575
rect 34931 16574 34943 16575
rect 34931 16546 34965 16574
rect 35710 16572 35716 16584
rect 34931 16541 34943 16546
rect 35671 16544 35716 16572
rect 34885 16535 34943 16541
rect 35710 16532 35716 16544
rect 35768 16532 35774 16584
rect 35989 16575 36047 16581
rect 35989 16572 36001 16575
rect 35866 16544 36001 16572
rect 23017 16507 23075 16513
rect 23017 16473 23029 16507
rect 23063 16504 23075 16507
rect 23658 16504 23664 16516
rect 23063 16476 23664 16504
rect 23063 16473 23075 16476
rect 23017 16467 23075 16473
rect 23658 16464 23664 16476
rect 23716 16464 23722 16516
rect 22741 16439 22799 16445
rect 22741 16436 22753 16439
rect 22388 16408 22753 16436
rect 22741 16405 22753 16408
rect 22787 16405 22799 16439
rect 22741 16399 22799 16405
rect 32677 16439 32735 16445
rect 32677 16405 32689 16439
rect 32723 16436 32735 16439
rect 33226 16436 33232 16448
rect 32723 16408 33232 16436
rect 32723 16405 32735 16408
rect 32677 16399 32735 16405
rect 33226 16396 33232 16408
rect 33284 16396 33290 16448
rect 34149 16439 34207 16445
rect 34149 16405 34161 16439
rect 34195 16436 34207 16439
rect 35866 16436 35894 16544
rect 35989 16541 36001 16544
rect 36035 16541 36047 16575
rect 35989 16535 36047 16541
rect 34195 16408 35894 16436
rect 34195 16405 34207 16408
rect 34149 16399 34207 16405
rect 1104 16346 38824 16368
rect 1104 16294 10398 16346
rect 10450 16294 10462 16346
rect 10514 16294 10526 16346
rect 10578 16294 10590 16346
rect 10642 16294 10654 16346
rect 10706 16294 19846 16346
rect 19898 16294 19910 16346
rect 19962 16294 19974 16346
rect 20026 16294 20038 16346
rect 20090 16294 20102 16346
rect 20154 16294 29294 16346
rect 29346 16294 29358 16346
rect 29410 16294 29422 16346
rect 29474 16294 29486 16346
rect 29538 16294 29550 16346
rect 29602 16294 38824 16346
rect 1104 16272 38824 16294
rect 2958 16232 2964 16244
rect 2919 16204 2964 16232
rect 2958 16192 2964 16204
rect 3016 16192 3022 16244
rect 10505 16235 10563 16241
rect 10505 16201 10517 16235
rect 10551 16232 10563 16235
rect 10778 16232 10784 16244
rect 10551 16204 10784 16232
rect 10551 16201 10563 16204
rect 10505 16195 10563 16201
rect 10778 16192 10784 16204
rect 10836 16192 10842 16244
rect 11517 16235 11575 16241
rect 11517 16201 11529 16235
rect 11563 16232 11575 16235
rect 11698 16232 11704 16244
rect 11563 16204 11704 16232
rect 11563 16201 11575 16204
rect 11517 16195 11575 16201
rect 11698 16192 11704 16204
rect 11756 16192 11762 16244
rect 19797 16235 19855 16241
rect 19797 16201 19809 16235
rect 19843 16232 19855 16235
rect 20622 16232 20628 16244
rect 19843 16204 20628 16232
rect 19843 16201 19855 16204
rect 19797 16195 19855 16201
rect 20622 16192 20628 16204
rect 20680 16192 20686 16244
rect 25866 16232 25872 16244
rect 25827 16204 25872 16232
rect 25866 16192 25872 16204
rect 25924 16192 25930 16244
rect 35897 16235 35955 16241
rect 35897 16201 35909 16235
rect 35943 16232 35955 16235
rect 36446 16232 36452 16244
rect 35943 16204 36452 16232
rect 35943 16201 35955 16204
rect 35897 16195 35955 16201
rect 36446 16192 36452 16204
rect 36504 16232 36510 16244
rect 36630 16232 36636 16244
rect 36504 16204 36636 16232
rect 36504 16192 36510 16204
rect 36630 16192 36636 16204
rect 36688 16192 36694 16244
rect 7837 16167 7895 16173
rect 7837 16133 7849 16167
rect 7883 16164 7895 16167
rect 8294 16164 8300 16176
rect 7883 16136 8300 16164
rect 7883 16133 7895 16136
rect 7837 16127 7895 16133
rect 8294 16124 8300 16136
rect 8352 16124 8358 16176
rect 11054 16124 11060 16176
rect 11112 16164 11118 16176
rect 12253 16167 12311 16173
rect 12253 16164 12265 16167
rect 11112 16136 12265 16164
rect 11112 16124 11118 16136
rect 12253 16133 12265 16136
rect 12299 16164 12311 16167
rect 14826 16164 14832 16176
rect 12299 16136 14832 16164
rect 12299 16133 12311 16136
rect 12253 16127 12311 16133
rect 14826 16124 14832 16136
rect 14884 16124 14890 16176
rect 26234 16124 26240 16176
rect 26292 16164 26298 16176
rect 26292 16136 26464 16164
rect 26292 16124 26298 16136
rect 2774 16096 2780 16108
rect 2735 16068 2780 16096
rect 2774 16056 2780 16068
rect 2832 16056 2838 16108
rect 9398 16056 9404 16108
rect 9456 16096 9462 16108
rect 10229 16099 10287 16105
rect 10229 16096 10241 16099
rect 9456 16068 10241 16096
rect 9456 16056 9462 16068
rect 10229 16065 10241 16068
rect 10275 16065 10287 16099
rect 10229 16059 10287 16065
rect 12342 16056 12348 16108
rect 12400 16096 12406 16108
rect 19613 16099 19671 16105
rect 19613 16096 19625 16099
rect 12400 16068 19625 16096
rect 12400 16056 12406 16068
rect 19613 16065 19625 16068
rect 19659 16065 19671 16099
rect 19613 16059 19671 16065
rect 25130 16056 25136 16108
rect 25188 16096 25194 16108
rect 26053 16099 26111 16105
rect 26053 16096 26065 16099
rect 25188 16068 26065 16096
rect 25188 16056 25194 16068
rect 26053 16065 26065 16068
rect 26099 16065 26111 16099
rect 26053 16059 26111 16065
rect 26145 16099 26203 16105
rect 26145 16065 26157 16099
rect 26191 16065 26203 16099
rect 26326 16096 26332 16108
rect 26287 16068 26332 16096
rect 26145 16059 26203 16065
rect 10134 16028 10140 16040
rect 10095 16000 10140 16028
rect 10134 15988 10140 16000
rect 10192 15988 10198 16040
rect 10318 15988 10324 16040
rect 10376 16028 10382 16040
rect 11698 16028 11704 16040
rect 10376 16000 11704 16028
rect 10376 15988 10382 16000
rect 11698 15988 11704 16000
rect 11756 15988 11762 16040
rect 11793 16031 11851 16037
rect 11793 15997 11805 16031
rect 11839 15997 11851 16031
rect 11793 15991 11851 15997
rect 8846 15920 8852 15972
rect 8904 15960 8910 15972
rect 11330 15960 11336 15972
rect 8904 15932 11336 15960
rect 8904 15920 8910 15932
rect 11330 15920 11336 15932
rect 11388 15960 11394 15972
rect 11808 15960 11836 15991
rect 24486 15988 24492 16040
rect 24544 16028 24550 16040
rect 26160 16028 26188 16059
rect 26326 16056 26332 16068
rect 26384 16056 26390 16108
rect 26436 16105 26464 16136
rect 26421 16099 26479 16105
rect 26421 16065 26433 16099
rect 26467 16065 26479 16099
rect 29733 16099 29791 16105
rect 29733 16096 29745 16099
rect 26421 16059 26479 16065
rect 27172 16068 29745 16096
rect 24544 16000 26188 16028
rect 26344 16028 26372 16056
rect 27172 16028 27200 16068
rect 29733 16065 29745 16068
rect 29779 16065 29791 16099
rect 29733 16059 29791 16065
rect 34514 16056 34520 16108
rect 34572 16096 34578 16108
rect 35710 16096 35716 16108
rect 34572 16068 35716 16096
rect 34572 16056 34578 16068
rect 35710 16056 35716 16068
rect 35768 16056 35774 16108
rect 26344 16000 27200 16028
rect 29549 16031 29607 16037
rect 24544 15988 24550 16000
rect 29549 15997 29561 16031
rect 29595 15997 29607 16031
rect 29549 15991 29607 15997
rect 12250 15960 12256 15972
rect 11388 15932 11836 15960
rect 12163 15932 12256 15960
rect 11388 15920 11394 15932
rect 12250 15920 12256 15932
rect 12308 15960 12314 15972
rect 16114 15960 16120 15972
rect 12308 15932 16120 15960
rect 12308 15920 12314 15932
rect 16114 15920 16120 15932
rect 16172 15920 16178 15972
rect 24302 15920 24308 15972
rect 24360 15960 24366 15972
rect 28997 15963 29055 15969
rect 28997 15960 29009 15963
rect 24360 15932 29009 15960
rect 24360 15920 24366 15932
rect 28997 15929 29009 15932
rect 29043 15960 29055 15963
rect 29564 15960 29592 15991
rect 34517 15963 34575 15969
rect 34517 15960 34529 15963
rect 29043 15932 34529 15960
rect 29043 15929 29055 15932
rect 28997 15923 29055 15929
rect 34517 15929 34529 15932
rect 34563 15960 34575 15963
rect 34606 15960 34612 15972
rect 34563 15932 34612 15960
rect 34563 15929 34575 15932
rect 34517 15923 34575 15929
rect 34606 15920 34612 15932
rect 34664 15920 34670 15972
rect 9030 15852 9036 15904
rect 9088 15892 9094 15904
rect 9125 15895 9183 15901
rect 9125 15892 9137 15895
rect 9088 15864 9137 15892
rect 9088 15852 9094 15864
rect 9125 15861 9137 15864
rect 9171 15892 9183 15895
rect 9490 15892 9496 15904
rect 9171 15864 9496 15892
rect 9171 15861 9183 15864
rect 9125 15855 9183 15861
rect 9490 15852 9496 15864
rect 9548 15852 9554 15904
rect 29917 15895 29975 15901
rect 29917 15861 29929 15895
rect 29963 15892 29975 15895
rect 30190 15892 30196 15904
rect 29963 15864 30196 15892
rect 29963 15861 29975 15864
rect 29917 15855 29975 15861
rect 30190 15852 30196 15864
rect 30248 15852 30254 15904
rect 1104 15802 38824 15824
rect 1104 15750 5674 15802
rect 5726 15750 5738 15802
rect 5790 15750 5802 15802
rect 5854 15750 5866 15802
rect 5918 15750 5930 15802
rect 5982 15750 15122 15802
rect 15174 15750 15186 15802
rect 15238 15750 15250 15802
rect 15302 15750 15314 15802
rect 15366 15750 15378 15802
rect 15430 15750 24570 15802
rect 24622 15750 24634 15802
rect 24686 15750 24698 15802
rect 24750 15750 24762 15802
rect 24814 15750 24826 15802
rect 24878 15750 34018 15802
rect 34070 15750 34082 15802
rect 34134 15750 34146 15802
rect 34198 15750 34210 15802
rect 34262 15750 34274 15802
rect 34326 15750 38824 15802
rect 1104 15728 38824 15750
rect 9674 15648 9680 15700
rect 9732 15688 9738 15700
rect 9861 15691 9919 15697
rect 9861 15688 9873 15691
rect 9732 15660 9873 15688
rect 9732 15648 9738 15660
rect 9861 15657 9873 15660
rect 9907 15657 9919 15691
rect 9861 15651 9919 15657
rect 24489 15691 24547 15697
rect 24489 15657 24501 15691
rect 24535 15688 24547 15691
rect 24946 15688 24952 15700
rect 24535 15660 24952 15688
rect 24535 15657 24547 15660
rect 24489 15651 24547 15657
rect 24946 15648 24952 15660
rect 25004 15648 25010 15700
rect 30742 15688 30748 15700
rect 30703 15660 30748 15688
rect 30742 15648 30748 15660
rect 30800 15648 30806 15700
rect 37458 15688 37464 15700
rect 37419 15660 37464 15688
rect 37458 15648 37464 15660
rect 37516 15648 37522 15700
rect 8386 15580 8392 15632
rect 8444 15620 8450 15632
rect 9125 15623 9183 15629
rect 9125 15620 9137 15623
rect 8444 15592 9137 15620
rect 8444 15580 8450 15592
rect 9125 15589 9137 15592
rect 9171 15620 9183 15623
rect 9398 15620 9404 15632
rect 9171 15592 9404 15620
rect 9171 15589 9183 15592
rect 9125 15583 9183 15589
rect 9398 15580 9404 15592
rect 9456 15620 9462 15632
rect 11425 15623 11483 15629
rect 11425 15620 11437 15623
rect 9456 15592 11437 15620
rect 9456 15580 9462 15592
rect 11425 15589 11437 15592
rect 11471 15589 11483 15623
rect 11425 15583 11483 15589
rect 11698 15580 11704 15632
rect 11756 15620 11762 15632
rect 14093 15623 14151 15629
rect 14093 15620 14105 15623
rect 11756 15592 14105 15620
rect 11756 15580 11762 15592
rect 14093 15589 14105 15592
rect 14139 15620 14151 15623
rect 15838 15620 15844 15632
rect 14139 15592 15844 15620
rect 14139 15589 14151 15592
rect 14093 15583 14151 15589
rect 15838 15580 15844 15592
rect 15896 15580 15902 15632
rect 27062 15620 27068 15632
rect 22066 15592 27068 15620
rect 2225 15555 2283 15561
rect 2225 15521 2237 15555
rect 2271 15552 2283 15555
rect 22066 15552 22094 15592
rect 27062 15580 27068 15592
rect 27120 15580 27126 15632
rect 2271 15524 22094 15552
rect 2271 15521 2283 15524
rect 2225 15515 2283 15521
rect 1673 15487 1731 15493
rect 1673 15453 1685 15487
rect 1719 15484 1731 15487
rect 2240 15484 2268 15515
rect 26234 15512 26240 15564
rect 26292 15552 26298 15564
rect 29733 15555 29791 15561
rect 29733 15552 29745 15555
rect 26292 15524 29745 15552
rect 26292 15512 26298 15524
rect 29733 15521 29745 15524
rect 29779 15521 29791 15555
rect 36446 15552 36452 15564
rect 36407 15524 36452 15552
rect 29733 15515 29791 15521
rect 36446 15512 36452 15524
rect 36504 15512 36510 15564
rect 1719 15456 2268 15484
rect 11609 15487 11667 15493
rect 1719 15453 1731 15456
rect 1673 15447 1731 15453
rect 11609 15453 11621 15487
rect 11655 15484 11667 15487
rect 12250 15484 12256 15496
rect 11655 15456 12256 15484
rect 11655 15453 11667 15456
rect 11609 15447 11667 15453
rect 12250 15444 12256 15456
rect 12308 15444 12314 15496
rect 14366 15484 14372 15496
rect 14327 15456 14372 15484
rect 14366 15444 14372 15456
rect 14424 15444 14430 15496
rect 14550 15484 14556 15496
rect 14511 15456 14556 15484
rect 14550 15444 14556 15456
rect 14608 15444 14614 15496
rect 14826 15484 14832 15496
rect 14787 15456 14832 15484
rect 14826 15444 14832 15456
rect 14884 15444 14890 15496
rect 15105 15487 15163 15493
rect 15105 15453 15117 15487
rect 15151 15484 15163 15487
rect 15746 15484 15752 15496
rect 15151 15456 15752 15484
rect 15151 15453 15163 15456
rect 15105 15447 15163 15453
rect 15746 15444 15752 15456
rect 15804 15444 15810 15496
rect 30006 15484 30012 15496
rect 29967 15456 30012 15484
rect 30006 15444 30012 15456
rect 30064 15444 30070 15496
rect 36722 15484 36728 15496
rect 36683 15456 36728 15484
rect 36722 15444 36728 15456
rect 36780 15444 36786 15496
rect 8846 15376 8852 15428
rect 8904 15416 8910 15428
rect 9125 15419 9183 15425
rect 9125 15416 9137 15419
rect 8904 15388 9137 15416
rect 8904 15376 8910 15388
rect 9125 15385 9137 15388
rect 9171 15385 9183 15419
rect 9125 15379 9183 15385
rect 9585 15419 9643 15425
rect 9585 15385 9597 15419
rect 9631 15416 9643 15419
rect 11054 15416 11060 15428
rect 9631 15388 11060 15416
rect 9631 15385 9643 15388
rect 9585 15379 9643 15385
rect 11054 15376 11060 15388
rect 11112 15376 11118 15428
rect 24486 15376 24492 15428
rect 24544 15416 24550 15428
rect 24673 15419 24731 15425
rect 24673 15416 24685 15419
rect 24544 15388 24685 15416
rect 24544 15376 24550 15388
rect 24673 15385 24685 15388
rect 24719 15385 24731 15419
rect 24673 15379 24731 15385
rect 24857 15419 24915 15425
rect 24857 15385 24869 15419
rect 24903 15416 24915 15419
rect 26050 15416 26056 15428
rect 24903 15388 26056 15416
rect 24903 15385 24915 15388
rect 24857 15379 24915 15385
rect 26050 15376 26056 15388
rect 26108 15376 26114 15428
rect 1486 15348 1492 15360
rect 1447 15320 1492 15348
rect 1486 15308 1492 15320
rect 1544 15308 1550 15360
rect 9674 15348 9680 15360
rect 9635 15320 9680 15348
rect 9674 15308 9680 15320
rect 9732 15308 9738 15360
rect 1104 15258 38824 15280
rect 1104 15206 10398 15258
rect 10450 15206 10462 15258
rect 10514 15206 10526 15258
rect 10578 15206 10590 15258
rect 10642 15206 10654 15258
rect 10706 15206 19846 15258
rect 19898 15206 19910 15258
rect 19962 15206 19974 15258
rect 20026 15206 20038 15258
rect 20090 15206 20102 15258
rect 20154 15206 29294 15258
rect 29346 15206 29358 15258
rect 29410 15206 29422 15258
rect 29474 15206 29486 15258
rect 29538 15206 29550 15258
rect 29602 15206 38824 15258
rect 1104 15184 38824 15206
rect 18782 15144 18788 15156
rect 18743 15116 18788 15144
rect 18782 15104 18788 15116
rect 18840 15104 18846 15156
rect 26237 15147 26295 15153
rect 26237 15113 26249 15147
rect 26283 15144 26295 15147
rect 27706 15144 27712 15156
rect 26283 15116 27712 15144
rect 26283 15113 26295 15116
rect 26237 15107 26295 15113
rect 27706 15104 27712 15116
rect 27764 15104 27770 15156
rect 30006 15144 30012 15156
rect 29967 15116 30012 15144
rect 30006 15104 30012 15116
rect 30064 15104 30070 15156
rect 35529 15147 35587 15153
rect 35529 15113 35541 15147
rect 35575 15144 35587 15147
rect 37458 15144 37464 15156
rect 35575 15116 37464 15144
rect 35575 15113 35587 15116
rect 35529 15107 35587 15113
rect 37458 15104 37464 15116
rect 37516 15104 37522 15156
rect 13814 15036 13820 15088
rect 13872 15076 13878 15088
rect 14550 15076 14556 15088
rect 13872 15048 14556 15076
rect 13872 15036 13878 15048
rect 14550 15036 14556 15048
rect 14608 15076 14614 15088
rect 25869 15079 25927 15085
rect 14608 15048 19012 15076
rect 14608 15036 14614 15048
rect 10413 15011 10471 15017
rect 10413 14977 10425 15011
rect 10459 15008 10471 15011
rect 11054 15008 11060 15020
rect 10459 14980 11060 15008
rect 10459 14977 10471 14980
rect 10413 14971 10471 14977
rect 11054 14968 11060 14980
rect 11112 14968 11118 15020
rect 14826 14968 14832 15020
rect 14884 15008 14890 15020
rect 16025 15011 16083 15017
rect 14884 14980 15884 15008
rect 14884 14968 14890 14980
rect 10134 14940 10140 14952
rect 10095 14912 10140 14940
rect 10134 14900 10140 14912
rect 10192 14900 10198 14952
rect 15746 14940 15752 14952
rect 15707 14912 15752 14940
rect 15746 14900 15752 14912
rect 15804 14900 15810 14952
rect 15856 14940 15884 14980
rect 16025 14977 16037 15011
rect 16071 15008 16083 15011
rect 16114 15008 16120 15020
rect 16071 14980 16120 15008
rect 16071 14977 16083 14980
rect 16025 14971 16083 14977
rect 16114 14968 16120 14980
rect 16172 14968 16178 15020
rect 17678 14968 17684 15020
rect 17736 15008 17742 15020
rect 18984 15017 19012 15048
rect 25869 15045 25881 15079
rect 25915 15076 25927 15079
rect 26418 15076 26424 15088
rect 25915 15048 26424 15076
rect 25915 15045 25927 15048
rect 25869 15039 25927 15045
rect 26418 15036 26424 15048
rect 26476 15036 26482 15088
rect 17773 15011 17831 15017
rect 17773 15008 17785 15011
rect 17736 14980 17785 15008
rect 17736 14968 17742 14980
rect 17773 14977 17785 14980
rect 17819 14977 17831 15011
rect 17773 14971 17831 14977
rect 18969 15011 19027 15017
rect 18969 14977 18981 15011
rect 19015 15008 19027 15011
rect 22002 15008 22008 15020
rect 19015 14980 22008 15008
rect 19015 14977 19027 14980
rect 18969 14971 19027 14977
rect 22002 14968 22008 14980
rect 22060 14968 22066 15020
rect 23474 14968 23480 15020
rect 23532 15008 23538 15020
rect 25777 15011 25835 15017
rect 25777 15008 25789 15011
rect 23532 14980 25789 15008
rect 23532 14968 23538 14980
rect 25777 14977 25789 14980
rect 25823 14977 25835 15011
rect 26050 15008 26056 15020
rect 26011 14980 26056 15008
rect 25777 14971 25835 14977
rect 17494 14940 17500 14952
rect 15856 14912 17500 14940
rect 17494 14900 17500 14912
rect 17552 14900 17558 14952
rect 25792 14940 25820 14971
rect 26050 14968 26056 14980
rect 26108 14968 26114 15020
rect 30190 15008 30196 15020
rect 30151 14980 30196 15008
rect 30190 14968 30196 14980
rect 30248 14968 30254 15020
rect 31478 14968 31484 15020
rect 31536 15008 31542 15020
rect 32861 15011 32919 15017
rect 32861 15008 32873 15011
rect 31536 14980 32873 15008
rect 31536 14968 31542 14980
rect 32861 14977 32873 14980
rect 32907 14977 32919 15011
rect 32861 14971 32919 14977
rect 33686 14968 33692 15020
rect 33744 15008 33750 15020
rect 34793 15011 34851 15017
rect 34793 15008 34805 15011
rect 33744 14980 34805 15008
rect 33744 14968 33750 14980
rect 34793 14977 34805 14980
rect 34839 14977 34851 15011
rect 34793 14971 34851 14977
rect 26970 14940 26976 14952
rect 25792 14912 26976 14940
rect 26970 14900 26976 14912
rect 27028 14900 27034 14952
rect 27249 14943 27307 14949
rect 27249 14909 27261 14943
rect 27295 14909 27307 14943
rect 34514 14940 34520 14952
rect 34427 14912 34520 14940
rect 27249 14903 27307 14909
rect 24486 14832 24492 14884
rect 24544 14872 24550 14884
rect 27264 14872 27292 14903
rect 34514 14900 34520 14912
rect 34572 14900 34578 14952
rect 24544 14844 27292 14872
rect 33045 14875 33103 14881
rect 24544 14832 24550 14844
rect 33045 14841 33057 14875
rect 33091 14872 33103 14875
rect 34532 14872 34560 14900
rect 33091 14844 34560 14872
rect 33091 14841 33103 14844
rect 33045 14835 33103 14841
rect 8846 14804 8852 14816
rect 8807 14776 8852 14804
rect 8846 14764 8852 14776
rect 8904 14764 8910 14816
rect 1104 14714 38824 14736
rect 1104 14662 5674 14714
rect 5726 14662 5738 14714
rect 5790 14662 5802 14714
rect 5854 14662 5866 14714
rect 5918 14662 5930 14714
rect 5982 14662 15122 14714
rect 15174 14662 15186 14714
rect 15238 14662 15250 14714
rect 15302 14662 15314 14714
rect 15366 14662 15378 14714
rect 15430 14662 24570 14714
rect 24622 14662 24634 14714
rect 24686 14662 24698 14714
rect 24750 14662 24762 14714
rect 24814 14662 24826 14714
rect 24878 14662 34018 14714
rect 34070 14662 34082 14714
rect 34134 14662 34146 14714
rect 34198 14662 34210 14714
rect 34262 14662 34274 14714
rect 34326 14662 38824 14714
rect 1104 14640 38824 14662
rect 26973 14603 27031 14609
rect 26973 14569 26985 14603
rect 27019 14600 27031 14603
rect 27246 14600 27252 14612
rect 27019 14572 27252 14600
rect 27019 14569 27031 14572
rect 26973 14563 27031 14569
rect 27246 14560 27252 14572
rect 27304 14600 27310 14612
rect 31294 14600 31300 14612
rect 27304 14572 31300 14600
rect 27304 14560 27310 14572
rect 31294 14560 31300 14572
rect 31352 14560 31358 14612
rect 31478 14600 31484 14612
rect 31439 14572 31484 14600
rect 31478 14560 31484 14572
rect 31536 14560 31542 14612
rect 33686 14600 33692 14612
rect 33647 14572 33692 14600
rect 33686 14560 33692 14572
rect 33744 14560 33750 14612
rect 15746 14492 15752 14544
rect 15804 14532 15810 14544
rect 15804 14504 21956 14532
rect 15804 14492 15810 14504
rect 9030 14464 9036 14476
rect 5460 14436 9036 14464
rect 1670 14396 1676 14408
rect 1631 14368 1676 14396
rect 1670 14356 1676 14368
rect 1728 14396 1734 14408
rect 2133 14399 2191 14405
rect 2133 14396 2145 14399
rect 1728 14368 2145 14396
rect 1728 14356 1734 14368
rect 2133 14365 2145 14368
rect 2179 14365 2191 14399
rect 2133 14359 2191 14365
rect 3786 14356 3792 14408
rect 3844 14396 3850 14408
rect 5460 14405 5488 14436
rect 9030 14424 9036 14436
rect 9088 14424 9094 14476
rect 9953 14467 10011 14473
rect 9953 14433 9965 14467
rect 9999 14464 10011 14467
rect 10318 14464 10324 14476
rect 9999 14436 10324 14464
rect 9999 14433 10011 14436
rect 9953 14427 10011 14433
rect 10318 14424 10324 14436
rect 10376 14424 10382 14476
rect 15197 14467 15255 14473
rect 15197 14433 15209 14467
rect 15243 14464 15255 14467
rect 15764 14464 15792 14492
rect 15243 14436 15792 14464
rect 15243 14433 15255 14436
rect 15197 14427 15255 14433
rect 15838 14424 15844 14476
rect 15896 14464 15902 14476
rect 16485 14467 16543 14473
rect 16485 14464 16497 14467
rect 15896 14436 16497 14464
rect 15896 14424 15902 14436
rect 16485 14433 16497 14436
rect 16531 14433 16543 14467
rect 16485 14427 16543 14433
rect 17494 14424 17500 14476
rect 17552 14464 17558 14476
rect 17865 14467 17923 14473
rect 17865 14464 17877 14467
rect 17552 14436 17877 14464
rect 17552 14424 17558 14436
rect 17865 14433 17877 14436
rect 17911 14433 17923 14467
rect 21818 14464 21824 14476
rect 21779 14436 21824 14464
rect 17865 14427 17923 14433
rect 21818 14424 21824 14436
rect 21876 14424 21882 14476
rect 21928 14464 21956 14504
rect 22306 14467 22364 14473
rect 22306 14464 22318 14467
rect 21928 14436 22318 14464
rect 22306 14433 22318 14436
rect 22352 14464 22364 14467
rect 22462 14464 22468 14476
rect 22352 14436 22468 14464
rect 22352 14433 22364 14436
rect 22306 14427 22364 14433
rect 22462 14424 22468 14436
rect 22520 14424 22526 14476
rect 23658 14424 23664 14476
rect 23716 14464 23722 14476
rect 30650 14464 30656 14476
rect 23716 14436 30656 14464
rect 23716 14424 23722 14436
rect 30650 14424 30656 14436
rect 30708 14464 30714 14476
rect 31205 14467 31263 14473
rect 31205 14464 31217 14467
rect 30708 14436 31217 14464
rect 30708 14424 30714 14436
rect 31205 14433 31217 14436
rect 31251 14433 31263 14467
rect 31205 14427 31263 14433
rect 5445 14399 5503 14405
rect 5445 14396 5457 14399
rect 3844 14368 5457 14396
rect 3844 14356 3850 14368
rect 5445 14365 5457 14368
rect 5491 14365 5503 14399
rect 9674 14396 9680 14408
rect 5445 14359 5503 14365
rect 8496 14368 9680 14396
rect 5721 14331 5779 14337
rect 5721 14297 5733 14331
rect 5767 14328 5779 14331
rect 5994 14328 6000 14340
rect 5767 14300 6000 14328
rect 5767 14297 5779 14300
rect 5721 14291 5779 14297
rect 5994 14288 6000 14300
rect 6052 14288 6058 14340
rect 7742 14328 7748 14340
rect 6946 14300 7748 14328
rect 7742 14288 7748 14300
rect 7800 14288 7806 14340
rect 1486 14260 1492 14272
rect 1447 14232 1492 14260
rect 1486 14220 1492 14232
rect 1544 14220 1550 14272
rect 7190 14260 7196 14272
rect 7151 14232 7196 14260
rect 7190 14220 7196 14232
rect 7248 14260 7254 14272
rect 8496 14260 8524 14368
rect 9674 14356 9680 14368
rect 9732 14356 9738 14408
rect 15470 14396 15476 14408
rect 15431 14368 15476 14396
rect 15470 14356 15476 14368
rect 15528 14356 15534 14408
rect 16761 14399 16819 14405
rect 16761 14365 16773 14399
rect 16807 14396 16819 14399
rect 17586 14396 17592 14408
rect 16807 14368 17592 14396
rect 16807 14365 16819 14368
rect 16761 14359 16819 14365
rect 17586 14356 17592 14368
rect 17644 14356 17650 14408
rect 18141 14399 18199 14405
rect 18141 14365 18153 14399
rect 18187 14396 18199 14399
rect 19334 14396 19340 14408
rect 18187 14368 19340 14396
rect 18187 14365 18199 14368
rect 18141 14359 18199 14365
rect 19334 14356 19340 14368
rect 19392 14356 19398 14408
rect 22097 14399 22155 14405
rect 22097 14365 22109 14399
rect 22143 14396 22155 14399
rect 22186 14396 22192 14408
rect 22143 14368 22192 14396
rect 22143 14365 22155 14368
rect 22097 14359 22155 14365
rect 22186 14356 22192 14368
rect 22244 14356 22250 14408
rect 26789 14399 26847 14405
rect 26789 14365 26801 14399
rect 26835 14396 26847 14399
rect 26970 14396 26976 14408
rect 26835 14368 26976 14396
rect 26835 14365 26847 14368
rect 26789 14359 26847 14365
rect 26970 14356 26976 14368
rect 27028 14356 27034 14408
rect 31113 14399 31171 14405
rect 31113 14365 31125 14399
rect 31159 14365 31171 14399
rect 31113 14359 31171 14365
rect 31941 14399 31999 14405
rect 31941 14365 31953 14399
rect 31987 14365 31999 14399
rect 31941 14359 31999 14365
rect 26050 14288 26056 14340
rect 26108 14328 26114 14340
rect 31128 14328 31156 14359
rect 31956 14328 31984 14359
rect 32490 14356 32496 14408
rect 32548 14396 32554 14408
rect 33505 14399 33563 14405
rect 33505 14396 33517 14399
rect 32548 14368 33517 14396
rect 32548 14356 32554 14368
rect 33505 14365 33517 14368
rect 33551 14365 33563 14399
rect 33505 14359 33563 14365
rect 26108 14300 31984 14328
rect 26108 14288 26114 14300
rect 7248 14232 8524 14260
rect 7248 14220 7254 14232
rect 20714 14220 20720 14272
rect 20772 14260 20778 14272
rect 21910 14260 21916 14272
rect 20772 14232 21916 14260
rect 20772 14220 20778 14232
rect 21910 14220 21916 14232
rect 21968 14260 21974 14272
rect 22189 14263 22247 14269
rect 22189 14260 22201 14263
rect 21968 14232 22201 14260
rect 21968 14220 21974 14232
rect 22189 14229 22201 14232
rect 22235 14229 22247 14263
rect 22189 14223 22247 14229
rect 22465 14263 22523 14269
rect 22465 14229 22477 14263
rect 22511 14260 22523 14263
rect 22830 14260 22836 14272
rect 22511 14232 22836 14260
rect 22511 14229 22523 14232
rect 22465 14223 22523 14229
rect 22830 14220 22836 14232
rect 22888 14260 22894 14272
rect 32030 14260 32036 14272
rect 22888 14232 32036 14260
rect 22888 14220 22894 14232
rect 32030 14220 32036 14232
rect 32088 14220 32094 14272
rect 32125 14263 32183 14269
rect 32125 14229 32137 14263
rect 32171 14260 32183 14263
rect 35342 14260 35348 14272
rect 32171 14232 35348 14260
rect 32171 14229 32183 14232
rect 32125 14223 32183 14229
rect 35342 14220 35348 14232
rect 35400 14220 35406 14272
rect 1104 14170 38824 14192
rect 1104 14118 10398 14170
rect 10450 14118 10462 14170
rect 10514 14118 10526 14170
rect 10578 14118 10590 14170
rect 10642 14118 10654 14170
rect 10706 14118 19846 14170
rect 19898 14118 19910 14170
rect 19962 14118 19974 14170
rect 20026 14118 20038 14170
rect 20090 14118 20102 14170
rect 20154 14118 29294 14170
rect 29346 14118 29358 14170
rect 29410 14118 29422 14170
rect 29474 14118 29486 14170
rect 29538 14118 29550 14170
rect 29602 14118 38824 14170
rect 1104 14096 38824 14118
rect 7742 14056 7748 14068
rect 7703 14028 7748 14056
rect 7742 14016 7748 14028
rect 7800 14016 7806 14068
rect 8389 14059 8447 14065
rect 8389 14025 8401 14059
rect 8435 14056 8447 14059
rect 9582 14056 9588 14068
rect 8435 14028 9588 14056
rect 8435 14025 8447 14028
rect 8389 14019 8447 14025
rect 7837 13923 7895 13929
rect 7837 13889 7849 13923
rect 7883 13920 7895 13923
rect 8404 13920 8432 14019
rect 9582 14016 9588 14028
rect 9640 14016 9646 14068
rect 22002 14016 22008 14068
rect 22060 14056 22066 14068
rect 22060 14016 22094 14056
rect 22186 14016 22192 14068
rect 22244 14056 22250 14068
rect 22465 14059 22523 14065
rect 22244 14028 22289 14056
rect 22244 14016 22250 14028
rect 22465 14025 22477 14059
rect 22511 14056 22523 14059
rect 23477 14059 23535 14065
rect 22511 14028 23428 14056
rect 22511 14025 22523 14028
rect 22465 14019 22523 14025
rect 15470 13948 15476 14000
rect 15528 13988 15534 14000
rect 18230 13988 18236 14000
rect 15528 13960 18236 13988
rect 15528 13948 15534 13960
rect 18230 13948 18236 13960
rect 18288 13988 18294 14000
rect 20898 13988 20904 14000
rect 18288 13960 20904 13988
rect 18288 13948 18294 13960
rect 20898 13948 20904 13960
rect 20956 13988 20962 14000
rect 21082 13988 21088 14000
rect 20956 13960 21088 13988
rect 20956 13948 20962 13960
rect 21082 13948 21088 13960
rect 21140 13988 21146 14000
rect 21818 13988 21824 14000
rect 21140 13960 21824 13988
rect 21140 13948 21146 13960
rect 21818 13948 21824 13960
rect 21876 13948 21882 14000
rect 22066 13988 22094 14016
rect 22306 13991 22364 13997
rect 22306 13988 22318 13991
rect 22066 13960 22318 13988
rect 22306 13957 22318 13960
rect 22352 13957 22364 13991
rect 22306 13951 22364 13957
rect 22554 13948 22560 14000
rect 22612 13988 22618 14000
rect 23293 13991 23351 13997
rect 23293 13988 23305 13991
rect 22612 13960 23305 13988
rect 22612 13948 22618 13960
rect 23293 13957 23305 13960
rect 23339 13957 23351 13991
rect 23400 13988 23428 14028
rect 23477 14025 23489 14059
rect 23523 14056 23535 14059
rect 23658 14056 23664 14068
rect 23523 14028 23664 14056
rect 23523 14025 23535 14028
rect 23477 14019 23535 14025
rect 23658 14016 23664 14028
rect 23716 14016 23722 14068
rect 32490 14056 32496 14068
rect 32451 14028 32496 14056
rect 32490 14016 32496 14028
rect 32548 14016 32554 14068
rect 23566 13988 23572 14000
rect 23400 13960 23572 13988
rect 23293 13951 23351 13957
rect 23566 13948 23572 13960
rect 23624 13948 23630 14000
rect 26234 13948 26240 14000
rect 26292 13988 26298 14000
rect 26973 13991 27031 13997
rect 26973 13988 26985 13991
rect 26292 13960 26985 13988
rect 26292 13948 26298 13960
rect 26973 13957 26985 13960
rect 27019 13957 27031 13991
rect 26973 13951 27031 13957
rect 17586 13920 17592 13932
rect 7883 13892 8432 13920
rect 17547 13892 17592 13920
rect 7883 13889 7895 13892
rect 7837 13883 7895 13889
rect 17586 13880 17592 13892
rect 17644 13920 17650 13932
rect 20714 13920 20720 13932
rect 17644 13892 20720 13920
rect 17644 13880 17650 13892
rect 20714 13880 20720 13892
rect 20772 13880 20778 13932
rect 22097 13923 22155 13929
rect 22097 13889 22109 13923
rect 22143 13889 22155 13923
rect 23584 13920 23612 13948
rect 27157 13923 27215 13929
rect 27157 13920 27169 13923
rect 23584 13892 27169 13920
rect 22097 13883 22155 13889
rect 27157 13889 27169 13892
rect 27203 13889 27215 13923
rect 27157 13883 27215 13889
rect 27249 13923 27307 13929
rect 27249 13889 27261 13923
rect 27295 13889 27307 13923
rect 27249 13883 27307 13889
rect 17865 13855 17923 13861
rect 17865 13821 17877 13855
rect 17911 13821 17923 13855
rect 17865 13815 17923 13821
rect 17880 13784 17908 13815
rect 21818 13812 21824 13864
rect 21876 13852 21882 13864
rect 21876 13824 21921 13852
rect 21876 13812 21882 13824
rect 18046 13784 18052 13796
rect 17880 13756 18052 13784
rect 18046 13744 18052 13756
rect 18104 13784 18110 13796
rect 21174 13784 21180 13796
rect 18104 13756 21180 13784
rect 18104 13744 18110 13756
rect 21174 13744 21180 13756
rect 21232 13744 21238 13796
rect 21910 13676 21916 13728
rect 21968 13716 21974 13728
rect 22112 13716 22140 13883
rect 22278 13812 22284 13864
rect 22336 13852 22342 13864
rect 22925 13855 22983 13861
rect 22925 13852 22937 13855
rect 22336 13824 22937 13852
rect 22336 13812 22342 13824
rect 22925 13821 22937 13824
rect 22971 13821 22983 13855
rect 26326 13852 26332 13864
rect 26287 13824 26332 13852
rect 22925 13815 22983 13821
rect 26326 13812 26332 13824
rect 26384 13812 26390 13864
rect 26344 13784 26372 13812
rect 27264 13784 27292 13883
rect 32030 13880 32036 13932
rect 32088 13920 32094 13932
rect 32309 13923 32367 13929
rect 32309 13920 32321 13923
rect 32088 13892 32321 13920
rect 32088 13880 32094 13892
rect 32309 13889 32321 13892
rect 32355 13889 32367 13923
rect 32309 13883 32367 13889
rect 30282 13812 30288 13864
rect 30340 13852 30346 13864
rect 31481 13855 31539 13861
rect 31481 13852 31493 13855
rect 30340 13824 31493 13852
rect 30340 13812 30346 13824
rect 31481 13821 31493 13824
rect 31527 13852 31539 13855
rect 32125 13855 32183 13861
rect 32125 13852 32137 13855
rect 31527 13824 32137 13852
rect 31527 13821 31539 13824
rect 31481 13815 31539 13821
rect 32125 13821 32137 13824
rect 32171 13821 32183 13855
rect 32125 13815 32183 13821
rect 26344 13756 27292 13784
rect 23293 13719 23351 13725
rect 23293 13716 23305 13719
rect 21968 13688 23305 13716
rect 21968 13676 21974 13688
rect 23293 13685 23305 13688
rect 23339 13685 23351 13719
rect 27246 13716 27252 13728
rect 27207 13688 27252 13716
rect 23293 13679 23351 13685
rect 27246 13676 27252 13688
rect 27304 13676 27310 13728
rect 27430 13716 27436 13728
rect 27391 13688 27436 13716
rect 27430 13676 27436 13688
rect 27488 13676 27494 13728
rect 1104 13626 38824 13648
rect 1104 13574 5674 13626
rect 5726 13574 5738 13626
rect 5790 13574 5802 13626
rect 5854 13574 5866 13626
rect 5918 13574 5930 13626
rect 5982 13574 15122 13626
rect 15174 13574 15186 13626
rect 15238 13574 15250 13626
rect 15302 13574 15314 13626
rect 15366 13574 15378 13626
rect 15430 13574 24570 13626
rect 24622 13574 24634 13626
rect 24686 13574 24698 13626
rect 24750 13574 24762 13626
rect 24814 13574 24826 13626
rect 24878 13574 34018 13626
rect 34070 13574 34082 13626
rect 34134 13574 34146 13626
rect 34198 13574 34210 13626
rect 34262 13574 34274 13626
rect 34326 13574 38824 13626
rect 1104 13552 38824 13574
rect 5994 13472 6000 13524
rect 6052 13512 6058 13524
rect 6365 13515 6423 13521
rect 6365 13512 6377 13515
rect 6052 13484 6377 13512
rect 6052 13472 6058 13484
rect 6365 13481 6377 13484
rect 6411 13481 6423 13515
rect 6365 13475 6423 13481
rect 8846 13472 8852 13524
rect 8904 13512 8910 13524
rect 11517 13515 11575 13521
rect 11517 13512 11529 13515
rect 8904 13484 11529 13512
rect 8904 13472 8910 13484
rect 11517 13481 11529 13484
rect 11563 13481 11575 13515
rect 11517 13475 11575 13481
rect 21085 13515 21143 13521
rect 21085 13481 21097 13515
rect 21131 13512 21143 13515
rect 21174 13512 21180 13524
rect 21131 13484 21180 13512
rect 21131 13481 21143 13484
rect 21085 13475 21143 13481
rect 1854 13404 1860 13456
rect 1912 13444 1918 13456
rect 7193 13447 7251 13453
rect 7193 13444 7205 13447
rect 1912 13416 7205 13444
rect 1912 13404 1918 13416
rect 7193 13413 7205 13416
rect 7239 13413 7251 13447
rect 7193 13407 7251 13413
rect 6549 13311 6607 13317
rect 6549 13277 6561 13311
rect 6595 13308 6607 13311
rect 7282 13308 7288 13320
rect 6595 13280 7288 13308
rect 6595 13277 6607 13280
rect 6549 13271 6607 13277
rect 7282 13268 7288 13280
rect 7340 13268 7346 13320
rect 7374 13268 7380 13320
rect 7432 13308 7438 13320
rect 8021 13311 8079 13317
rect 8021 13308 8033 13311
rect 7432 13280 8033 13308
rect 7432 13268 7438 13280
rect 8021 13277 8033 13280
rect 8067 13308 8079 13311
rect 9306 13308 9312 13320
rect 8067 13280 9312 13308
rect 8067 13277 8079 13280
rect 8021 13271 8079 13277
rect 9306 13268 9312 13280
rect 9364 13268 9370 13320
rect 11532 13308 11560 13475
rect 21174 13472 21180 13484
rect 21232 13472 21238 13524
rect 21266 13472 21272 13524
rect 21324 13512 21330 13524
rect 26326 13512 26332 13524
rect 21324 13484 26332 13512
rect 21324 13472 21330 13484
rect 26326 13472 26332 13484
rect 26384 13472 26390 13524
rect 12345 13447 12403 13453
rect 12345 13413 12357 13447
rect 12391 13444 12403 13447
rect 13814 13444 13820 13456
rect 12391 13416 13820 13444
rect 12391 13413 12403 13416
rect 12345 13407 12403 13413
rect 13814 13404 13820 13416
rect 13872 13404 13878 13456
rect 24302 13444 24308 13456
rect 13924 13416 24308 13444
rect 12161 13311 12219 13317
rect 12161 13308 12173 13311
rect 11532 13280 12173 13308
rect 12161 13277 12173 13280
rect 12207 13277 12219 13311
rect 12161 13271 12219 13277
rect 6886 13212 7880 13240
rect 2038 13132 2044 13184
rect 2096 13172 2102 13184
rect 6886 13172 6914 13212
rect 7852 13181 7880 13212
rect 2096 13144 6914 13172
rect 7837 13175 7895 13181
rect 2096 13132 2102 13144
rect 7837 13141 7849 13175
rect 7883 13141 7895 13175
rect 7837 13135 7895 13141
rect 8938 13132 8944 13184
rect 8996 13172 9002 13184
rect 9125 13175 9183 13181
rect 9125 13172 9137 13175
rect 8996 13144 9137 13172
rect 8996 13132 9002 13144
rect 9125 13141 9137 13144
rect 9171 13172 9183 13175
rect 13924 13172 13952 13416
rect 24302 13404 24308 13416
rect 24360 13404 24366 13456
rect 25041 13447 25099 13453
rect 25041 13413 25053 13447
rect 25087 13444 25099 13447
rect 26050 13444 26056 13456
rect 25087 13416 26056 13444
rect 25087 13413 25099 13416
rect 25041 13407 25099 13413
rect 26050 13404 26056 13416
rect 26108 13404 26114 13456
rect 16482 13336 16488 13388
rect 16540 13376 16546 13388
rect 17773 13379 17831 13385
rect 17773 13376 17785 13379
rect 16540 13348 17785 13376
rect 16540 13336 16546 13348
rect 14550 13268 14556 13320
rect 14608 13308 14614 13320
rect 17052 13317 17080 13348
rect 17773 13345 17785 13348
rect 17819 13345 17831 13379
rect 17773 13339 17831 13345
rect 19245 13379 19303 13385
rect 19245 13345 19257 13379
rect 19291 13376 19303 13379
rect 19610 13376 19616 13388
rect 19291 13348 19616 13376
rect 19291 13345 19303 13348
rect 19245 13339 19303 13345
rect 19610 13336 19616 13348
rect 19668 13336 19674 13388
rect 16853 13311 16911 13317
rect 16853 13308 16865 13311
rect 14608 13280 16865 13308
rect 14608 13268 14614 13280
rect 16853 13277 16865 13280
rect 16899 13277 16911 13311
rect 16853 13271 16911 13277
rect 17037 13311 17095 13317
rect 17037 13277 17049 13311
rect 17083 13277 17095 13311
rect 17037 13271 17095 13277
rect 17497 13311 17555 13317
rect 17497 13277 17509 13311
rect 17543 13308 17555 13311
rect 17678 13308 17684 13320
rect 17543 13280 17684 13308
rect 17543 13277 17555 13280
rect 17497 13271 17555 13277
rect 17678 13268 17684 13280
rect 17736 13268 17742 13320
rect 19518 13308 19524 13320
rect 19479 13280 19524 13308
rect 19518 13268 19524 13280
rect 19576 13268 19582 13320
rect 20824 13280 21496 13308
rect 16945 13243 17003 13249
rect 16945 13209 16957 13243
rect 16991 13240 17003 13243
rect 20824 13240 20852 13280
rect 16991 13212 20852 13240
rect 16991 13209 17003 13212
rect 16945 13203 17003 13209
rect 20898 13200 20904 13252
rect 20956 13240 20962 13252
rect 21468 13240 21496 13280
rect 21910 13268 21916 13320
rect 21968 13308 21974 13320
rect 22005 13311 22063 13317
rect 22005 13308 22017 13311
rect 21968 13280 22017 13308
rect 21968 13268 21974 13280
rect 22005 13277 22017 13280
rect 22051 13277 22063 13311
rect 22186 13308 22192 13320
rect 22147 13280 22192 13308
rect 22005 13271 22063 13277
rect 22186 13268 22192 13280
rect 22244 13268 22250 13320
rect 22462 13308 22468 13320
rect 22423 13280 22468 13308
rect 22462 13268 22468 13280
rect 22520 13268 22526 13320
rect 25130 13308 25136 13320
rect 24044 13280 25136 13308
rect 24044 13240 24072 13280
rect 25130 13268 25136 13280
rect 25188 13268 25194 13320
rect 20956 13212 21001 13240
rect 21468 13212 24072 13240
rect 24857 13243 24915 13249
rect 20956 13200 20962 13212
rect 24857 13209 24869 13243
rect 24903 13240 24915 13243
rect 25038 13240 25044 13252
rect 24903 13212 25044 13240
rect 24903 13209 24915 13212
rect 24857 13203 24915 13209
rect 25038 13200 25044 13212
rect 25096 13200 25102 13252
rect 9171 13144 13952 13172
rect 9171 13141 9183 13144
rect 9125 13135 9183 13141
rect 18782 13132 18788 13184
rect 18840 13172 18846 13184
rect 20990 13172 20996 13184
rect 18840 13144 20996 13172
rect 18840 13132 18846 13144
rect 20990 13132 20996 13144
rect 21048 13132 21054 13184
rect 21101 13175 21159 13181
rect 21101 13141 21113 13175
rect 21147 13172 21159 13175
rect 21910 13172 21916 13184
rect 21147 13144 21916 13172
rect 21147 13141 21159 13144
rect 21101 13135 21159 13141
rect 21910 13132 21916 13144
rect 21968 13132 21974 13184
rect 22649 13175 22707 13181
rect 22649 13141 22661 13175
rect 22695 13172 22707 13175
rect 23750 13172 23756 13184
rect 22695 13144 23756 13172
rect 22695 13141 22707 13144
rect 22649 13135 22707 13141
rect 23750 13132 23756 13144
rect 23808 13132 23814 13184
rect 1104 13082 38824 13104
rect 1104 13030 10398 13082
rect 10450 13030 10462 13082
rect 10514 13030 10526 13082
rect 10578 13030 10590 13082
rect 10642 13030 10654 13082
rect 10706 13030 19846 13082
rect 19898 13030 19910 13082
rect 19962 13030 19974 13082
rect 20026 13030 20038 13082
rect 20090 13030 20102 13082
rect 20154 13030 29294 13082
rect 29346 13030 29358 13082
rect 29410 13030 29422 13082
rect 29474 13030 29486 13082
rect 29538 13030 29550 13082
rect 29602 13030 38824 13082
rect 1104 13008 38824 13030
rect 3326 12928 3332 12980
rect 3384 12968 3390 12980
rect 3513 12971 3571 12977
rect 3513 12968 3525 12971
rect 3384 12940 3525 12968
rect 3384 12928 3390 12940
rect 3513 12937 3525 12940
rect 3559 12937 3571 12971
rect 3513 12931 3571 12937
rect 9306 12928 9312 12980
rect 9364 12968 9370 12980
rect 19518 12968 19524 12980
rect 9364 12940 19524 12968
rect 9364 12928 9370 12940
rect 19518 12928 19524 12940
rect 19576 12928 19582 12980
rect 21910 12968 21916 12980
rect 21823 12940 21916 12968
rect 21910 12928 21916 12940
rect 21968 12968 21974 12980
rect 26234 12968 26240 12980
rect 21968 12940 26240 12968
rect 21968 12928 21974 12940
rect 26234 12928 26240 12940
rect 26292 12928 26298 12980
rect 27154 12928 27160 12980
rect 27212 12977 27218 12980
rect 27212 12971 27231 12977
rect 27219 12937 27231 12971
rect 27212 12931 27231 12937
rect 27212 12928 27218 12931
rect 30558 12928 30564 12980
rect 30616 12968 30622 12980
rect 30653 12971 30711 12977
rect 30653 12968 30665 12971
rect 30616 12940 30665 12968
rect 30616 12928 30622 12940
rect 30653 12937 30665 12940
rect 30699 12968 30711 12971
rect 31110 12968 31116 12980
rect 30699 12940 31116 12968
rect 30699 12937 30711 12940
rect 30653 12931 30711 12937
rect 31110 12928 31116 12940
rect 31168 12968 31174 12980
rect 31573 12971 31631 12977
rect 31168 12940 31248 12968
rect 31168 12928 31174 12940
rect 2225 12903 2283 12909
rect 2225 12869 2237 12903
rect 2271 12900 2283 12903
rect 18782 12900 18788 12912
rect 2271 12872 18788 12900
rect 2271 12869 2283 12872
rect 2225 12863 2283 12869
rect 1673 12835 1731 12841
rect 1673 12801 1685 12835
rect 1719 12832 1731 12835
rect 2240 12832 2268 12863
rect 18782 12860 18788 12872
rect 18840 12860 18846 12912
rect 19058 12860 19064 12912
rect 19116 12900 19122 12912
rect 19245 12903 19303 12909
rect 19245 12900 19257 12903
rect 19116 12872 19257 12900
rect 19116 12860 19122 12872
rect 19245 12869 19257 12872
rect 19291 12869 19303 12903
rect 22186 12900 22192 12912
rect 19245 12863 19303 12869
rect 21836 12872 22192 12900
rect 1719 12804 2268 12832
rect 1719 12801 1731 12804
rect 1673 12795 1731 12801
rect 3142 12792 3148 12844
rect 3200 12832 3206 12844
rect 3421 12835 3479 12841
rect 3421 12832 3433 12835
rect 3200 12804 3433 12832
rect 3200 12792 3206 12804
rect 3421 12801 3433 12804
rect 3467 12801 3479 12835
rect 3421 12795 3479 12801
rect 3697 12835 3755 12841
rect 3697 12801 3709 12835
rect 3743 12832 3755 12835
rect 14185 12835 14243 12841
rect 3743 12804 4292 12832
rect 3743 12801 3755 12804
rect 3697 12795 3755 12801
rect 1486 12628 1492 12640
rect 1447 12600 1492 12628
rect 1486 12588 1492 12600
rect 1544 12588 1550 12640
rect 2961 12631 3019 12637
rect 2961 12597 2973 12631
rect 3007 12628 3019 12631
rect 3142 12628 3148 12640
rect 3007 12600 3148 12628
rect 3007 12597 3019 12600
rect 2961 12591 3019 12597
rect 3142 12588 3148 12600
rect 3200 12588 3206 12640
rect 3602 12588 3608 12640
rect 3660 12628 3666 12640
rect 4264 12637 4292 12804
rect 14185 12801 14197 12835
rect 14231 12832 14243 12835
rect 14458 12832 14464 12844
rect 14231 12804 14464 12832
rect 14231 12801 14243 12804
rect 14185 12795 14243 12801
rect 14458 12792 14464 12804
rect 14516 12792 14522 12844
rect 18601 12835 18659 12841
rect 18601 12832 18613 12835
rect 18340 12804 18613 12832
rect 13998 12764 14004 12776
rect 13959 12736 14004 12764
rect 13998 12724 14004 12736
rect 14056 12724 14062 12776
rect 14093 12767 14151 12773
rect 14093 12733 14105 12767
rect 14139 12733 14151 12767
rect 14093 12727 14151 12733
rect 14277 12767 14335 12773
rect 14277 12733 14289 12767
rect 14323 12764 14335 12767
rect 14366 12764 14372 12776
rect 14323 12736 14372 12764
rect 14323 12733 14335 12736
rect 14277 12727 14335 12733
rect 14108 12696 14136 12727
rect 14366 12724 14372 12736
rect 14424 12764 14430 12776
rect 18046 12764 18052 12776
rect 14424 12736 18052 12764
rect 14424 12724 14430 12736
rect 18046 12724 18052 12736
rect 18104 12724 18110 12776
rect 14642 12696 14648 12708
rect 14108 12668 14648 12696
rect 14642 12656 14648 12668
rect 14700 12656 14706 12708
rect 3697 12631 3755 12637
rect 3697 12628 3709 12631
rect 3660 12600 3709 12628
rect 3660 12588 3666 12600
rect 3697 12597 3709 12600
rect 3743 12597 3755 12631
rect 3697 12591 3755 12597
rect 4249 12631 4307 12637
rect 4249 12597 4261 12631
rect 4295 12628 4307 12631
rect 13262 12628 13268 12640
rect 4295 12600 13268 12628
rect 4295 12597 4307 12600
rect 4249 12591 4307 12597
rect 13262 12588 13268 12600
rect 13320 12628 13326 12640
rect 13630 12628 13636 12640
rect 13320 12600 13636 12628
rect 13320 12588 13326 12600
rect 13630 12588 13636 12600
rect 13688 12588 13694 12640
rect 13814 12628 13820 12640
rect 13775 12600 13820 12628
rect 13814 12588 13820 12600
rect 13872 12588 13878 12640
rect 14826 12628 14832 12640
rect 14787 12600 14832 12628
rect 14826 12588 14832 12600
rect 14884 12588 14890 12640
rect 17957 12631 18015 12637
rect 17957 12597 17969 12631
rect 18003 12628 18015 12631
rect 18340 12628 18368 12804
rect 18601 12801 18613 12804
rect 18647 12801 18659 12835
rect 19334 12832 19340 12844
rect 19295 12804 19340 12832
rect 18601 12795 18659 12801
rect 19334 12792 19340 12804
rect 19392 12832 19398 12844
rect 21836 12841 21864 12872
rect 22186 12860 22192 12872
rect 22244 12860 22250 12912
rect 31220 12909 31248 12940
rect 31573 12937 31585 12971
rect 31619 12968 31631 12971
rect 33505 12971 33563 12977
rect 31619 12940 33456 12968
rect 31619 12937 31631 12940
rect 31573 12931 31631 12937
rect 26973 12903 27031 12909
rect 26973 12900 26985 12903
rect 26344 12872 26985 12900
rect 21821 12835 21879 12841
rect 21821 12832 21833 12835
rect 19392 12804 21833 12832
rect 19392 12792 19398 12804
rect 21821 12801 21833 12804
rect 21867 12801 21879 12835
rect 22002 12832 22008 12844
rect 21963 12804 22008 12832
rect 21821 12795 21879 12801
rect 22002 12792 22008 12804
rect 22060 12792 22066 12844
rect 23750 12832 23756 12844
rect 23711 12804 23756 12832
rect 23750 12792 23756 12804
rect 23808 12792 23814 12844
rect 18417 12767 18475 12773
rect 18417 12733 18429 12767
rect 18463 12764 18475 12767
rect 19426 12764 19432 12776
rect 18463 12736 19432 12764
rect 18463 12733 18475 12736
rect 18417 12727 18475 12733
rect 19426 12724 19432 12736
rect 19484 12724 19490 12776
rect 23937 12699 23995 12705
rect 23937 12665 23949 12699
rect 23983 12696 23995 12699
rect 25038 12696 25044 12708
rect 23983 12668 25044 12696
rect 23983 12665 23995 12668
rect 23937 12659 23995 12665
rect 25038 12656 25044 12668
rect 25096 12656 25102 12708
rect 19610 12628 19616 12640
rect 18003 12600 19616 12628
rect 18003 12597 18015 12600
rect 17957 12591 18015 12597
rect 19610 12588 19616 12600
rect 19668 12628 19674 12640
rect 20165 12631 20223 12637
rect 20165 12628 20177 12631
rect 19668 12600 20177 12628
rect 19668 12588 19674 12600
rect 20165 12597 20177 12600
rect 20211 12597 20223 12631
rect 20165 12591 20223 12597
rect 22462 12588 22468 12640
rect 22520 12628 22526 12640
rect 26344 12637 26372 12872
rect 26973 12869 26985 12872
rect 27019 12869 27031 12903
rect 26973 12863 27031 12869
rect 31205 12903 31263 12909
rect 31205 12869 31217 12903
rect 31251 12869 31263 12903
rect 31205 12863 31263 12869
rect 26988 12832 27016 12863
rect 31294 12860 31300 12912
rect 31352 12900 31358 12912
rect 31410 12903 31468 12909
rect 31410 12900 31422 12903
rect 31352 12872 31422 12900
rect 31352 12860 31358 12872
rect 31410 12869 31422 12872
rect 31456 12900 31468 12903
rect 31456 12872 31524 12900
rect 31456 12869 31468 12872
rect 31410 12863 31468 12869
rect 30282 12832 30288 12844
rect 26988 12804 30288 12832
rect 30282 12792 30288 12804
rect 30340 12792 30346 12844
rect 31496 12832 31524 12872
rect 31662 12860 31668 12912
rect 31720 12900 31726 12912
rect 31938 12900 31944 12912
rect 31720 12872 31944 12900
rect 31720 12860 31726 12872
rect 31938 12860 31944 12872
rect 31996 12900 32002 12912
rect 32125 12903 32183 12909
rect 32125 12900 32137 12903
rect 31996 12872 32137 12900
rect 31996 12860 32002 12872
rect 32125 12869 32137 12872
rect 32171 12869 32183 12903
rect 32325 12903 32383 12909
rect 32325 12900 32337 12903
rect 32125 12863 32183 12869
rect 32232 12872 32337 12900
rect 32232 12832 32260 12872
rect 32325 12869 32337 12872
rect 32371 12869 32383 12903
rect 32325 12863 32383 12869
rect 33321 12835 33379 12841
rect 33321 12832 33333 12835
rect 31496 12804 32260 12832
rect 32508 12804 33333 12832
rect 32508 12705 32536 12804
rect 33321 12801 33333 12804
rect 33367 12801 33379 12835
rect 33428 12832 33456 12940
rect 33505 12937 33517 12971
rect 33551 12937 33563 12971
rect 33505 12931 33563 12937
rect 33520 12900 33548 12931
rect 33520 12872 35664 12900
rect 34609 12835 34667 12841
rect 34609 12832 34621 12835
rect 33428 12804 34621 12832
rect 33321 12795 33379 12801
rect 34609 12801 34621 12804
rect 34655 12801 34667 12835
rect 35342 12832 35348 12844
rect 35303 12804 35348 12832
rect 34609 12795 34667 12801
rect 35342 12792 35348 12804
rect 35400 12792 35406 12844
rect 35636 12841 35664 12872
rect 35621 12835 35679 12841
rect 35621 12801 35633 12835
rect 35667 12801 35679 12835
rect 35621 12795 35679 12801
rect 32493 12699 32551 12705
rect 31404 12668 31754 12696
rect 26329 12631 26387 12637
rect 26329 12628 26341 12631
rect 22520 12600 26341 12628
rect 22520 12588 22526 12600
rect 26329 12597 26341 12600
rect 26375 12597 26387 12631
rect 26329 12591 26387 12597
rect 26418 12588 26424 12640
rect 26476 12628 26482 12640
rect 27157 12631 27215 12637
rect 27157 12628 27169 12631
rect 26476 12600 27169 12628
rect 26476 12588 26482 12600
rect 27157 12597 27169 12600
rect 27203 12597 27215 12631
rect 27338 12628 27344 12640
rect 27299 12600 27344 12628
rect 27157 12591 27215 12597
rect 27338 12588 27344 12600
rect 27396 12588 27402 12640
rect 31404 12637 31432 12668
rect 31726 12640 31754 12668
rect 32493 12665 32505 12699
rect 32539 12665 32551 12699
rect 32493 12659 32551 12665
rect 31389 12631 31447 12637
rect 31389 12597 31401 12631
rect 31435 12597 31447 12631
rect 31726 12600 31760 12640
rect 31389 12591 31447 12597
rect 31754 12588 31760 12600
rect 31812 12628 31818 12640
rect 32309 12631 32367 12637
rect 32309 12628 32321 12631
rect 31812 12600 32321 12628
rect 31812 12588 31818 12600
rect 32309 12597 32321 12600
rect 32355 12597 32367 12631
rect 32309 12591 32367 12597
rect 34793 12631 34851 12637
rect 34793 12597 34805 12631
rect 34839 12628 34851 12631
rect 36078 12628 36084 12640
rect 34839 12600 36084 12628
rect 34839 12597 34851 12600
rect 34793 12591 34851 12597
rect 36078 12588 36084 12600
rect 36136 12588 36142 12640
rect 36354 12628 36360 12640
rect 36315 12600 36360 12628
rect 36354 12588 36360 12600
rect 36412 12588 36418 12640
rect 1104 12538 38824 12560
rect 1104 12486 5674 12538
rect 5726 12486 5738 12538
rect 5790 12486 5802 12538
rect 5854 12486 5866 12538
rect 5918 12486 5930 12538
rect 5982 12486 15122 12538
rect 15174 12486 15186 12538
rect 15238 12486 15250 12538
rect 15302 12486 15314 12538
rect 15366 12486 15378 12538
rect 15430 12486 24570 12538
rect 24622 12486 24634 12538
rect 24686 12486 24698 12538
rect 24750 12486 24762 12538
rect 24814 12486 24826 12538
rect 24878 12486 34018 12538
rect 34070 12486 34082 12538
rect 34134 12486 34146 12538
rect 34198 12486 34210 12538
rect 34262 12486 34274 12538
rect 34326 12486 38824 12538
rect 1104 12464 38824 12486
rect 5534 12424 5540 12436
rect 5493 12396 5540 12424
rect 5534 12384 5540 12396
rect 5592 12433 5598 12436
rect 5592 12427 5641 12433
rect 5592 12393 5595 12427
rect 5629 12424 5641 12427
rect 8846 12424 8852 12436
rect 5629 12396 8852 12424
rect 5629 12393 5641 12396
rect 5592 12387 5641 12393
rect 5592 12384 5598 12387
rect 8846 12384 8852 12396
rect 8904 12384 8910 12436
rect 31938 12424 31944 12436
rect 31899 12396 31944 12424
rect 31938 12384 31944 12396
rect 31996 12384 32002 12436
rect 13998 12356 14004 12368
rect 4908 12328 14004 12356
rect 3786 12288 3792 12300
rect 3747 12260 3792 12288
rect 3786 12248 3792 12260
rect 3844 12248 3850 12300
rect 4908 12288 4936 12328
rect 13998 12316 14004 12328
rect 14056 12356 14062 12368
rect 14826 12356 14832 12368
rect 14056 12328 14832 12356
rect 14056 12316 14062 12328
rect 3988 12260 4936 12288
rect 3053 12223 3111 12229
rect 3053 12220 3065 12223
rect 2746 12192 3065 12220
rect 2746 12152 2774 12192
rect 3053 12189 3065 12192
rect 3099 12220 3111 12223
rect 3988 12220 4016 12260
rect 7282 12248 7288 12300
rect 7340 12288 7346 12300
rect 12710 12288 12716 12300
rect 7340 12260 12716 12288
rect 7340 12248 7346 12260
rect 12710 12248 12716 12260
rect 12768 12248 12774 12300
rect 13541 12291 13599 12297
rect 13541 12257 13553 12291
rect 13587 12288 13599 12291
rect 13722 12288 13728 12300
rect 13587 12260 13728 12288
rect 13587 12257 13599 12260
rect 13541 12251 13599 12257
rect 13722 12248 13728 12260
rect 13780 12248 13786 12300
rect 14366 12288 14372 12300
rect 14327 12260 14372 12288
rect 14366 12248 14372 12260
rect 14424 12248 14430 12300
rect 14752 12297 14780 12328
rect 14826 12316 14832 12328
rect 14884 12356 14890 12368
rect 15197 12359 15255 12365
rect 15197 12356 15209 12359
rect 14884 12328 15209 12356
rect 14884 12316 14890 12328
rect 15197 12325 15209 12328
rect 15243 12325 15255 12359
rect 15197 12319 15255 12325
rect 14737 12291 14795 12297
rect 14737 12257 14749 12291
rect 14783 12257 14795 12291
rect 14737 12251 14795 12257
rect 34790 12248 34796 12300
rect 34848 12288 34854 12300
rect 35342 12288 35348 12300
rect 34848 12260 35348 12288
rect 34848 12248 34854 12260
rect 35342 12248 35348 12260
rect 35400 12288 35406 12300
rect 35805 12291 35863 12297
rect 35805 12288 35817 12291
rect 35400 12260 35817 12288
rect 35400 12248 35406 12260
rect 35805 12257 35817 12260
rect 35851 12257 35863 12291
rect 35805 12251 35863 12257
rect 4154 12220 4160 12232
rect 3099 12192 4016 12220
rect 4115 12192 4160 12220
rect 3099 12189 3111 12192
rect 3053 12183 3111 12189
rect 4154 12180 4160 12192
rect 4212 12180 4218 12232
rect 9401 12223 9459 12229
rect 5276 12192 6592 12220
rect 2424 12124 2774 12152
rect 2130 12044 2136 12096
rect 2188 12084 2194 12096
rect 2424 12093 2452 12124
rect 5166 12112 5172 12164
rect 5224 12112 5230 12164
rect 2409 12087 2467 12093
rect 2409 12084 2421 12087
rect 2188 12056 2421 12084
rect 2188 12044 2194 12056
rect 2409 12053 2421 12056
rect 2455 12053 2467 12087
rect 3142 12084 3148 12096
rect 3055 12056 3148 12084
rect 2409 12047 2467 12053
rect 3142 12044 3148 12056
rect 3200 12084 3206 12096
rect 3418 12084 3424 12096
rect 3200 12056 3424 12084
rect 3200 12044 3206 12056
rect 3418 12044 3424 12056
rect 3476 12084 3482 12096
rect 5276 12084 5304 12192
rect 6564 12152 6592 12192
rect 9401 12189 9413 12223
rect 9447 12220 9459 12223
rect 9582 12220 9588 12232
rect 9447 12192 9588 12220
rect 9447 12189 9459 12192
rect 9401 12183 9459 12189
rect 9582 12180 9588 12192
rect 9640 12220 9646 12232
rect 9861 12223 9919 12229
rect 9861 12220 9873 12223
rect 9640 12192 9873 12220
rect 9640 12180 9646 12192
rect 9861 12189 9873 12192
rect 9907 12189 9919 12223
rect 13262 12220 13268 12232
rect 13223 12192 13268 12220
rect 9861 12183 9919 12189
rect 13262 12180 13268 12192
rect 13320 12180 13326 12232
rect 13630 12180 13636 12232
rect 13688 12220 13694 12232
rect 14277 12223 14335 12229
rect 14277 12220 14289 12223
rect 13688 12192 14289 12220
rect 13688 12180 13694 12192
rect 14277 12189 14289 12192
rect 14323 12189 14335 12223
rect 14277 12183 14335 12189
rect 25041 12223 25099 12229
rect 25041 12189 25053 12223
rect 25087 12220 25099 12223
rect 26234 12220 26240 12232
rect 25087 12192 26240 12220
rect 25087 12189 25099 12192
rect 25041 12183 25099 12189
rect 26234 12180 26240 12192
rect 26292 12180 26298 12232
rect 27338 12220 27344 12232
rect 27299 12192 27344 12220
rect 27338 12180 27344 12192
rect 27396 12180 27402 12232
rect 36078 12220 36084 12232
rect 36039 12192 36084 12220
rect 36078 12180 36084 12192
rect 36136 12180 36142 12232
rect 14366 12152 14372 12164
rect 6564 12124 14372 12152
rect 14366 12112 14372 12124
rect 14424 12112 14430 12164
rect 16482 12152 16488 12164
rect 14568 12124 16488 12152
rect 9214 12084 9220 12096
rect 3476 12056 5304 12084
rect 9175 12056 9220 12084
rect 3476 12044 3482 12056
rect 9214 12044 9220 12056
rect 9272 12044 9278 12096
rect 13170 12044 13176 12096
rect 13228 12084 13234 12096
rect 14093 12087 14151 12093
rect 14093 12084 14105 12087
rect 13228 12056 14105 12084
rect 13228 12044 13234 12056
rect 14093 12053 14105 12056
rect 14139 12053 14151 12087
rect 14093 12047 14151 12053
rect 14458 12044 14464 12096
rect 14516 12084 14522 12096
rect 14568 12093 14596 12124
rect 16482 12112 16488 12124
rect 16540 12112 16546 12164
rect 31754 12152 31760 12164
rect 26206 12124 31760 12152
rect 14553 12087 14611 12093
rect 14553 12084 14565 12087
rect 14516 12056 14565 12084
rect 14516 12044 14522 12056
rect 14553 12053 14565 12056
rect 14599 12053 14611 12087
rect 14553 12047 14611 12053
rect 14642 12044 14648 12096
rect 14700 12084 14706 12096
rect 25222 12084 25228 12096
rect 14700 12056 14745 12084
rect 25183 12056 25228 12084
rect 14700 12044 14706 12056
rect 25222 12044 25228 12056
rect 25280 12084 25286 12096
rect 26206 12084 26234 12124
rect 31754 12112 31760 12124
rect 31812 12112 31818 12164
rect 25280 12056 26234 12084
rect 27157 12087 27215 12093
rect 25280 12044 25286 12056
rect 27157 12053 27169 12087
rect 27203 12084 27215 12087
rect 27246 12084 27252 12096
rect 27203 12056 27252 12084
rect 27203 12053 27215 12056
rect 27157 12047 27215 12053
rect 27246 12044 27252 12056
rect 27304 12044 27310 12096
rect 34514 12044 34520 12096
rect 34572 12084 34578 12096
rect 35802 12084 35808 12096
rect 34572 12056 35808 12084
rect 34572 12044 34578 12056
rect 35802 12044 35808 12056
rect 35860 12084 35866 12096
rect 36354 12084 36360 12096
rect 35860 12056 36360 12084
rect 35860 12044 35866 12056
rect 36354 12044 36360 12056
rect 36412 12084 36418 12096
rect 36817 12087 36875 12093
rect 36817 12084 36829 12087
rect 36412 12056 36829 12084
rect 36412 12044 36418 12056
rect 36817 12053 36829 12056
rect 36863 12053 36875 12087
rect 36817 12047 36875 12053
rect 1104 11994 38824 12016
rect 1104 11942 10398 11994
rect 10450 11942 10462 11994
rect 10514 11942 10526 11994
rect 10578 11942 10590 11994
rect 10642 11942 10654 11994
rect 10706 11942 19846 11994
rect 19898 11942 19910 11994
rect 19962 11942 19974 11994
rect 20026 11942 20038 11994
rect 20090 11942 20102 11994
rect 20154 11942 29294 11994
rect 29346 11942 29358 11994
rect 29410 11942 29422 11994
rect 29474 11942 29486 11994
rect 29538 11942 29550 11994
rect 29602 11942 38824 11994
rect 1104 11920 38824 11942
rect 3789 11883 3847 11889
rect 3789 11849 3801 11883
rect 3835 11880 3847 11883
rect 4154 11880 4160 11892
rect 3835 11852 4160 11880
rect 3835 11849 3847 11852
rect 3789 11843 3847 11849
rect 4154 11840 4160 11852
rect 4212 11840 4218 11892
rect 5166 11840 5172 11892
rect 5224 11880 5230 11892
rect 6457 11883 6515 11889
rect 6457 11880 6469 11883
rect 5224 11852 6469 11880
rect 5224 11840 5230 11852
rect 6457 11849 6469 11852
rect 6503 11849 6515 11883
rect 6457 11843 6515 11849
rect 8573 11883 8631 11889
rect 8573 11849 8585 11883
rect 8619 11880 8631 11883
rect 9122 11880 9128 11892
rect 8619 11852 9128 11880
rect 8619 11849 8631 11852
rect 8573 11843 8631 11849
rect 9122 11840 9128 11852
rect 9180 11880 9186 11892
rect 12710 11880 12716 11892
rect 9180 11852 10824 11880
rect 12671 11852 12716 11880
rect 9180 11840 9186 11852
rect 10042 11772 10048 11824
rect 10100 11772 10106 11824
rect 1673 11747 1731 11753
rect 1673 11713 1685 11747
rect 1719 11744 1731 11747
rect 2869 11747 2927 11753
rect 1719 11716 2268 11744
rect 1719 11713 1731 11716
rect 1673 11707 1731 11713
rect 2240 11552 2268 11716
rect 2869 11713 2881 11747
rect 2915 11744 2927 11747
rect 3418 11744 3424 11756
rect 2915 11716 3424 11744
rect 2915 11713 2927 11716
rect 2869 11707 2927 11713
rect 3418 11704 3424 11716
rect 3476 11704 3482 11756
rect 3602 11744 3608 11756
rect 3563 11716 3608 11744
rect 3602 11704 3608 11716
rect 3660 11704 3666 11756
rect 6549 11747 6607 11753
rect 6549 11713 6561 11747
rect 6595 11744 6607 11747
rect 9214 11744 9220 11756
rect 6595 11716 9220 11744
rect 6595 11713 6607 11716
rect 6549 11707 6607 11713
rect 9214 11704 9220 11716
rect 9272 11704 9278 11756
rect 10796 11753 10824 11852
rect 12710 11840 12716 11852
rect 12768 11840 12774 11892
rect 14458 11880 14464 11892
rect 14419 11852 14464 11880
rect 14458 11840 14464 11852
rect 14516 11840 14522 11892
rect 14550 11840 14556 11892
rect 14608 11880 14614 11892
rect 14608 11852 14653 11880
rect 14608 11840 14614 11852
rect 13170 11812 13176 11824
rect 13131 11784 13176 11812
rect 13170 11772 13176 11784
rect 13228 11772 13234 11824
rect 25038 11772 25044 11824
rect 25096 11812 25102 11824
rect 25096 11784 28488 11812
rect 25096 11772 25102 11784
rect 10781 11747 10839 11753
rect 10781 11713 10793 11747
rect 10827 11744 10839 11747
rect 11790 11744 11796 11756
rect 10827 11716 11796 11744
rect 10827 11713 10839 11716
rect 10781 11707 10839 11713
rect 11790 11704 11796 11716
rect 11848 11704 11854 11756
rect 13630 11704 13636 11756
rect 13688 11744 13694 11756
rect 14185 11747 14243 11753
rect 14185 11744 14197 11747
rect 13688 11716 14197 11744
rect 13688 11704 13694 11716
rect 14185 11713 14197 11716
rect 14231 11713 14243 11747
rect 14185 11707 14243 11713
rect 14366 11704 14372 11756
rect 14424 11744 14430 11756
rect 14645 11747 14703 11753
rect 14645 11744 14657 11747
rect 14424 11716 14657 11744
rect 14424 11704 14430 11716
rect 14645 11713 14657 11716
rect 14691 11744 14703 11747
rect 14734 11744 14740 11756
rect 14691 11716 14740 11744
rect 14691 11713 14703 11716
rect 14645 11707 14703 11713
rect 14734 11704 14740 11716
rect 14792 11744 14798 11756
rect 15105 11747 15163 11753
rect 15105 11744 15117 11747
rect 14792 11716 15117 11744
rect 14792 11704 14798 11716
rect 15105 11713 15117 11716
rect 15151 11713 15163 11747
rect 18046 11744 18052 11756
rect 18007 11716 18052 11744
rect 15105 11707 15163 11713
rect 18046 11704 18052 11716
rect 18104 11704 18110 11756
rect 18230 11744 18236 11756
rect 18191 11716 18236 11744
rect 18230 11704 18236 11716
rect 18288 11704 18294 11756
rect 26988 11753 27016 11784
rect 26973 11747 27031 11753
rect 26973 11713 26985 11747
rect 27019 11713 27031 11747
rect 27246 11744 27252 11756
rect 27207 11716 27252 11744
rect 26973 11707 27031 11713
rect 27246 11704 27252 11716
rect 27304 11704 27310 11756
rect 28460 11753 28488 11784
rect 28445 11747 28503 11753
rect 28445 11713 28457 11747
rect 28491 11713 28503 11747
rect 28718 11744 28724 11756
rect 28679 11716 28724 11744
rect 28445 11707 28503 11713
rect 28718 11704 28724 11716
rect 28776 11704 28782 11756
rect 3326 11676 3332 11688
rect 3287 11648 3332 11676
rect 3326 11636 3332 11648
rect 3384 11636 3390 11688
rect 9232 11676 9260 11704
rect 10134 11676 10140 11688
rect 9232 11648 10140 11676
rect 10134 11636 10140 11648
rect 10192 11636 10198 11688
rect 10505 11679 10563 11685
rect 10505 11645 10517 11679
rect 10551 11676 10563 11679
rect 10551 11648 14228 11676
rect 10551 11645 10563 11648
rect 10505 11639 10563 11645
rect 12897 11611 12955 11617
rect 12897 11577 12909 11611
rect 12943 11608 12955 11611
rect 13814 11608 13820 11620
rect 12943 11580 13820 11608
rect 12943 11577 12955 11580
rect 12897 11571 12955 11577
rect 13814 11568 13820 11580
rect 13872 11568 13878 11620
rect 14200 11617 14228 11648
rect 14185 11611 14243 11617
rect 14185 11577 14197 11611
rect 14231 11577 14243 11611
rect 14185 11571 14243 11577
rect 16666 11568 16672 11620
rect 16724 11608 16730 11620
rect 16724 11580 26234 11608
rect 16724 11568 16730 11580
rect 1486 11540 1492 11552
rect 1447 11512 1492 11540
rect 1486 11500 1492 11512
rect 1544 11500 1550 11552
rect 2222 11540 2228 11552
rect 2183 11512 2228 11540
rect 2222 11500 2228 11512
rect 2280 11500 2286 11552
rect 6270 11500 6276 11552
rect 6328 11540 6334 11552
rect 9033 11543 9091 11549
rect 9033 11540 9045 11543
rect 6328 11512 9045 11540
rect 6328 11500 6334 11512
rect 9033 11509 9045 11512
rect 9079 11540 9091 11543
rect 9950 11540 9956 11552
rect 9079 11512 9956 11540
rect 9079 11509 9091 11512
rect 9033 11503 9091 11509
rect 9950 11500 9956 11512
rect 10008 11500 10014 11552
rect 14274 11500 14280 11552
rect 14332 11540 14338 11552
rect 18046 11540 18052 11552
rect 14332 11512 14377 11540
rect 18007 11512 18052 11540
rect 14332 11500 14338 11512
rect 18046 11500 18052 11512
rect 18104 11500 18110 11552
rect 26206 11540 26234 11580
rect 27985 11543 28043 11549
rect 27985 11540 27997 11543
rect 26206 11512 27997 11540
rect 27985 11509 27997 11512
rect 28031 11540 28043 11543
rect 29457 11543 29515 11549
rect 29457 11540 29469 11543
rect 28031 11512 29469 11540
rect 28031 11509 28043 11512
rect 27985 11503 28043 11509
rect 29457 11509 29469 11512
rect 29503 11540 29515 11543
rect 34514 11540 34520 11552
rect 29503 11512 34520 11540
rect 29503 11509 29515 11512
rect 29457 11503 29515 11509
rect 34514 11500 34520 11512
rect 34572 11500 34578 11552
rect 1104 11450 38824 11472
rect 1104 11398 5674 11450
rect 5726 11398 5738 11450
rect 5790 11398 5802 11450
rect 5854 11398 5866 11450
rect 5918 11398 5930 11450
rect 5982 11398 15122 11450
rect 15174 11398 15186 11450
rect 15238 11398 15250 11450
rect 15302 11398 15314 11450
rect 15366 11398 15378 11450
rect 15430 11398 24570 11450
rect 24622 11398 24634 11450
rect 24686 11398 24698 11450
rect 24750 11398 24762 11450
rect 24814 11398 24826 11450
rect 24878 11398 34018 11450
rect 34070 11398 34082 11450
rect 34134 11398 34146 11450
rect 34198 11398 34210 11450
rect 34262 11398 34274 11450
rect 34326 11398 38824 11450
rect 1104 11376 38824 11398
rect 10042 11336 10048 11348
rect 10003 11308 10048 11336
rect 10042 11296 10048 11308
rect 10100 11296 10106 11348
rect 13541 11339 13599 11345
rect 13541 11305 13553 11339
rect 13587 11336 13599 11339
rect 13630 11336 13636 11348
rect 13587 11308 13636 11336
rect 13587 11305 13599 11308
rect 13541 11299 13599 11305
rect 13630 11296 13636 11308
rect 13688 11296 13694 11348
rect 14274 11296 14280 11348
rect 14332 11336 14338 11348
rect 16485 11339 16543 11345
rect 16485 11336 16497 11339
rect 14332 11308 16497 11336
rect 14332 11296 14338 11308
rect 16485 11305 16497 11308
rect 16531 11305 16543 11339
rect 16485 11299 16543 11305
rect 24581 11339 24639 11345
rect 24581 11305 24593 11339
rect 24627 11336 24639 11339
rect 25222 11336 25228 11348
rect 24627 11308 25228 11336
rect 24627 11305 24639 11308
rect 24581 11299 24639 11305
rect 25222 11296 25228 11308
rect 25280 11296 25286 11348
rect 26973 11339 27031 11345
rect 26973 11305 26985 11339
rect 27019 11336 27031 11339
rect 28718 11336 28724 11348
rect 27019 11308 28724 11336
rect 27019 11305 27031 11308
rect 26973 11299 27031 11305
rect 28718 11296 28724 11308
rect 28776 11296 28782 11348
rect 31665 11339 31723 11345
rect 31665 11305 31677 11339
rect 31711 11336 31723 11339
rect 31754 11336 31760 11348
rect 31711 11308 31760 11336
rect 31711 11305 31723 11308
rect 31665 11299 31723 11305
rect 31754 11296 31760 11308
rect 31812 11336 31818 11348
rect 32493 11339 32551 11345
rect 32493 11336 32505 11339
rect 31812 11308 32505 11336
rect 31812 11296 31818 11308
rect 32493 11305 32505 11308
rect 32539 11305 32551 11339
rect 32493 11299 32551 11305
rect 2222 11228 2228 11280
rect 2280 11268 2286 11280
rect 2280 11240 2774 11268
rect 2280 11228 2286 11240
rect 2746 11200 2774 11240
rect 14550 11228 14556 11280
rect 14608 11268 14614 11280
rect 14737 11271 14795 11277
rect 14737 11268 14749 11271
rect 14608 11240 14749 11268
rect 14608 11228 14614 11240
rect 14737 11237 14749 11240
rect 14783 11237 14795 11271
rect 14737 11231 14795 11237
rect 14826 11228 14832 11280
rect 14884 11268 14890 11280
rect 24765 11271 24823 11277
rect 14884 11240 16804 11268
rect 14884 11228 14890 11240
rect 16666 11200 16672 11212
rect 2746 11172 16672 11200
rect 16666 11160 16672 11172
rect 16724 11160 16730 11212
rect 10134 11132 10140 11144
rect 10095 11104 10140 11132
rect 10134 11092 10140 11104
rect 10192 11092 10198 11144
rect 13262 11092 13268 11144
rect 13320 11132 13326 11144
rect 14553 11135 14611 11141
rect 14553 11132 14565 11135
rect 13320 11104 14565 11132
rect 13320 11092 13326 11104
rect 14553 11101 14565 11104
rect 14599 11132 14611 11135
rect 14642 11132 14648 11144
rect 14599 11104 14648 11132
rect 14599 11101 14611 11104
rect 14553 11095 14611 11101
rect 14642 11092 14648 11104
rect 14700 11132 14706 11144
rect 16022 11132 16028 11144
rect 14700 11104 16028 11132
rect 14700 11092 14706 11104
rect 16022 11092 16028 11104
rect 16080 11092 16086 11144
rect 16482 11132 16488 11144
rect 16443 11104 16488 11132
rect 16482 11092 16488 11104
rect 16540 11092 16546 11144
rect 16776 11141 16804 11240
rect 24765 11237 24777 11271
rect 24811 11268 24823 11271
rect 32677 11271 32735 11277
rect 24811 11240 26234 11268
rect 24811 11237 24823 11240
rect 24765 11231 24823 11237
rect 16761 11135 16819 11141
rect 16761 11101 16773 11135
rect 16807 11132 16819 11135
rect 26206 11132 26234 11240
rect 32677 11237 32689 11271
rect 32723 11268 32735 11271
rect 33686 11268 33692 11280
rect 32723 11240 33692 11268
rect 32723 11237 32735 11240
rect 32677 11231 32735 11237
rect 33686 11228 33692 11240
rect 33744 11228 33750 11280
rect 31021 11203 31079 11209
rect 31021 11169 31033 11203
rect 31067 11200 31079 11203
rect 31478 11200 31484 11212
rect 31067 11172 31484 11200
rect 31067 11169 31079 11172
rect 31021 11163 31079 11169
rect 31478 11160 31484 11172
rect 31536 11200 31542 11212
rect 32214 11200 32220 11212
rect 31536 11172 32220 11200
rect 31536 11160 31542 11172
rect 32214 11160 32220 11172
rect 32272 11160 32278 11212
rect 26789 11135 26847 11141
rect 26789 11132 26801 11135
rect 16807 11104 17356 11132
rect 26206 11104 26801 11132
rect 16807 11101 16819 11104
rect 16761 11095 16819 11101
rect 17328 11073 17356 11104
rect 26789 11101 26801 11104
rect 26835 11101 26847 11135
rect 26789 11095 26847 11101
rect 31420 11104 32444 11132
rect 17313 11067 17371 11073
rect 17313 11033 17325 11067
rect 17359 11064 17371 11067
rect 23566 11064 23572 11076
rect 17359 11036 23572 11064
rect 17359 11033 17371 11036
rect 17313 11027 17371 11033
rect 23566 11024 23572 11036
rect 23624 11024 23630 11076
rect 23750 11024 23756 11076
rect 23808 11064 23814 11076
rect 24397 11067 24455 11073
rect 24397 11064 24409 11067
rect 23808 11036 24409 11064
rect 23808 11024 23814 11036
rect 24397 11033 24409 11036
rect 24443 11033 24455 11067
rect 24397 11027 24455 11033
rect 24486 11024 24492 11076
rect 24544 11064 24550 11076
rect 24613 11067 24671 11073
rect 24613 11064 24625 11067
rect 24544 11036 24625 11064
rect 24544 11024 24550 11036
rect 24613 11033 24625 11036
rect 24659 11064 24671 11067
rect 31420 11064 31448 11104
rect 24659 11036 31448 11064
rect 24659 11033 24671 11036
rect 24613 11027 24671 11033
rect 31478 11024 31484 11076
rect 31536 11064 31542 11076
rect 31680 11073 31708 11104
rect 31680 11067 31739 11073
rect 31536 11036 31581 11064
rect 31680 11036 31693 11067
rect 31536 11024 31542 11036
rect 31681 11033 31693 11036
rect 31727 11033 31739 11067
rect 31681 11027 31739 11033
rect 32030 11024 32036 11076
rect 32088 11064 32094 11076
rect 32309 11067 32367 11073
rect 32309 11064 32321 11067
rect 32088 11036 32321 11064
rect 32088 11024 32094 11036
rect 32309 11033 32321 11036
rect 32355 11033 32367 11067
rect 32416 11064 32444 11104
rect 32509 11067 32567 11073
rect 32509 11064 32521 11067
rect 32416 11036 32521 11064
rect 32309 11027 32367 11033
rect 32509 11033 32521 11036
rect 32555 11033 32567 11067
rect 32509 11027 32567 11033
rect 16666 10996 16672 11008
rect 16627 10968 16672 10996
rect 16666 10956 16672 10968
rect 16724 10956 16730 11008
rect 31846 10996 31852 11008
rect 31807 10968 31852 10996
rect 31846 10956 31852 10968
rect 31904 10956 31910 11008
rect 1104 10906 38824 10928
rect 1104 10854 10398 10906
rect 10450 10854 10462 10906
rect 10514 10854 10526 10906
rect 10578 10854 10590 10906
rect 10642 10854 10654 10906
rect 10706 10854 19846 10906
rect 19898 10854 19910 10906
rect 19962 10854 19974 10906
rect 20026 10854 20038 10906
rect 20090 10854 20102 10906
rect 20154 10854 29294 10906
rect 29346 10854 29358 10906
rect 29410 10854 29422 10906
rect 29474 10854 29486 10906
rect 29538 10854 29550 10906
rect 29602 10854 38824 10906
rect 1104 10832 38824 10854
rect 3326 10752 3332 10804
rect 3384 10792 3390 10804
rect 18046 10792 18052 10804
rect 3384 10764 7328 10792
rect 18007 10764 18052 10792
rect 3384 10752 3390 10764
rect 7098 10733 7104 10736
rect 7085 10727 7104 10733
rect 7085 10693 7097 10727
rect 7085 10687 7104 10693
rect 7098 10684 7104 10687
rect 7156 10684 7162 10736
rect 7300 10733 7328 10764
rect 18046 10752 18052 10764
rect 18104 10752 18110 10804
rect 22922 10792 22928 10804
rect 22296 10764 22928 10792
rect 7285 10727 7343 10733
rect 7285 10693 7297 10727
rect 7331 10724 7343 10727
rect 14550 10724 14556 10736
rect 7331 10696 14556 10724
rect 7331 10693 7343 10696
rect 7285 10687 7343 10693
rect 14550 10684 14556 10696
rect 14608 10684 14614 10736
rect 16666 10684 16672 10736
rect 16724 10724 16730 10736
rect 17862 10724 17868 10736
rect 16724 10696 17868 10724
rect 16724 10684 16730 10696
rect 17862 10684 17868 10696
rect 17920 10724 17926 10736
rect 18233 10727 18291 10733
rect 18233 10724 18245 10727
rect 17920 10696 18245 10724
rect 17920 10684 17926 10696
rect 18233 10693 18245 10696
rect 18279 10693 18291 10727
rect 18233 10687 18291 10693
rect 18417 10727 18475 10733
rect 18417 10693 18429 10727
rect 18463 10724 18475 10727
rect 19058 10724 19064 10736
rect 18463 10696 19064 10724
rect 18463 10693 18475 10696
rect 18417 10687 18475 10693
rect 19058 10684 19064 10696
rect 19116 10684 19122 10736
rect 22296 10733 22324 10764
rect 22922 10752 22928 10764
rect 22980 10752 22986 10804
rect 32030 10752 32036 10804
rect 32088 10792 32094 10804
rect 32125 10795 32183 10801
rect 32125 10792 32137 10795
rect 32088 10764 32137 10792
rect 32088 10752 32094 10764
rect 32125 10761 32137 10764
rect 32171 10761 32183 10795
rect 32125 10755 32183 10761
rect 33229 10795 33287 10801
rect 33229 10761 33241 10795
rect 33275 10761 33287 10795
rect 35802 10792 35808 10804
rect 35763 10764 35808 10792
rect 33229 10755 33287 10761
rect 22281 10727 22339 10733
rect 22281 10693 22293 10727
rect 22327 10693 22339 10727
rect 22462 10724 22468 10736
rect 22423 10696 22468 10724
rect 22281 10687 22339 10693
rect 22462 10684 22468 10696
rect 22520 10684 22526 10736
rect 33244 10724 33272 10755
rect 35802 10752 35808 10764
rect 35860 10752 35866 10804
rect 33244 10696 35112 10724
rect 18141 10659 18199 10665
rect 18141 10625 18153 10659
rect 18187 10656 18199 10659
rect 18966 10656 18972 10668
rect 18187 10628 18972 10656
rect 18187 10625 18199 10628
rect 18141 10619 18199 10625
rect 18966 10616 18972 10628
rect 19024 10616 19030 10668
rect 31846 10616 31852 10668
rect 31904 10656 31910 10668
rect 33045 10659 33103 10665
rect 33045 10656 33057 10659
rect 31904 10628 33057 10656
rect 31904 10616 31910 10628
rect 33045 10625 33057 10628
rect 33091 10625 33103 10659
rect 33686 10656 33692 10668
rect 33647 10628 33692 10656
rect 33045 10619 33103 10625
rect 33686 10616 33692 10628
rect 33744 10616 33750 10668
rect 34790 10656 34796 10668
rect 34751 10628 34796 10656
rect 34790 10616 34796 10628
rect 34848 10616 34854 10668
rect 35084 10665 35112 10696
rect 35069 10659 35127 10665
rect 35069 10625 35081 10659
rect 35115 10625 35127 10659
rect 35069 10619 35127 10625
rect 4890 10412 4896 10464
rect 4948 10452 4954 10464
rect 6917 10455 6975 10461
rect 6917 10452 6929 10455
rect 4948 10424 6929 10452
rect 4948 10412 4954 10424
rect 6917 10421 6929 10424
rect 6963 10421 6975 10455
rect 6917 10415 6975 10421
rect 7101 10455 7159 10461
rect 7101 10421 7113 10455
rect 7147 10452 7159 10455
rect 7374 10452 7380 10464
rect 7147 10424 7380 10452
rect 7147 10421 7159 10424
rect 7101 10415 7159 10421
rect 7374 10412 7380 10424
rect 7432 10412 7438 10464
rect 17586 10412 17592 10464
rect 17644 10452 17650 10464
rect 17865 10455 17923 10461
rect 17865 10452 17877 10455
rect 17644 10424 17877 10452
rect 17644 10412 17650 10424
rect 17865 10421 17877 10424
rect 17911 10421 17923 10455
rect 18966 10452 18972 10464
rect 18927 10424 18972 10452
rect 17865 10415 17923 10421
rect 18966 10412 18972 10424
rect 19024 10412 19030 10464
rect 33873 10455 33931 10461
rect 33873 10421 33885 10455
rect 33919 10452 33931 10455
rect 35710 10452 35716 10464
rect 33919 10424 35716 10452
rect 33919 10421 33931 10424
rect 33873 10415 33931 10421
rect 35710 10412 35716 10424
rect 35768 10412 35774 10464
rect 1104 10362 38824 10384
rect 1104 10310 5674 10362
rect 5726 10310 5738 10362
rect 5790 10310 5802 10362
rect 5854 10310 5866 10362
rect 5918 10310 5930 10362
rect 5982 10310 15122 10362
rect 15174 10310 15186 10362
rect 15238 10310 15250 10362
rect 15302 10310 15314 10362
rect 15366 10310 15378 10362
rect 15430 10310 24570 10362
rect 24622 10310 24634 10362
rect 24686 10310 24698 10362
rect 24750 10310 24762 10362
rect 24814 10310 24826 10362
rect 24878 10310 34018 10362
rect 34070 10310 34082 10362
rect 34134 10310 34146 10362
rect 34198 10310 34210 10362
rect 34262 10310 34274 10362
rect 34326 10310 38824 10362
rect 1104 10288 38824 10310
rect 35802 10208 35808 10260
rect 35860 10248 35866 10260
rect 36541 10251 36599 10257
rect 36541 10248 36553 10251
rect 35860 10220 36553 10248
rect 35860 10208 35866 10220
rect 36541 10217 36553 10220
rect 36587 10217 36599 10251
rect 36541 10211 36599 10217
rect 16022 10112 16028 10124
rect 15983 10084 16028 10112
rect 16022 10072 16028 10084
rect 16080 10072 16086 10124
rect 16301 10115 16359 10121
rect 16301 10081 16313 10115
rect 16347 10112 16359 10115
rect 16666 10112 16672 10124
rect 16347 10084 16672 10112
rect 16347 10081 16359 10084
rect 16301 10075 16359 10081
rect 16666 10072 16672 10084
rect 16724 10072 16730 10124
rect 34790 10072 34796 10124
rect 34848 10112 34854 10124
rect 35529 10115 35587 10121
rect 35529 10112 35541 10115
rect 34848 10084 35541 10112
rect 34848 10072 34854 10084
rect 35529 10081 35541 10084
rect 35575 10081 35587 10115
rect 35529 10075 35587 10081
rect 1673 10047 1731 10053
rect 1673 10013 1685 10047
rect 1719 10044 1731 10047
rect 4890 10044 4896 10056
rect 1719 10016 2268 10044
rect 4851 10016 4896 10044
rect 1719 10013 1731 10016
rect 1673 10007 1731 10013
rect 2240 9985 2268 10016
rect 4890 10004 4896 10016
rect 4948 10004 4954 10056
rect 27430 10044 27436 10056
rect 27391 10016 27436 10044
rect 27430 10004 27436 10016
rect 27488 10004 27494 10056
rect 35710 10004 35716 10056
rect 35768 10044 35774 10056
rect 35805 10047 35863 10053
rect 35805 10044 35817 10047
rect 35768 10016 35817 10044
rect 35768 10004 35774 10016
rect 35805 10013 35817 10016
rect 35851 10013 35863 10047
rect 35805 10007 35863 10013
rect 2225 9979 2283 9985
rect 2225 9945 2237 9979
rect 2271 9976 2283 9979
rect 20806 9976 20812 9988
rect 2271 9948 20812 9976
rect 2271 9945 2283 9948
rect 2225 9939 2283 9945
rect 20806 9936 20812 9948
rect 20864 9936 20870 9988
rect 1486 9908 1492 9920
rect 1447 9880 1492 9908
rect 1486 9868 1492 9880
rect 1544 9868 1550 9920
rect 4706 9908 4712 9920
rect 4667 9880 4712 9908
rect 4706 9868 4712 9880
rect 4764 9868 4770 9920
rect 27249 9911 27307 9917
rect 27249 9877 27261 9911
rect 27295 9908 27307 9911
rect 27430 9908 27436 9920
rect 27295 9880 27436 9908
rect 27295 9877 27307 9880
rect 27249 9871 27307 9877
rect 27430 9868 27436 9880
rect 27488 9868 27494 9920
rect 1104 9818 38824 9840
rect 1104 9766 10398 9818
rect 10450 9766 10462 9818
rect 10514 9766 10526 9818
rect 10578 9766 10590 9818
rect 10642 9766 10654 9818
rect 10706 9766 19846 9818
rect 19898 9766 19910 9818
rect 19962 9766 19974 9818
rect 20026 9766 20038 9818
rect 20090 9766 20102 9818
rect 20154 9766 29294 9818
rect 29346 9766 29358 9818
rect 29410 9766 29422 9818
rect 29474 9766 29486 9818
rect 29538 9766 29550 9818
rect 29602 9766 38824 9818
rect 1104 9744 38824 9766
rect 7193 9639 7251 9645
rect 7193 9605 7205 9639
rect 7239 9636 7251 9639
rect 13262 9636 13268 9648
rect 7239 9608 13268 9636
rect 7239 9605 7251 9608
rect 7193 9599 7251 9605
rect 13262 9596 13268 9608
rect 13320 9596 13326 9648
rect 18966 9596 18972 9648
rect 19024 9636 19030 9648
rect 22462 9636 22468 9648
rect 19024 9608 22468 9636
rect 19024 9596 19030 9608
rect 22462 9596 22468 9608
rect 22520 9596 22526 9648
rect 22002 9528 22008 9580
rect 22060 9568 22066 9580
rect 22097 9571 22155 9577
rect 22097 9568 22109 9571
rect 22060 9540 22109 9568
rect 22060 9528 22066 9540
rect 22097 9537 22109 9540
rect 22143 9537 22155 9571
rect 22922 9568 22928 9580
rect 22883 9540 22928 9568
rect 22097 9531 22155 9537
rect 22922 9528 22928 9540
rect 22980 9528 22986 9580
rect 24394 9568 24400 9580
rect 24355 9540 24400 9568
rect 24394 9528 24400 9540
rect 24452 9528 24458 9580
rect 20254 9460 20260 9512
rect 20312 9500 20318 9512
rect 21821 9503 21879 9509
rect 21821 9500 21833 9503
rect 20312 9472 21833 9500
rect 20312 9460 20318 9472
rect 21821 9469 21833 9472
rect 21867 9469 21879 9503
rect 21821 9463 21879 9469
rect 26786 9460 26792 9512
rect 26844 9500 26850 9512
rect 30650 9500 30656 9512
rect 26844 9472 30656 9500
rect 26844 9460 26850 9472
rect 30650 9460 30656 9472
rect 30708 9460 30714 9512
rect 1946 9392 1952 9444
rect 2004 9432 2010 9444
rect 3694 9432 3700 9444
rect 2004 9404 3700 9432
rect 2004 9392 2010 9404
rect 3694 9392 3700 9404
rect 3752 9392 3758 9444
rect 6914 9432 6920 9444
rect 6875 9404 6920 9432
rect 6914 9392 6920 9404
rect 6972 9392 6978 9444
rect 30374 9432 30380 9444
rect 22388 9404 30380 9432
rect 3237 9367 3295 9373
rect 3237 9333 3249 9367
rect 3283 9364 3295 9367
rect 4982 9364 4988 9376
rect 3283 9336 4988 9364
rect 3283 9333 3295 9336
rect 3237 9327 3295 9333
rect 4982 9324 4988 9336
rect 5040 9324 5046 9376
rect 6638 9324 6644 9376
rect 6696 9364 6702 9376
rect 6733 9367 6791 9373
rect 6733 9364 6745 9367
rect 6696 9336 6745 9364
rect 6696 9324 6702 9336
rect 6733 9333 6745 9336
rect 6779 9333 6791 9367
rect 6733 9327 6791 9333
rect 20622 9324 20628 9376
rect 20680 9364 20686 9376
rect 22388 9364 22416 9404
rect 30374 9392 30380 9404
rect 30432 9392 30438 9444
rect 20680 9336 22416 9364
rect 24581 9367 24639 9373
rect 20680 9324 20686 9336
rect 24581 9333 24593 9367
rect 24627 9364 24639 9367
rect 27154 9364 27160 9376
rect 24627 9336 27160 9364
rect 24627 9333 24639 9336
rect 24581 9327 24639 9333
rect 27154 9324 27160 9336
rect 27212 9324 27218 9376
rect 30466 9324 30472 9376
rect 30524 9364 30530 9376
rect 31021 9367 31079 9373
rect 31021 9364 31033 9367
rect 30524 9336 31033 9364
rect 30524 9324 30530 9336
rect 31021 9333 31033 9336
rect 31067 9333 31079 9367
rect 31021 9327 31079 9333
rect 1104 9274 38824 9296
rect 1104 9222 5674 9274
rect 5726 9222 5738 9274
rect 5790 9222 5802 9274
rect 5854 9222 5866 9274
rect 5918 9222 5930 9274
rect 5982 9222 15122 9274
rect 15174 9222 15186 9274
rect 15238 9222 15250 9274
rect 15302 9222 15314 9274
rect 15366 9222 15378 9274
rect 15430 9222 24570 9274
rect 24622 9222 24634 9274
rect 24686 9222 24698 9274
rect 24750 9222 24762 9274
rect 24814 9222 24826 9274
rect 24878 9222 34018 9274
rect 34070 9222 34082 9274
rect 34134 9222 34146 9274
rect 34198 9222 34210 9274
rect 34262 9222 34274 9274
rect 34326 9222 38824 9274
rect 1104 9200 38824 9222
rect 2869 9163 2927 9169
rect 2869 9129 2881 9163
rect 2915 9160 2927 9163
rect 22002 9160 22008 9172
rect 2915 9132 3556 9160
rect 21963 9132 22008 9160
rect 2915 9129 2927 9132
rect 2869 9123 2927 9129
rect 2225 9027 2283 9033
rect 2225 9024 2237 9027
rect 1688 8996 2237 9024
rect 1688 8965 1716 8996
rect 2225 8993 2237 8996
rect 2271 9024 2283 9027
rect 2866 9024 2872 9036
rect 2271 8996 2872 9024
rect 2271 8993 2283 8996
rect 2225 8987 2283 8993
rect 2866 8984 2872 8996
rect 2924 8984 2930 9036
rect 3528 9024 3556 9132
rect 22002 9120 22008 9132
rect 22060 9120 22066 9172
rect 22462 9120 22468 9172
rect 22520 9160 22526 9172
rect 22649 9163 22707 9169
rect 22649 9160 22661 9163
rect 22520 9132 22661 9160
rect 22520 9120 22526 9132
rect 22649 9129 22661 9132
rect 22695 9129 22707 9163
rect 22649 9123 22707 9129
rect 22833 9163 22891 9169
rect 22833 9129 22845 9163
rect 22879 9160 22891 9163
rect 24394 9160 24400 9172
rect 22879 9132 24400 9160
rect 22879 9129 22891 9132
rect 22833 9123 22891 9129
rect 24394 9120 24400 9132
rect 24452 9120 24458 9172
rect 26786 9160 26792 9172
rect 24504 9132 26792 9160
rect 3694 9052 3700 9104
rect 3752 9092 3758 9104
rect 3752 9064 22416 9092
rect 3752 9052 3758 9064
rect 3528 8996 3924 9024
rect 1673 8959 1731 8965
rect 1673 8925 1685 8959
rect 1719 8925 1731 8959
rect 1673 8919 1731 8925
rect 2682 8888 2688 8900
rect 2643 8860 2688 8888
rect 2682 8848 2688 8860
rect 2740 8848 2746 8900
rect 3896 8897 3924 8996
rect 4982 8984 4988 9036
rect 5040 9024 5046 9036
rect 21082 9024 21088 9036
rect 5040 8996 21088 9024
rect 5040 8984 5046 8996
rect 21082 8984 21088 8996
rect 21140 8984 21146 9036
rect 6638 8956 6644 8968
rect 6599 8928 6644 8956
rect 6638 8916 6644 8928
rect 6696 8916 6702 8968
rect 17862 8916 17868 8968
rect 17920 8956 17926 8968
rect 20806 8956 20812 8968
rect 17920 8928 20812 8956
rect 17920 8916 17926 8928
rect 20806 8916 20812 8928
rect 20864 8956 20870 8968
rect 20901 8959 20959 8965
rect 20901 8956 20913 8959
rect 20864 8928 20913 8956
rect 20864 8916 20870 8928
rect 20901 8925 20913 8928
rect 20947 8925 20959 8959
rect 20901 8919 20959 8925
rect 22005 8959 22063 8965
rect 22005 8925 22017 8959
rect 22051 8956 22063 8959
rect 22278 8956 22284 8968
rect 22051 8928 22284 8956
rect 22051 8925 22063 8928
rect 22005 8919 22063 8925
rect 3881 8891 3939 8897
rect 3881 8857 3893 8891
rect 3927 8888 3939 8891
rect 13814 8888 13820 8900
rect 3927 8860 13820 8888
rect 3927 8857 3939 8860
rect 3881 8851 3939 8857
rect 13814 8848 13820 8860
rect 13872 8848 13878 8900
rect 20916 8888 20944 8919
rect 22278 8916 22284 8928
rect 22336 8916 22342 8968
rect 22388 8956 22416 9064
rect 22462 8984 22468 9036
rect 22520 9024 22526 9036
rect 23293 9027 23351 9033
rect 23293 9024 23305 9027
rect 22520 8996 23305 9024
rect 22520 8984 22526 8996
rect 23293 8993 23305 8996
rect 23339 8993 23351 9027
rect 23293 8987 23351 8993
rect 24504 8956 24532 9132
rect 26786 9120 26792 9132
rect 26844 9120 26850 9172
rect 31389 9163 31447 9169
rect 26896 9132 30512 9160
rect 26896 9092 26924 9132
rect 26206 9064 26924 9092
rect 30484 9092 30512 9132
rect 31389 9129 31401 9163
rect 31435 9160 31447 9163
rect 31938 9160 31944 9172
rect 31435 9132 31944 9160
rect 31435 9129 31447 9132
rect 31389 9123 31447 9129
rect 31938 9120 31944 9132
rect 31996 9120 32002 9172
rect 31662 9092 31668 9104
rect 30484 9064 31668 9092
rect 22388 8928 22600 8956
rect 22465 8891 22523 8897
rect 22465 8888 22477 8891
rect 20916 8860 22477 8888
rect 22465 8857 22477 8860
rect 22511 8857 22523 8891
rect 22465 8851 22523 8857
rect 1486 8820 1492 8832
rect 1447 8792 1492 8820
rect 1486 8780 1492 8792
rect 1544 8780 1550 8832
rect 2866 8780 2872 8832
rect 2924 8829 2930 8832
rect 2924 8823 2943 8829
rect 2931 8789 2943 8823
rect 2924 8783 2943 8789
rect 3053 8823 3111 8829
rect 3053 8789 3065 8823
rect 3099 8820 3111 8823
rect 3694 8820 3700 8832
rect 3099 8792 3700 8820
rect 3099 8789 3111 8792
rect 3053 8783 3111 8789
rect 2924 8780 2930 8783
rect 3694 8780 3700 8792
rect 3752 8780 3758 8832
rect 6178 8780 6184 8832
rect 6236 8820 6242 8832
rect 6549 8823 6607 8829
rect 6549 8820 6561 8823
rect 6236 8792 6561 8820
rect 6236 8780 6242 8792
rect 6549 8789 6561 8792
rect 6595 8789 6607 8823
rect 7374 8820 7380 8832
rect 7335 8792 7380 8820
rect 6549 8783 6607 8789
rect 7374 8780 7380 8792
rect 7432 8780 7438 8832
rect 8846 8780 8852 8832
rect 8904 8820 8910 8832
rect 20622 8820 20628 8832
rect 8904 8792 20628 8820
rect 8904 8780 8910 8792
rect 20622 8780 20628 8792
rect 20680 8780 20686 8832
rect 22572 8820 22600 8928
rect 23308 8928 24532 8956
rect 22681 8891 22739 8897
rect 22681 8857 22693 8891
rect 22727 8888 22739 8891
rect 23308 8888 23336 8928
rect 24762 8916 24768 8968
rect 24820 8956 24826 8968
rect 26206 8956 26234 9064
rect 31662 9052 31668 9064
rect 31720 9092 31726 9104
rect 32033 9095 32091 9101
rect 32033 9092 32045 9095
rect 31720 9064 32045 9092
rect 31720 9052 31726 9064
rect 32033 9061 32045 9064
rect 32079 9061 32091 9095
rect 32033 9055 32091 9061
rect 27430 8984 27436 9036
rect 27488 9024 27494 9036
rect 27488 8996 27533 9024
rect 27488 8984 27494 8996
rect 27154 8956 27160 8968
rect 24820 8928 26234 8956
rect 27115 8928 27160 8956
rect 24820 8916 24826 8928
rect 27154 8916 27160 8928
rect 27212 8916 27218 8968
rect 30561 8959 30619 8965
rect 30561 8925 30573 8959
rect 30607 8956 30619 8959
rect 30650 8956 30656 8968
rect 30607 8928 30656 8956
rect 30607 8925 30619 8928
rect 30561 8919 30619 8925
rect 30650 8916 30656 8928
rect 30708 8916 30714 8968
rect 31205 8959 31263 8965
rect 31205 8956 31217 8959
rect 30760 8928 31217 8956
rect 22727 8860 23336 8888
rect 22727 8857 22739 8860
rect 22681 8851 22739 8857
rect 24854 8848 24860 8900
rect 24912 8888 24918 8900
rect 30466 8888 30472 8900
rect 24912 8860 30472 8888
rect 24912 8848 24918 8860
rect 30466 8848 30472 8860
rect 30524 8888 30530 8900
rect 30760 8888 30788 8928
rect 31205 8925 31217 8928
rect 31251 8925 31263 8959
rect 31205 8919 31263 8925
rect 30524 8860 30788 8888
rect 30524 8848 30530 8860
rect 26421 8823 26479 8829
rect 26421 8820 26433 8823
rect 22572 8792 26433 8820
rect 26421 8789 26433 8792
rect 26467 8820 26479 8823
rect 28718 8820 28724 8832
rect 26467 8792 28724 8820
rect 26467 8789 26479 8792
rect 26421 8783 26479 8789
rect 28718 8780 28724 8792
rect 28776 8780 28782 8832
rect 30742 8820 30748 8832
rect 30703 8792 30748 8820
rect 30742 8780 30748 8792
rect 30800 8780 30806 8832
rect 1104 8730 38824 8752
rect 1104 8678 10398 8730
rect 10450 8678 10462 8730
rect 10514 8678 10526 8730
rect 10578 8678 10590 8730
rect 10642 8678 10654 8730
rect 10706 8678 19846 8730
rect 19898 8678 19910 8730
rect 19962 8678 19974 8730
rect 20026 8678 20038 8730
rect 20090 8678 20102 8730
rect 20154 8678 29294 8730
rect 29346 8678 29358 8730
rect 29410 8678 29422 8730
rect 29474 8678 29486 8730
rect 29538 8678 29550 8730
rect 29602 8678 38824 8730
rect 1104 8656 38824 8678
rect 2682 8576 2688 8628
rect 2740 8616 2746 8628
rect 4982 8616 4988 8628
rect 2740 8588 4988 8616
rect 2740 8576 2746 8588
rect 2884 8557 2912 8588
rect 4982 8576 4988 8588
rect 5040 8576 5046 8628
rect 7006 8625 7012 8628
rect 6993 8619 7012 8625
rect 6993 8585 7005 8619
rect 7064 8616 7070 8628
rect 8087 8619 8145 8625
rect 8087 8616 8099 8619
rect 7064 8588 8099 8616
rect 6993 8579 7012 8585
rect 7006 8576 7012 8579
rect 7064 8576 7070 8588
rect 8087 8585 8099 8588
rect 8133 8585 8145 8619
rect 8846 8616 8852 8628
rect 8087 8579 8145 8585
rect 8312 8588 8852 8616
rect 2869 8551 2927 8557
rect 2869 8517 2881 8551
rect 2915 8517 2927 8551
rect 2869 8511 2927 8517
rect 2958 8508 2964 8560
rect 3016 8548 3022 8560
rect 3085 8551 3143 8557
rect 3085 8548 3097 8551
rect 3016 8520 3097 8548
rect 3016 8508 3022 8520
rect 3085 8517 3097 8520
rect 3131 8548 3143 8551
rect 7098 8548 7104 8560
rect 3131 8520 7104 8548
rect 3131 8517 3143 8520
rect 3085 8511 3143 8517
rect 7098 8508 7104 8520
rect 7156 8508 7162 8560
rect 7193 8551 7251 8557
rect 7193 8517 7205 8551
rect 7239 8548 7251 8551
rect 7374 8548 7380 8560
rect 7239 8520 7380 8548
rect 7239 8517 7251 8520
rect 7193 8511 7251 8517
rect 7374 8508 7380 8520
rect 7432 8548 7438 8560
rect 8312 8557 8340 8588
rect 8846 8576 8852 8588
rect 8904 8576 8910 8628
rect 9401 8619 9459 8625
rect 9401 8585 9413 8619
rect 9447 8616 9459 8619
rect 18966 8616 18972 8628
rect 9447 8588 18972 8616
rect 9447 8585 9459 8588
rect 9401 8579 9459 8585
rect 8297 8551 8355 8557
rect 8297 8548 8309 8551
rect 7432 8520 8309 8548
rect 7432 8508 7438 8520
rect 8297 8517 8309 8520
rect 8343 8517 8355 8551
rect 8297 8511 8355 8517
rect 3694 8480 3700 8492
rect 3655 8452 3700 8480
rect 3694 8440 3700 8452
rect 3752 8440 3758 8492
rect 4430 8344 4436 8356
rect 3068 8316 4436 8344
rect 3068 8285 3096 8316
rect 4430 8304 4436 8316
rect 4488 8304 4494 8356
rect 6825 8347 6883 8353
rect 6825 8313 6837 8347
rect 6871 8344 6883 8347
rect 6914 8344 6920 8356
rect 6871 8316 6920 8344
rect 6871 8313 6883 8316
rect 6825 8307 6883 8313
rect 6914 8304 6920 8316
rect 6972 8304 6978 8356
rect 7742 8304 7748 8356
rect 7800 8344 7806 8356
rect 7929 8347 7987 8353
rect 7929 8344 7941 8347
rect 7800 8316 7941 8344
rect 7800 8304 7806 8316
rect 7929 8313 7941 8316
rect 7975 8313 7987 8347
rect 9416 8344 9444 8579
rect 18966 8576 18972 8588
rect 19024 8576 19030 8628
rect 19061 8619 19119 8625
rect 19061 8585 19073 8619
rect 19107 8585 19119 8619
rect 19061 8579 19119 8585
rect 19797 8619 19855 8625
rect 19797 8585 19809 8619
rect 19843 8616 19855 8619
rect 30282 8616 30288 8628
rect 19843 8588 30288 8616
rect 19843 8585 19855 8588
rect 19797 8579 19855 8585
rect 13814 8508 13820 8560
rect 13872 8548 13878 8560
rect 19076 8548 19104 8579
rect 13872 8520 19104 8548
rect 13872 8508 13878 8520
rect 10134 8440 10140 8492
rect 10192 8480 10198 8492
rect 13173 8483 13231 8489
rect 13173 8480 13185 8483
rect 10192 8452 13185 8480
rect 10192 8440 10198 8452
rect 13173 8449 13185 8452
rect 13219 8480 13231 8483
rect 13722 8480 13728 8492
rect 13219 8452 13728 8480
rect 13219 8449 13231 8452
rect 13173 8443 13231 8449
rect 13722 8440 13728 8452
rect 13780 8440 13786 8492
rect 17770 8480 17776 8492
rect 17731 8452 17776 8480
rect 17770 8440 17776 8452
rect 17828 8440 17834 8492
rect 19245 8483 19303 8489
rect 19245 8449 19257 8483
rect 19291 8480 19303 8483
rect 19812 8480 19840 8579
rect 30282 8576 30288 8588
rect 30340 8576 30346 8628
rect 30466 8616 30472 8628
rect 30427 8588 30472 8616
rect 30466 8576 30472 8588
rect 30524 8576 30530 8628
rect 31389 8619 31447 8625
rect 31389 8585 31401 8619
rect 31435 8616 31447 8619
rect 34422 8616 34428 8628
rect 31435 8588 34428 8616
rect 31435 8585 31447 8588
rect 31389 8579 31447 8585
rect 34422 8576 34428 8588
rect 34480 8576 34486 8628
rect 20622 8548 20628 8560
rect 20583 8520 20628 8548
rect 20622 8508 20628 8520
rect 20680 8508 20686 8560
rect 20806 8548 20812 8560
rect 20767 8520 20812 8548
rect 20806 8508 20812 8520
rect 20864 8508 20870 8560
rect 21082 8508 21088 8560
rect 21140 8548 21146 8560
rect 23474 8548 23480 8560
rect 21140 8520 23480 8548
rect 21140 8508 21146 8520
rect 23474 8508 23480 8520
rect 23532 8548 23538 8560
rect 23569 8551 23627 8557
rect 23569 8548 23581 8551
rect 23532 8520 23581 8548
rect 23532 8508 23538 8520
rect 23569 8517 23581 8520
rect 23615 8517 23627 8551
rect 23569 8511 23627 8517
rect 23785 8551 23843 8557
rect 23785 8517 23797 8551
rect 23831 8548 23843 8551
rect 30009 8551 30067 8557
rect 23831 8520 29960 8548
rect 23831 8517 23843 8520
rect 23785 8511 23843 8517
rect 22278 8480 22284 8492
rect 19291 8452 19840 8480
rect 22191 8452 22284 8480
rect 19291 8449 19303 8452
rect 19245 8443 19303 8449
rect 17494 8412 17500 8424
rect 17455 8384 17500 8412
rect 17494 8372 17500 8384
rect 17552 8372 17558 8424
rect 7929 8307 7987 8313
rect 8680 8316 9444 8344
rect 18509 8347 18567 8353
rect 3053 8279 3111 8285
rect 3053 8245 3065 8279
rect 3099 8245 3111 8279
rect 3234 8276 3240 8288
rect 3195 8248 3240 8276
rect 3053 8239 3111 8245
rect 3234 8236 3240 8248
rect 3292 8236 3298 8288
rect 3881 8279 3939 8285
rect 3881 8245 3893 8279
rect 3927 8276 3939 8279
rect 4062 8276 4068 8288
rect 3927 8248 4068 8276
rect 3927 8245 3939 8248
rect 3881 8239 3939 8245
rect 4062 8236 4068 8248
rect 4120 8236 4126 8288
rect 7009 8279 7067 8285
rect 7009 8245 7021 8279
rect 7055 8276 7067 8279
rect 7558 8276 7564 8288
rect 7055 8248 7564 8276
rect 7055 8245 7067 8248
rect 7009 8239 7067 8245
rect 7558 8236 7564 8248
rect 7616 8236 7622 8288
rect 8113 8279 8171 8285
rect 8113 8245 8125 8279
rect 8159 8276 8171 8279
rect 8680 8276 8708 8316
rect 18509 8313 18521 8347
rect 18555 8344 18567 8347
rect 19260 8344 19288 8443
rect 22278 8440 22284 8452
rect 22336 8480 22342 8492
rect 22462 8480 22468 8492
rect 22336 8452 22468 8480
rect 22336 8440 22342 8452
rect 22462 8440 22468 8452
rect 22520 8440 22526 8492
rect 23584 8480 23612 8511
rect 24762 8480 24768 8492
rect 23584 8452 24768 8480
rect 24762 8440 24768 8452
rect 24820 8440 24826 8492
rect 26973 8483 27031 8489
rect 26973 8480 26985 8483
rect 26206 8452 26985 8480
rect 20254 8372 20260 8424
rect 20312 8412 20318 8424
rect 22005 8415 22063 8421
rect 22005 8412 22017 8415
rect 20312 8384 22017 8412
rect 20312 8372 20318 8384
rect 22005 8381 22017 8384
rect 22051 8381 22063 8415
rect 24854 8412 24860 8424
rect 22005 8375 22063 8381
rect 23032 8384 24860 8412
rect 23032 8356 23060 8384
rect 24854 8372 24860 8384
rect 24912 8372 24918 8424
rect 23014 8344 23020 8356
rect 18555 8316 19288 8344
rect 22975 8316 23020 8344
rect 18555 8313 18567 8316
rect 18509 8307 18567 8313
rect 23014 8304 23020 8316
rect 23072 8304 23078 8356
rect 23937 8347 23995 8353
rect 23937 8313 23949 8347
rect 23983 8344 23995 8347
rect 26206 8344 26234 8452
rect 26973 8449 26985 8452
rect 27019 8449 27031 8483
rect 27893 8483 27951 8489
rect 27893 8480 27905 8483
rect 26973 8443 27031 8449
rect 27172 8452 27905 8480
rect 27172 8353 27200 8452
rect 27893 8449 27905 8452
rect 27939 8449 27951 8483
rect 29932 8480 29960 8520
rect 30009 8517 30021 8551
rect 30055 8548 30067 8551
rect 30374 8548 30380 8560
rect 30055 8520 30380 8548
rect 30055 8517 30067 8520
rect 30009 8511 30067 8517
rect 30374 8508 30380 8520
rect 30432 8548 30438 8560
rect 31021 8551 31079 8557
rect 31021 8548 31033 8551
rect 30432 8520 31033 8548
rect 30432 8508 30438 8520
rect 31021 8517 31033 8520
rect 31067 8517 31079 8551
rect 31221 8551 31279 8557
rect 31221 8548 31233 8551
rect 31021 8511 31079 8517
rect 31128 8520 31233 8548
rect 30742 8480 30748 8492
rect 29932 8452 30748 8480
rect 27893 8443 27951 8449
rect 30742 8440 30748 8452
rect 30800 8480 30806 8492
rect 31128 8480 31156 8520
rect 31221 8517 31233 8520
rect 31267 8517 31279 8551
rect 31221 8511 31279 8517
rect 31662 8508 31668 8560
rect 31720 8548 31726 8560
rect 32125 8551 32183 8557
rect 32125 8548 32137 8551
rect 31720 8520 32137 8548
rect 31720 8508 31726 8520
rect 32125 8517 32137 8520
rect 32171 8517 32183 8551
rect 32325 8551 32383 8557
rect 32325 8548 32337 8551
rect 32125 8511 32183 8517
rect 32232 8520 32337 8548
rect 32232 8480 32260 8520
rect 32325 8517 32337 8520
rect 32371 8517 32383 8551
rect 32325 8511 32383 8517
rect 30800 8452 32260 8480
rect 30800 8440 30806 8452
rect 27430 8372 27436 8424
rect 27488 8412 27494 8424
rect 27614 8412 27620 8424
rect 27488 8384 27620 8412
rect 27488 8372 27494 8384
rect 27614 8372 27620 8384
rect 27672 8372 27678 8424
rect 28718 8372 28724 8424
rect 28776 8412 28782 8424
rect 33134 8412 33140 8424
rect 28776 8384 33140 8412
rect 28776 8372 28782 8384
rect 33134 8372 33140 8384
rect 33192 8372 33198 8424
rect 23983 8316 26234 8344
rect 27157 8347 27215 8353
rect 23983 8313 23995 8316
rect 23937 8307 23995 8313
rect 27157 8313 27169 8347
rect 27203 8313 27215 8347
rect 27157 8307 27215 8313
rect 28629 8347 28687 8353
rect 28629 8313 28641 8347
rect 28675 8344 28687 8347
rect 28736 8344 28764 8372
rect 28675 8316 28764 8344
rect 28675 8313 28687 8316
rect 28629 8307 28687 8313
rect 30282 8304 30288 8356
rect 30340 8344 30346 8356
rect 32493 8347 32551 8353
rect 30340 8316 32076 8344
rect 30340 8304 30346 8316
rect 32048 8288 32076 8316
rect 32493 8313 32505 8347
rect 32539 8344 32551 8347
rect 33778 8344 33784 8356
rect 32539 8316 33784 8344
rect 32539 8313 32551 8316
rect 32493 8307 32551 8313
rect 33778 8304 33784 8316
rect 33836 8304 33842 8356
rect 13078 8276 13084 8288
rect 8159 8248 8708 8276
rect 13039 8248 13084 8276
rect 8159 8245 8171 8248
rect 8113 8239 8171 8245
rect 13078 8236 13084 8248
rect 13136 8236 13142 8288
rect 23750 8276 23756 8288
rect 23711 8248 23756 8276
rect 23750 8236 23756 8248
rect 23808 8236 23814 8288
rect 30466 8236 30472 8288
rect 30524 8276 30530 8288
rect 31205 8279 31263 8285
rect 31205 8276 31217 8279
rect 30524 8248 31217 8276
rect 30524 8236 30530 8248
rect 31205 8245 31217 8248
rect 31251 8245 31263 8279
rect 31205 8239 31263 8245
rect 32030 8236 32036 8288
rect 32088 8276 32094 8288
rect 32309 8279 32367 8285
rect 32309 8276 32321 8279
rect 32088 8248 32321 8276
rect 32088 8236 32094 8248
rect 32309 8245 32321 8248
rect 32355 8245 32367 8279
rect 32309 8239 32367 8245
rect 1104 8186 38824 8208
rect 1104 8134 5674 8186
rect 5726 8134 5738 8186
rect 5790 8134 5802 8186
rect 5854 8134 5866 8186
rect 5918 8134 5930 8186
rect 5982 8134 15122 8186
rect 15174 8134 15186 8186
rect 15238 8134 15250 8186
rect 15302 8134 15314 8186
rect 15366 8134 15378 8186
rect 15430 8134 24570 8186
rect 24622 8134 24634 8186
rect 24686 8134 24698 8186
rect 24750 8134 24762 8186
rect 24814 8134 24826 8186
rect 24878 8134 34018 8186
rect 34070 8134 34082 8186
rect 34134 8134 34146 8186
rect 34198 8134 34210 8186
rect 34262 8134 34274 8186
rect 34326 8134 38824 8186
rect 1104 8112 38824 8134
rect 6365 8075 6423 8081
rect 6365 8041 6377 8075
rect 6411 8072 6423 8075
rect 7282 8072 7288 8084
rect 6411 8044 7288 8072
rect 6411 8041 6423 8044
rect 6365 8035 6423 8041
rect 7282 8032 7288 8044
rect 7340 8032 7346 8084
rect 23474 8072 23480 8084
rect 23435 8044 23480 8072
rect 23474 8032 23480 8044
rect 23532 8032 23538 8084
rect 31110 8072 31116 8084
rect 31071 8044 31116 8072
rect 31110 8032 31116 8044
rect 31168 8032 31174 8084
rect 31849 8075 31907 8081
rect 31849 8041 31861 8075
rect 31895 8072 31907 8075
rect 32030 8072 32036 8084
rect 31895 8044 32036 8072
rect 31895 8041 31907 8044
rect 31849 8035 31907 8041
rect 32030 8032 32036 8044
rect 32088 8032 32094 8084
rect 27893 8007 27951 8013
rect 27893 7973 27905 8007
rect 27939 8004 27951 8007
rect 32122 8004 32128 8016
rect 27939 7976 32128 8004
rect 27939 7973 27951 7976
rect 27893 7967 27951 7973
rect 32122 7964 32128 7976
rect 32180 7964 32186 8016
rect 9030 7896 9036 7948
rect 9088 7936 9094 7948
rect 9125 7939 9183 7945
rect 9125 7936 9137 7939
rect 9088 7908 9137 7936
rect 9088 7896 9094 7908
rect 9125 7905 9137 7908
rect 9171 7905 9183 7939
rect 11790 7936 11796 7948
rect 11751 7908 11796 7936
rect 9125 7899 9183 7905
rect 11790 7896 11796 7908
rect 11848 7896 11854 7948
rect 13541 7939 13599 7945
rect 13541 7905 13553 7939
rect 13587 7936 13599 7939
rect 18230 7936 18236 7948
rect 13587 7908 18236 7936
rect 13587 7905 13599 7908
rect 13541 7899 13599 7905
rect 18230 7896 18236 7908
rect 18288 7896 18294 7948
rect 3053 7871 3111 7877
rect 3053 7837 3065 7871
rect 3099 7868 3111 7871
rect 3234 7868 3240 7880
rect 3099 7840 3240 7868
rect 3099 7837 3111 7840
rect 3053 7831 3111 7837
rect 3234 7828 3240 7840
rect 3292 7828 3298 7880
rect 3786 7868 3792 7880
rect 3747 7840 3792 7868
rect 3786 7828 3792 7840
rect 3844 7828 3850 7880
rect 4062 7868 4068 7880
rect 4023 7840 4068 7868
rect 4062 7828 4068 7840
rect 4120 7828 4126 7880
rect 13722 7828 13728 7880
rect 13780 7868 13786 7880
rect 14093 7871 14151 7877
rect 14093 7868 14105 7871
rect 13780 7840 14105 7868
rect 13780 7828 13786 7840
rect 14093 7837 14105 7840
rect 14139 7837 14151 7871
rect 14093 7831 14151 7837
rect 27614 7828 27620 7880
rect 27672 7868 27678 7880
rect 27709 7871 27767 7877
rect 27709 7868 27721 7871
rect 27672 7840 27721 7868
rect 27672 7828 27678 7840
rect 27709 7837 27721 7840
rect 27755 7837 27767 7871
rect 30929 7871 30987 7877
rect 30929 7868 30941 7871
rect 27709 7831 27767 7837
rect 30392 7840 30941 7868
rect 3142 7760 3148 7812
rect 3200 7800 3206 7812
rect 6549 7803 6607 7809
rect 3200 7772 4844 7800
rect 3200 7760 3206 7772
rect 3237 7735 3295 7741
rect 3237 7701 3249 7735
rect 3283 7732 3295 7735
rect 3602 7732 3608 7744
rect 3283 7704 3608 7732
rect 3283 7701 3295 7704
rect 3237 7695 3295 7701
rect 3602 7692 3608 7704
rect 3660 7692 3666 7744
rect 4816 7741 4844 7772
rect 6549 7769 6561 7803
rect 6595 7800 6607 7803
rect 7374 7800 7380 7812
rect 6595 7772 7380 7800
rect 6595 7769 6607 7772
rect 6549 7763 6607 7769
rect 7374 7760 7380 7772
rect 7432 7760 7438 7812
rect 9401 7803 9459 7809
rect 9401 7769 9413 7803
rect 9447 7800 9459 7803
rect 9490 7800 9496 7812
rect 9447 7772 9496 7800
rect 9447 7769 9459 7772
rect 9401 7763 9459 7769
rect 9490 7760 9496 7772
rect 9548 7760 9554 7812
rect 9950 7760 9956 7812
rect 10008 7760 10014 7812
rect 12066 7800 12072 7812
rect 12027 7772 12072 7800
rect 12066 7760 12072 7772
rect 12124 7760 12130 7812
rect 13078 7760 13084 7812
rect 13136 7760 13142 7812
rect 18046 7800 18052 7812
rect 13740 7772 18052 7800
rect 4801 7735 4859 7741
rect 4801 7701 4813 7735
rect 4847 7701 4859 7735
rect 4801 7695 4859 7701
rect 6086 7692 6092 7744
rect 6144 7732 6150 7744
rect 6181 7735 6239 7741
rect 6181 7732 6193 7735
rect 6144 7704 6193 7732
rect 6144 7692 6150 7704
rect 6181 7701 6193 7704
rect 6227 7701 6239 7735
rect 6181 7695 6239 7701
rect 6349 7735 6407 7741
rect 6349 7701 6361 7735
rect 6395 7732 6407 7735
rect 7098 7732 7104 7744
rect 6395 7704 7104 7732
rect 6395 7701 6407 7704
rect 6349 7695 6407 7701
rect 7098 7692 7104 7704
rect 7156 7692 7162 7744
rect 7558 7732 7564 7744
rect 7519 7704 7564 7732
rect 7558 7692 7564 7704
rect 7616 7692 7622 7744
rect 10873 7735 10931 7741
rect 10873 7701 10885 7735
rect 10919 7732 10931 7735
rect 13740 7732 13768 7772
rect 18046 7760 18052 7772
rect 18104 7760 18110 7812
rect 10919 7704 13768 7732
rect 10919 7701 10931 7704
rect 10873 7695 10931 7701
rect 14090 7692 14096 7744
rect 14148 7732 14154 7744
rect 14185 7735 14243 7741
rect 14185 7732 14197 7735
rect 14148 7704 14197 7732
rect 14148 7692 14154 7704
rect 14185 7701 14197 7704
rect 14231 7701 14243 7735
rect 14185 7695 14243 7701
rect 30098 7692 30104 7744
rect 30156 7732 30162 7744
rect 30392 7741 30420 7840
rect 30929 7837 30941 7840
rect 30975 7837 30987 7871
rect 33778 7868 33784 7880
rect 33739 7840 33784 7868
rect 30929 7831 30987 7837
rect 33778 7828 33784 7840
rect 33836 7828 33842 7880
rect 34422 7828 34428 7880
rect 34480 7868 34486 7880
rect 34701 7871 34759 7877
rect 34701 7868 34713 7871
rect 34480 7840 34713 7868
rect 34480 7828 34486 7840
rect 34701 7837 34713 7840
rect 34747 7837 34759 7871
rect 34701 7831 34759 7837
rect 35434 7828 35440 7880
rect 35492 7868 35498 7880
rect 35713 7871 35771 7877
rect 35713 7868 35725 7871
rect 35492 7840 35725 7868
rect 35492 7828 35498 7840
rect 35713 7837 35725 7840
rect 35759 7837 35771 7871
rect 35989 7871 36047 7877
rect 35989 7868 36001 7871
rect 35713 7831 35771 7837
rect 35866 7840 36001 7868
rect 30377 7735 30435 7741
rect 30377 7732 30389 7735
rect 30156 7704 30389 7732
rect 30156 7692 30162 7704
rect 30377 7701 30389 7704
rect 30423 7701 30435 7735
rect 33962 7732 33968 7744
rect 33923 7704 33968 7732
rect 30377 7695 30435 7701
rect 33962 7692 33968 7704
rect 34020 7692 34026 7744
rect 34885 7735 34943 7741
rect 34885 7701 34897 7735
rect 34931 7732 34943 7735
rect 35866 7732 35894 7840
rect 35989 7837 36001 7840
rect 36035 7837 36047 7871
rect 35989 7831 36047 7837
rect 36722 7732 36728 7744
rect 34931 7704 35894 7732
rect 36683 7704 36728 7732
rect 34931 7701 34943 7704
rect 34885 7695 34943 7701
rect 36722 7692 36728 7704
rect 36780 7692 36786 7744
rect 1104 7642 38824 7664
rect 1104 7590 10398 7642
rect 10450 7590 10462 7642
rect 10514 7590 10526 7642
rect 10578 7590 10590 7642
rect 10642 7590 10654 7642
rect 10706 7590 19846 7642
rect 19898 7590 19910 7642
rect 19962 7590 19974 7642
rect 20026 7590 20038 7642
rect 20090 7590 20102 7642
rect 20154 7590 29294 7642
rect 29346 7590 29358 7642
rect 29410 7590 29422 7642
rect 29474 7590 29486 7642
rect 29538 7590 29550 7642
rect 29602 7590 38824 7642
rect 1104 7568 38824 7590
rect 7374 7528 7380 7540
rect 7335 7500 7380 7528
rect 7374 7488 7380 7500
rect 7432 7488 7438 7540
rect 9950 7528 9956 7540
rect 9911 7500 9956 7528
rect 9950 7488 9956 7500
rect 10008 7488 10014 7540
rect 11701 7531 11759 7537
rect 11701 7497 11713 7531
rect 11747 7528 11759 7531
rect 11790 7528 11796 7540
rect 11747 7500 11796 7528
rect 11747 7497 11759 7500
rect 11701 7491 11759 7497
rect 11790 7488 11796 7500
rect 11848 7528 11854 7540
rect 12161 7531 12219 7537
rect 12161 7528 12173 7531
rect 11848 7500 12173 7528
rect 11848 7488 11854 7500
rect 12161 7497 12173 7500
rect 12207 7528 12219 7531
rect 12207 7500 12434 7528
rect 12207 7497 12219 7500
rect 12161 7491 12219 7497
rect 1673 7395 1731 7401
rect 1673 7361 1685 7395
rect 1719 7392 1731 7395
rect 2225 7395 2283 7401
rect 2225 7392 2237 7395
rect 1719 7364 2237 7392
rect 1719 7361 1731 7364
rect 1673 7355 1731 7361
rect 2225 7361 2237 7364
rect 2271 7392 2283 7395
rect 9861 7395 9919 7401
rect 2271 7364 2774 7392
rect 2271 7361 2283 7364
rect 2225 7355 2283 7361
rect 2746 7324 2774 7364
rect 9861 7361 9873 7395
rect 9907 7392 9919 7395
rect 10134 7392 10140 7404
rect 9907 7364 10140 7392
rect 9907 7361 9919 7364
rect 9861 7355 9919 7361
rect 10134 7352 10140 7364
rect 10192 7352 10198 7404
rect 12406 7392 12434 7500
rect 30742 7488 30748 7540
rect 30800 7528 30806 7540
rect 30853 7531 30911 7537
rect 30853 7528 30865 7531
rect 30800 7500 30865 7528
rect 30800 7488 30806 7500
rect 30853 7497 30865 7500
rect 30899 7497 30911 7531
rect 36446 7528 36452 7540
rect 36359 7500 36452 7528
rect 30853 7491 30911 7497
rect 36446 7488 36452 7500
rect 36504 7528 36510 7540
rect 36722 7528 36728 7540
rect 36504 7500 36728 7528
rect 36504 7488 36510 7500
rect 36722 7488 36728 7500
rect 36780 7488 36786 7540
rect 17402 7420 17408 7472
rect 17460 7460 17466 7472
rect 23014 7460 23020 7472
rect 17460 7432 23020 7460
rect 17460 7420 17466 7432
rect 23014 7420 23020 7432
rect 23072 7420 23078 7472
rect 30374 7420 30380 7472
rect 30432 7460 30438 7472
rect 30653 7463 30711 7469
rect 30653 7460 30665 7463
rect 30432 7432 30665 7460
rect 30432 7420 30438 7432
rect 30653 7429 30665 7432
rect 30699 7429 30711 7463
rect 30653 7423 30711 7429
rect 12713 7395 12771 7401
rect 12713 7392 12725 7395
rect 12406 7364 12725 7392
rect 12713 7361 12725 7364
rect 12759 7361 12771 7395
rect 12713 7355 12771 7361
rect 14090 7352 14096 7404
rect 14148 7352 14154 7404
rect 18230 7392 18236 7404
rect 18191 7364 18236 7392
rect 18230 7352 18236 7364
rect 18288 7352 18294 7404
rect 33962 7352 33968 7404
rect 34020 7392 34026 7404
rect 35713 7395 35771 7401
rect 35713 7392 35725 7395
rect 34020 7364 35725 7392
rect 34020 7352 34026 7364
rect 35713 7361 35725 7364
rect 35759 7361 35771 7395
rect 35713 7355 35771 7361
rect 12158 7324 12164 7336
rect 2746 7296 12164 7324
rect 12158 7284 12164 7296
rect 12216 7284 12222 7336
rect 12986 7324 12992 7336
rect 12947 7296 12992 7324
rect 12986 7284 12992 7296
rect 13044 7284 13050 7336
rect 14461 7327 14519 7333
rect 14461 7293 14473 7327
rect 14507 7324 14519 7327
rect 17957 7327 18015 7333
rect 17957 7324 17969 7327
rect 14507 7296 17969 7324
rect 14507 7293 14519 7296
rect 14461 7287 14519 7293
rect 17957 7293 17969 7296
rect 18003 7324 18015 7327
rect 22002 7324 22008 7336
rect 18003 7296 22008 7324
rect 18003 7293 18015 7296
rect 17957 7287 18015 7293
rect 22002 7284 22008 7296
rect 22060 7284 22066 7336
rect 35434 7324 35440 7336
rect 35395 7296 35440 7324
rect 35434 7284 35440 7296
rect 35492 7284 35498 7336
rect 17681 7259 17739 7265
rect 17681 7225 17693 7259
rect 17727 7256 17739 7259
rect 17727 7228 18000 7256
rect 17727 7225 17739 7228
rect 17681 7219 17739 7225
rect 17972 7200 18000 7228
rect 1486 7188 1492 7200
rect 1447 7160 1492 7188
rect 1486 7148 1492 7160
rect 1544 7148 1550 7200
rect 6917 7191 6975 7197
rect 6917 7157 6929 7191
rect 6963 7188 6975 7191
rect 7282 7188 7288 7200
rect 6963 7160 7288 7188
rect 6963 7157 6975 7160
rect 6917 7151 6975 7157
rect 7282 7148 7288 7160
rect 7340 7148 7346 7200
rect 17954 7148 17960 7200
rect 18012 7148 18018 7200
rect 18046 7148 18052 7200
rect 18104 7188 18110 7200
rect 30098 7188 30104 7200
rect 18104 7160 18149 7188
rect 30059 7160 30104 7188
rect 18104 7148 18110 7160
rect 30098 7148 30104 7160
rect 30156 7188 30162 7200
rect 30837 7191 30895 7197
rect 30837 7188 30849 7191
rect 30156 7160 30849 7188
rect 30156 7148 30162 7160
rect 30837 7157 30849 7160
rect 30883 7157 30895 7191
rect 30837 7151 30895 7157
rect 31021 7191 31079 7197
rect 31021 7157 31033 7191
rect 31067 7188 31079 7191
rect 32030 7188 32036 7200
rect 31067 7160 32036 7188
rect 31067 7157 31079 7160
rect 31021 7151 31079 7157
rect 32030 7148 32036 7160
rect 32088 7148 32094 7200
rect 1104 7098 38824 7120
rect 1104 7046 5674 7098
rect 5726 7046 5738 7098
rect 5790 7046 5802 7098
rect 5854 7046 5866 7098
rect 5918 7046 5930 7098
rect 5982 7046 15122 7098
rect 15174 7046 15186 7098
rect 15238 7046 15250 7098
rect 15302 7046 15314 7098
rect 15366 7046 15378 7098
rect 15430 7046 24570 7098
rect 24622 7046 24634 7098
rect 24686 7046 24698 7098
rect 24750 7046 24762 7098
rect 24814 7046 24826 7098
rect 24878 7046 34018 7098
rect 34070 7046 34082 7098
rect 34134 7046 34146 7098
rect 34198 7046 34210 7098
rect 34262 7046 34274 7098
rect 34326 7046 38824 7098
rect 1104 7024 38824 7046
rect 12986 6944 12992 6996
rect 13044 6984 13050 6996
rect 25777 6987 25835 6993
rect 25777 6984 25789 6987
rect 13044 6956 25789 6984
rect 13044 6944 13050 6956
rect 25777 6953 25789 6956
rect 25823 6953 25835 6987
rect 25777 6947 25835 6953
rect 30374 6944 30380 6996
rect 30432 6984 30438 6996
rect 30469 6987 30527 6993
rect 30469 6984 30481 6987
rect 30432 6956 30481 6984
rect 30432 6944 30438 6956
rect 30469 6953 30481 6956
rect 30515 6953 30527 6987
rect 30469 6947 30527 6953
rect 30834 6944 30840 6996
rect 30892 6984 30898 6996
rect 31389 6987 31447 6993
rect 31389 6984 31401 6987
rect 30892 6956 31401 6984
rect 30892 6944 30898 6956
rect 31389 6953 31401 6956
rect 31435 6984 31447 6987
rect 31478 6984 31484 6996
rect 31435 6956 31484 6984
rect 31435 6953 31447 6956
rect 31389 6947 31447 6953
rect 31478 6944 31484 6956
rect 31536 6944 31542 6996
rect 7558 6876 7564 6928
rect 7616 6916 7622 6928
rect 17402 6916 17408 6928
rect 7616 6888 17408 6916
rect 7616 6876 7622 6888
rect 17402 6876 17408 6888
rect 17460 6876 17466 6928
rect 17494 6876 17500 6928
rect 17552 6916 17558 6928
rect 19702 6916 19708 6928
rect 17552 6888 19708 6916
rect 17552 6876 17558 6888
rect 19702 6876 19708 6888
rect 19760 6876 19766 6928
rect 18046 6808 18052 6860
rect 18104 6848 18110 6860
rect 19245 6851 19303 6857
rect 19245 6848 19257 6851
rect 18104 6820 19257 6848
rect 18104 6808 18110 6820
rect 19245 6817 19257 6820
rect 19291 6817 19303 6851
rect 19245 6811 19303 6817
rect 6914 6780 6920 6792
rect 6875 6752 6920 6780
rect 6914 6740 6920 6752
rect 6972 6740 6978 6792
rect 17954 6780 17960 6792
rect 17915 6752 17960 6780
rect 17954 6740 17960 6752
rect 18012 6740 18018 6792
rect 18417 6783 18475 6789
rect 18417 6749 18429 6783
rect 18463 6749 18475 6783
rect 19518 6780 19524 6792
rect 19479 6752 19524 6780
rect 18417 6743 18475 6749
rect 18432 6712 18460 6743
rect 19518 6740 19524 6752
rect 19576 6740 19582 6792
rect 26510 6780 26516 6792
rect 26471 6752 26516 6780
rect 26510 6740 26516 6752
rect 26568 6740 26574 6792
rect 26789 6783 26847 6789
rect 26789 6749 26801 6783
rect 26835 6780 26847 6783
rect 26878 6780 26884 6792
rect 26835 6752 26884 6780
rect 26835 6749 26847 6752
rect 26789 6743 26847 6749
rect 26878 6740 26884 6752
rect 26936 6740 26942 6792
rect 31662 6780 31668 6792
rect 31220 6752 31668 6780
rect 31220 6721 31248 6752
rect 31662 6740 31668 6752
rect 31720 6740 31726 6792
rect 32030 6780 32036 6792
rect 31991 6752 32036 6780
rect 32030 6740 32036 6752
rect 32088 6740 32094 6792
rect 34701 6783 34759 6789
rect 34701 6749 34713 6783
rect 34747 6749 34759 6783
rect 34701 6743 34759 6749
rect 17788 6684 18460 6712
rect 31205 6715 31263 6721
rect 17788 6656 17816 6684
rect 31205 6681 31217 6715
rect 31251 6681 31263 6715
rect 34716 6712 34744 6743
rect 31205 6675 31263 6681
rect 31588 6684 34744 6712
rect 6638 6604 6644 6656
rect 6696 6644 6702 6656
rect 6733 6647 6791 6653
rect 6733 6644 6745 6647
rect 6696 6616 6745 6644
rect 6696 6604 6702 6616
rect 6733 6613 6745 6616
rect 6779 6613 6791 6647
rect 17770 6644 17776 6656
rect 17731 6616 17776 6644
rect 6733 6607 6791 6613
rect 17770 6604 17776 6616
rect 17828 6604 17834 6656
rect 18322 6604 18328 6656
rect 18380 6644 18386 6656
rect 18509 6647 18567 6653
rect 18509 6644 18521 6647
rect 18380 6616 18521 6644
rect 18380 6604 18386 6616
rect 18509 6613 18521 6616
rect 18555 6613 18567 6647
rect 18509 6607 18567 6613
rect 30742 6604 30748 6656
rect 30800 6644 30806 6656
rect 31588 6653 31616 6684
rect 31405 6647 31463 6653
rect 31405 6644 31417 6647
rect 30800 6616 31417 6644
rect 30800 6604 30806 6616
rect 31405 6613 31417 6616
rect 31451 6613 31463 6647
rect 31405 6607 31463 6613
rect 31573 6647 31631 6653
rect 31573 6613 31585 6647
rect 31619 6613 31631 6647
rect 31573 6607 31631 6613
rect 32217 6647 32275 6653
rect 32217 6613 32229 6647
rect 32263 6644 32275 6647
rect 32398 6644 32404 6656
rect 32263 6616 32404 6644
rect 32263 6613 32275 6616
rect 32217 6607 32275 6613
rect 32398 6604 32404 6616
rect 32456 6604 32462 6656
rect 34882 6644 34888 6656
rect 34843 6616 34888 6644
rect 34882 6604 34888 6616
rect 34940 6604 34946 6656
rect 1104 6554 38824 6576
rect 1104 6502 10398 6554
rect 10450 6502 10462 6554
rect 10514 6502 10526 6554
rect 10578 6502 10590 6554
rect 10642 6502 10654 6554
rect 10706 6502 19846 6554
rect 19898 6502 19910 6554
rect 19962 6502 19974 6554
rect 20026 6502 20038 6554
rect 20090 6502 20102 6554
rect 20154 6502 29294 6554
rect 29346 6502 29358 6554
rect 29410 6502 29422 6554
rect 29474 6502 29486 6554
rect 29538 6502 29550 6554
rect 29602 6502 38824 6554
rect 1104 6480 38824 6502
rect 31481 6443 31539 6449
rect 31481 6409 31493 6443
rect 31527 6440 31539 6443
rect 31662 6440 31668 6452
rect 31527 6412 31668 6440
rect 31527 6409 31539 6412
rect 31481 6403 31539 6409
rect 31662 6400 31668 6412
rect 31720 6400 31726 6452
rect 33134 6440 33140 6452
rect 33047 6412 33140 6440
rect 33134 6400 33140 6412
rect 33192 6440 33198 6452
rect 36446 6440 36452 6452
rect 33192 6412 36452 6440
rect 33192 6400 33198 6412
rect 36446 6400 36452 6412
rect 36504 6400 36510 6452
rect 3786 6332 3792 6384
rect 3844 6372 3850 6384
rect 3844 6344 3924 6372
rect 3844 6332 3850 6344
rect 1578 6264 1584 6316
rect 1636 6304 1642 6316
rect 1673 6307 1731 6313
rect 1673 6304 1685 6307
rect 1636 6276 1685 6304
rect 1636 6264 1642 6276
rect 1673 6273 1685 6276
rect 1719 6304 1731 6307
rect 2133 6307 2191 6313
rect 2133 6304 2145 6307
rect 1719 6276 2145 6304
rect 1719 6273 1731 6276
rect 1673 6267 1731 6273
rect 2133 6273 2145 6276
rect 2179 6273 2191 6307
rect 3602 6304 3608 6316
rect 3563 6276 3608 6304
rect 2133 6267 2191 6273
rect 3602 6264 3608 6276
rect 3660 6264 3666 6316
rect 3896 6313 3924 6344
rect 18230 6332 18236 6384
rect 18288 6372 18294 6384
rect 18969 6375 19027 6381
rect 18969 6372 18981 6375
rect 18288 6344 18981 6372
rect 18288 6332 18294 6344
rect 18969 6341 18981 6344
rect 19015 6341 19027 6375
rect 18969 6335 19027 6341
rect 32140 6344 33824 6372
rect 32140 6316 32168 6344
rect 3881 6307 3939 6313
rect 3881 6273 3893 6307
rect 3927 6304 3939 6307
rect 6178 6304 6184 6316
rect 3927 6276 6184 6304
rect 3927 6273 3939 6276
rect 3881 6267 3939 6273
rect 6178 6264 6184 6276
rect 6236 6264 6242 6316
rect 32122 6304 32128 6316
rect 32083 6276 32128 6304
rect 32122 6264 32128 6276
rect 32180 6264 32186 6316
rect 32398 6304 32404 6316
rect 32359 6276 32404 6304
rect 32398 6264 32404 6276
rect 32456 6264 32462 6316
rect 33796 6236 33824 6344
rect 34882 6264 34888 6316
rect 34940 6304 34946 6316
rect 35713 6307 35771 6313
rect 35713 6304 35725 6307
rect 34940 6276 35725 6304
rect 34940 6264 34946 6276
rect 35713 6273 35725 6276
rect 35759 6273 35771 6307
rect 35713 6267 35771 6273
rect 35434 6236 35440 6248
rect 33796 6208 35440 6236
rect 35434 6196 35440 6208
rect 35492 6196 35498 6248
rect 19153 6171 19211 6177
rect 19153 6137 19165 6171
rect 19199 6168 19211 6171
rect 20530 6168 20536 6180
rect 19199 6140 20536 6168
rect 19199 6137 19211 6140
rect 19153 6131 19211 6137
rect 20530 6128 20536 6140
rect 20588 6128 20594 6180
rect 1486 6100 1492 6112
rect 1447 6072 1492 6100
rect 1486 6060 1492 6072
rect 1544 6060 1550 6112
rect 2869 6103 2927 6109
rect 2869 6069 2881 6103
rect 2915 6100 2927 6103
rect 3142 6100 3148 6112
rect 2915 6072 3148 6100
rect 2915 6069 2927 6072
rect 2869 6063 2927 6069
rect 3142 6060 3148 6072
rect 3200 6060 3206 6112
rect 30834 6100 30840 6112
rect 30795 6072 30840 6100
rect 30834 6060 30840 6072
rect 30892 6060 30898 6112
rect 1104 6010 38824 6032
rect 1104 5958 5674 6010
rect 5726 5958 5738 6010
rect 5790 5958 5802 6010
rect 5854 5958 5866 6010
rect 5918 5958 5930 6010
rect 5982 5958 15122 6010
rect 15174 5958 15186 6010
rect 15238 5958 15250 6010
rect 15302 5958 15314 6010
rect 15366 5958 15378 6010
rect 15430 5958 24570 6010
rect 24622 5958 24634 6010
rect 24686 5958 24698 6010
rect 24750 5958 24762 6010
rect 24814 5958 24826 6010
rect 24878 5958 34018 6010
rect 34070 5958 34082 6010
rect 34134 5958 34146 6010
rect 34198 5958 34210 6010
rect 34262 5958 34274 6010
rect 34326 5958 38824 6010
rect 1104 5936 38824 5958
rect 7282 5856 7288 5908
rect 7340 5896 7346 5908
rect 28353 5899 28411 5905
rect 28353 5896 28365 5899
rect 7340 5868 28365 5896
rect 7340 5856 7346 5868
rect 28353 5865 28365 5868
rect 28399 5896 28411 5899
rect 30098 5896 30104 5908
rect 28399 5868 30104 5896
rect 28399 5865 28411 5868
rect 28353 5859 28411 5865
rect 30098 5856 30104 5868
rect 30156 5856 30162 5908
rect 19702 5788 19708 5840
rect 19760 5828 19766 5840
rect 19981 5831 20039 5837
rect 19981 5828 19993 5831
rect 19760 5800 19993 5828
rect 19760 5788 19766 5800
rect 19981 5797 19993 5800
rect 20027 5797 20039 5831
rect 23198 5828 23204 5840
rect 23159 5800 23204 5828
rect 19981 5791 20039 5797
rect 23198 5788 23204 5800
rect 23256 5788 23262 5840
rect 22002 5720 22008 5772
rect 22060 5760 22066 5772
rect 22465 5763 22523 5769
rect 22465 5760 22477 5763
rect 22060 5732 22477 5760
rect 22060 5720 22066 5732
rect 22465 5729 22477 5732
rect 22511 5760 22523 5763
rect 22925 5763 22983 5769
rect 22925 5760 22937 5763
rect 22511 5732 22937 5760
rect 22511 5729 22523 5732
rect 22465 5723 22523 5729
rect 22925 5729 22937 5732
rect 22971 5729 22983 5763
rect 22925 5723 22983 5729
rect 6178 5692 6184 5704
rect 6139 5664 6184 5692
rect 6178 5652 6184 5664
rect 6236 5652 6242 5704
rect 20165 5695 20223 5701
rect 20165 5661 20177 5695
rect 20211 5692 20223 5695
rect 20254 5692 20260 5704
rect 20211 5664 20260 5692
rect 20211 5661 20223 5664
rect 20165 5655 20223 5661
rect 20254 5652 20260 5664
rect 20312 5652 20318 5704
rect 22189 5695 22247 5701
rect 22189 5661 22201 5695
rect 22235 5692 22247 5695
rect 22370 5692 22376 5704
rect 22235 5664 22376 5692
rect 22235 5661 22247 5664
rect 22189 5655 22247 5661
rect 22370 5652 22376 5664
rect 22428 5652 22434 5704
rect 26878 5652 26884 5704
rect 26936 5692 26942 5704
rect 27341 5695 27399 5701
rect 27341 5692 27353 5695
rect 26936 5664 27353 5692
rect 26936 5652 26942 5664
rect 27341 5661 27353 5664
rect 27387 5661 27399 5695
rect 27614 5692 27620 5704
rect 27575 5664 27620 5692
rect 27341 5655 27399 5661
rect 27614 5652 27620 5664
rect 27672 5652 27678 5704
rect 6362 5556 6368 5568
rect 6323 5528 6368 5556
rect 6362 5516 6368 5528
rect 6420 5516 6426 5568
rect 23385 5559 23443 5565
rect 23385 5525 23397 5559
rect 23431 5556 23443 5559
rect 28534 5556 28540 5568
rect 23431 5528 28540 5556
rect 23431 5525 23443 5528
rect 23385 5519 23443 5525
rect 28534 5516 28540 5528
rect 28592 5516 28598 5568
rect 1104 5466 38824 5488
rect 1104 5414 10398 5466
rect 10450 5414 10462 5466
rect 10514 5414 10526 5466
rect 10578 5414 10590 5466
rect 10642 5414 10654 5466
rect 10706 5414 19846 5466
rect 19898 5414 19910 5466
rect 19962 5414 19974 5466
rect 20026 5414 20038 5466
rect 20090 5414 20102 5466
rect 20154 5414 29294 5466
rect 29346 5414 29358 5466
rect 29410 5414 29422 5466
rect 29474 5414 29486 5466
rect 29538 5414 29550 5466
rect 29602 5414 38824 5466
rect 1104 5392 38824 5414
rect 22462 5352 22468 5364
rect 22423 5324 22468 5352
rect 22462 5312 22468 5324
rect 22520 5312 22526 5364
rect 26510 5312 26516 5364
rect 26568 5352 26574 5364
rect 26973 5355 27031 5361
rect 26973 5352 26985 5355
rect 26568 5324 26985 5352
rect 26568 5312 26574 5324
rect 26973 5321 26985 5324
rect 27019 5321 27031 5355
rect 26973 5315 27031 5321
rect 19426 5284 19432 5296
rect 19339 5256 19432 5284
rect 19426 5244 19432 5256
rect 19484 5284 19490 5296
rect 20254 5284 20260 5296
rect 19484 5256 20260 5284
rect 19484 5244 19490 5256
rect 20254 5244 20260 5256
rect 20312 5244 20318 5296
rect 6178 5176 6184 5228
rect 6236 5216 6242 5228
rect 6365 5219 6423 5225
rect 6365 5216 6377 5219
rect 6236 5188 6377 5216
rect 6236 5176 6242 5188
rect 6365 5185 6377 5188
rect 6411 5185 6423 5219
rect 6638 5216 6644 5228
rect 6599 5188 6644 5216
rect 6365 5179 6423 5185
rect 6638 5176 6644 5188
rect 6696 5176 6702 5228
rect 20070 5216 20076 5228
rect 20031 5188 20076 5216
rect 20070 5176 20076 5188
rect 20128 5176 20134 5228
rect 20441 5219 20499 5225
rect 20441 5185 20453 5219
rect 20487 5216 20499 5219
rect 20530 5216 20536 5228
rect 20487 5188 20536 5216
rect 20487 5185 20499 5188
rect 20441 5179 20499 5185
rect 20530 5176 20536 5188
rect 20588 5176 20594 5228
rect 22370 5216 22376 5228
rect 22331 5188 22376 5216
rect 22370 5176 22376 5188
rect 22428 5176 22434 5228
rect 22554 5216 22560 5228
rect 22515 5188 22560 5216
rect 22554 5176 22560 5188
rect 22612 5176 22618 5228
rect 27154 5216 27160 5228
rect 27115 5188 27160 5216
rect 27154 5176 27160 5188
rect 27212 5176 27218 5228
rect 19518 5108 19524 5160
rect 19576 5148 19582 5160
rect 20254 5148 20260 5160
rect 19576 5120 20260 5148
rect 19576 5108 19582 5120
rect 20254 5108 20260 5120
rect 20312 5108 20318 5160
rect 19613 5083 19671 5089
rect 19613 5049 19625 5083
rect 19659 5080 19671 5083
rect 24394 5080 24400 5092
rect 19659 5052 24400 5080
rect 19659 5049 19671 5052
rect 19613 5043 19671 5049
rect 24394 5040 24400 5052
rect 24452 5040 24458 5092
rect 7377 5015 7435 5021
rect 7377 4981 7389 5015
rect 7423 5012 7435 5015
rect 7466 5012 7472 5024
rect 7423 4984 7472 5012
rect 7423 4981 7435 4984
rect 7377 4975 7435 4981
rect 7466 4972 7472 4984
rect 7524 4972 7530 5024
rect 20162 5012 20168 5024
rect 20123 4984 20168 5012
rect 20162 4972 20168 4984
rect 20220 4972 20226 5024
rect 1104 4922 38824 4944
rect 1104 4870 5674 4922
rect 5726 4870 5738 4922
rect 5790 4870 5802 4922
rect 5854 4870 5866 4922
rect 5918 4870 5930 4922
rect 5982 4870 15122 4922
rect 15174 4870 15186 4922
rect 15238 4870 15250 4922
rect 15302 4870 15314 4922
rect 15366 4870 15378 4922
rect 15430 4870 24570 4922
rect 24622 4870 24634 4922
rect 24686 4870 24698 4922
rect 24750 4870 24762 4922
rect 24814 4870 24826 4922
rect 24878 4870 34018 4922
rect 34070 4870 34082 4922
rect 34134 4870 34146 4922
rect 34198 4870 34210 4922
rect 34262 4870 34274 4922
rect 34326 4870 38824 4922
rect 1104 4848 38824 4870
rect 2866 4808 2872 4820
rect 2779 4780 2872 4808
rect 2866 4768 2872 4780
rect 2924 4808 2930 4820
rect 4246 4808 4252 4820
rect 2924 4780 4252 4808
rect 2924 4768 2930 4780
rect 4246 4768 4252 4780
rect 4304 4768 4310 4820
rect 19426 4808 19432 4820
rect 19387 4780 19432 4808
rect 19426 4768 19432 4780
rect 19484 4768 19490 4820
rect 20254 4808 20260 4820
rect 20215 4780 20260 4808
rect 20254 4768 20260 4780
rect 20312 4768 20318 4820
rect 22554 4768 22560 4820
rect 22612 4808 22618 4820
rect 22925 4811 22983 4817
rect 22925 4808 22937 4811
rect 22612 4780 22937 4808
rect 22612 4768 22618 4780
rect 22925 4777 22937 4780
rect 22971 4808 22983 4811
rect 22971 4780 26234 4808
rect 22971 4777 22983 4780
rect 22925 4771 22983 4777
rect 19981 4743 20039 4749
rect 19981 4740 19993 4743
rect 16546 4712 19993 4740
rect 15120 4644 15792 4672
rect 1673 4607 1731 4613
rect 1673 4573 1685 4607
rect 1719 4604 1731 4607
rect 3142 4604 3148 4616
rect 1719 4576 3148 4604
rect 1719 4573 1731 4576
rect 1673 4567 1731 4573
rect 3142 4564 3148 4576
rect 3200 4564 3206 4616
rect 6086 4604 6092 4616
rect 6047 4576 6092 4604
rect 6086 4564 6092 4576
rect 6144 4564 6150 4616
rect 7742 4604 7748 4616
rect 7703 4576 7748 4604
rect 7742 4564 7748 4576
rect 7800 4564 7806 4616
rect 14826 4604 14832 4616
rect 14787 4576 14832 4604
rect 14826 4564 14832 4576
rect 14884 4564 14890 4616
rect 15120 4613 15148 4644
rect 15764 4613 15792 4644
rect 15105 4607 15163 4613
rect 15105 4573 15117 4607
rect 15151 4573 15163 4607
rect 15105 4567 15163 4573
rect 15565 4607 15623 4613
rect 15565 4573 15577 4607
rect 15611 4573 15623 4607
rect 15565 4567 15623 4573
rect 15749 4607 15807 4613
rect 15749 4573 15761 4607
rect 15795 4604 15807 4607
rect 16546 4604 16574 4712
rect 19981 4709 19993 4712
rect 20027 4709 20039 4743
rect 19981 4703 20039 4709
rect 20272 4672 20300 4768
rect 26206 4740 26234 4780
rect 26789 4743 26847 4749
rect 26789 4740 26801 4743
rect 26206 4712 26801 4740
rect 26789 4709 26801 4712
rect 26835 4740 26847 4743
rect 31846 4740 31852 4752
rect 26835 4712 31852 4740
rect 26835 4709 26847 4712
rect 26789 4703 26847 4709
rect 31846 4700 31852 4712
rect 31904 4700 31910 4752
rect 22557 4675 22615 4681
rect 22557 4672 22569 4675
rect 20272 4644 22569 4672
rect 22557 4641 22569 4644
rect 22603 4672 22615 4675
rect 23198 4672 23204 4684
rect 22603 4644 23204 4672
rect 22603 4641 22615 4644
rect 22557 4635 22615 4641
rect 23198 4632 23204 4644
rect 23256 4632 23262 4684
rect 28169 4675 28227 4681
rect 28169 4672 28181 4675
rect 27632 4644 28181 4672
rect 27632 4616 27660 4644
rect 28169 4641 28181 4644
rect 28215 4641 28227 4675
rect 28169 4635 28227 4641
rect 15795 4576 16574 4604
rect 19521 4607 19579 4613
rect 15795 4573 15807 4576
rect 15749 4567 15807 4573
rect 19521 4573 19533 4607
rect 19567 4604 19579 4607
rect 20162 4604 20168 4616
rect 19567 4576 20168 4604
rect 19567 4573 19579 4576
rect 19521 4567 19579 4573
rect 15013 4539 15071 4545
rect 15013 4505 15025 4539
rect 15059 4536 15071 4539
rect 15580 4536 15608 4567
rect 19536 4536 19564 4567
rect 20162 4564 20168 4576
rect 20220 4564 20226 4616
rect 20257 4607 20315 4613
rect 20257 4573 20269 4607
rect 20303 4573 20315 4607
rect 20257 4567 20315 4573
rect 20349 4607 20407 4613
rect 20349 4573 20361 4607
rect 20395 4604 20407 4607
rect 20530 4604 20536 4616
rect 20395 4576 20536 4604
rect 20395 4573 20407 4576
rect 20349 4567 20407 4573
rect 15059 4508 19564 4536
rect 15059 4505 15071 4508
rect 15013 4499 15071 4505
rect 20070 4496 20076 4548
rect 20128 4536 20134 4548
rect 20272 4536 20300 4567
rect 20530 4564 20536 4576
rect 20588 4604 20594 4616
rect 26697 4607 26755 4613
rect 26697 4604 26709 4607
rect 20588 4576 26709 4604
rect 20588 4564 20594 4576
rect 26697 4573 26709 4576
rect 26743 4604 26755 4607
rect 27614 4604 27620 4616
rect 26743 4576 27476 4604
rect 27575 4576 27620 4604
rect 26743 4573 26755 4576
rect 26697 4567 26755 4573
rect 20438 4536 20444 4548
rect 20128 4508 20444 4536
rect 20128 4496 20134 4508
rect 20438 4496 20444 4508
rect 20496 4536 20502 4548
rect 22370 4536 22376 4548
rect 20496 4508 22376 4536
rect 20496 4496 20502 4508
rect 22370 4496 22376 4508
rect 22428 4536 22434 4548
rect 22925 4539 22983 4545
rect 22925 4536 22937 4539
rect 22428 4508 22937 4536
rect 22428 4496 22434 4508
rect 22925 4505 22937 4508
rect 22971 4505 22983 4539
rect 27338 4536 27344 4548
rect 27299 4508 27344 4536
rect 22925 4499 22983 4505
rect 27338 4496 27344 4508
rect 27396 4496 27402 4548
rect 27448 4536 27476 4576
rect 27614 4564 27620 4576
rect 27672 4564 27678 4616
rect 28077 4607 28135 4613
rect 28077 4573 28089 4607
rect 28123 4573 28135 4607
rect 28077 4567 28135 4573
rect 28261 4607 28319 4613
rect 28261 4573 28273 4607
rect 28307 4604 28319 4607
rect 28534 4604 28540 4616
rect 28307 4576 28540 4604
rect 28307 4573 28319 4576
rect 28261 4567 28319 4573
rect 28092 4536 28120 4567
rect 28534 4564 28540 4576
rect 28592 4564 28598 4616
rect 27448 4508 28120 4536
rect 27632 4480 27660 4508
rect 1486 4468 1492 4480
rect 1447 4440 1492 4468
rect 1486 4428 1492 4440
rect 1544 4428 1550 4480
rect 5534 4428 5540 4480
rect 5592 4468 5598 4480
rect 5905 4471 5963 4477
rect 5905 4468 5917 4471
rect 5592 4440 5917 4468
rect 5592 4428 5598 4440
rect 5905 4437 5917 4440
rect 5951 4437 5963 4471
rect 7558 4468 7564 4480
rect 7519 4440 7564 4468
rect 5905 4431 5963 4437
rect 7558 4428 7564 4440
rect 7616 4428 7622 4480
rect 14274 4428 14280 4480
rect 14332 4468 14338 4480
rect 14645 4471 14703 4477
rect 14645 4468 14657 4471
rect 14332 4440 14657 4468
rect 14332 4428 14338 4440
rect 14645 4437 14657 4440
rect 14691 4437 14703 4471
rect 15562 4468 15568 4480
rect 15523 4440 15568 4468
rect 14645 4431 14703 4437
rect 15562 4428 15568 4440
rect 15620 4428 15626 4480
rect 23109 4471 23167 4477
rect 23109 4437 23121 4471
rect 23155 4468 23167 4471
rect 23474 4468 23480 4480
rect 23155 4440 23480 4468
rect 23155 4437 23167 4440
rect 23109 4431 23167 4437
rect 23474 4428 23480 4440
rect 23532 4428 23538 4480
rect 27614 4428 27620 4480
rect 27672 4428 27678 4480
rect 1104 4378 38824 4400
rect 1104 4326 10398 4378
rect 10450 4326 10462 4378
rect 10514 4326 10526 4378
rect 10578 4326 10590 4378
rect 10642 4326 10654 4378
rect 10706 4326 19846 4378
rect 19898 4326 19910 4378
rect 19962 4326 19974 4378
rect 20026 4326 20038 4378
rect 20090 4326 20102 4378
rect 20154 4326 29294 4378
rect 29346 4326 29358 4378
rect 29410 4326 29422 4378
rect 29474 4326 29486 4378
rect 29538 4326 29550 4378
rect 29602 4326 38824 4378
rect 1104 4304 38824 4326
rect 3142 4264 3148 4276
rect 3055 4236 3148 4264
rect 3142 4224 3148 4236
rect 3200 4264 3206 4276
rect 4062 4264 4068 4276
rect 3200 4236 4068 4264
rect 3200 4224 3206 4236
rect 4062 4224 4068 4236
rect 4120 4224 4126 4276
rect 7466 4264 7472 4276
rect 7427 4236 7472 4264
rect 7466 4224 7472 4236
rect 7524 4224 7530 4276
rect 27154 4224 27160 4276
rect 27212 4264 27218 4276
rect 27249 4267 27307 4273
rect 27249 4264 27261 4267
rect 27212 4236 27261 4264
rect 27212 4224 27218 4236
rect 27249 4233 27261 4236
rect 27295 4233 27307 4267
rect 27249 4227 27307 4233
rect 27417 4267 27475 4273
rect 27417 4233 27429 4267
rect 27463 4264 27475 4267
rect 27522 4264 27528 4276
rect 27463 4236 27528 4264
rect 27463 4233 27475 4236
rect 27417 4227 27475 4233
rect 27522 4224 27528 4236
rect 27580 4224 27586 4276
rect 19613 4199 19671 4205
rect 5368 4168 5672 4196
rect 2501 4131 2559 4137
rect 2501 4097 2513 4131
rect 2547 4128 2559 4131
rect 3881 4131 3939 4137
rect 2547 4100 3556 4128
rect 2547 4097 2559 4100
rect 2501 4091 2559 4097
rect 2317 4063 2375 4069
rect 2317 4029 2329 4063
rect 2363 4060 2375 4063
rect 2866 4060 2872 4072
rect 2363 4032 2872 4060
rect 2363 4029 2375 4032
rect 2317 4023 2375 4029
rect 2866 4020 2872 4032
rect 2924 4020 2930 4072
rect 2685 3927 2743 3933
rect 2685 3893 2697 3927
rect 2731 3924 2743 3927
rect 2866 3924 2872 3936
rect 2731 3896 2872 3924
rect 2731 3893 2743 3896
rect 2685 3887 2743 3893
rect 2866 3884 2872 3896
rect 2924 3884 2930 3936
rect 3528 3924 3556 4100
rect 3881 4097 3893 4131
rect 3927 4128 3939 4131
rect 4706 4128 4712 4140
rect 3927 4100 4712 4128
rect 3927 4097 3939 4100
rect 3881 4091 3939 4097
rect 4706 4088 4712 4100
rect 4764 4088 4770 4140
rect 5368 4128 5396 4168
rect 5534 4128 5540 4140
rect 5092 4100 5396 4128
rect 5495 4100 5540 4128
rect 4157 4063 4215 4069
rect 4157 4029 4169 4063
rect 4203 4060 4215 4063
rect 5092 4060 5120 4100
rect 5534 4088 5540 4100
rect 5592 4088 5598 4140
rect 5644 4128 5672 4168
rect 14108 4168 14412 4196
rect 5813 4131 5871 4137
rect 5813 4128 5825 4131
rect 5644 4100 5825 4128
rect 5813 4097 5825 4100
rect 5859 4128 5871 4131
rect 6362 4128 6368 4140
rect 5859 4100 6368 4128
rect 5859 4097 5871 4100
rect 5813 4091 5871 4097
rect 6362 4088 6368 4100
rect 6420 4128 6426 4140
rect 6457 4131 6515 4137
rect 6457 4128 6469 4131
rect 6420 4100 6469 4128
rect 6420 4088 6426 4100
rect 6457 4097 6469 4100
rect 6503 4097 6515 4131
rect 6457 4091 6515 4097
rect 6733 4131 6791 4137
rect 6733 4097 6745 4131
rect 6779 4128 6791 4131
rect 7558 4128 7564 4140
rect 6779 4100 7564 4128
rect 6779 4097 6791 4100
rect 6733 4091 6791 4097
rect 7558 4088 7564 4100
rect 7616 4088 7622 4140
rect 10229 4131 10287 4137
rect 10229 4097 10241 4131
rect 10275 4128 10287 4131
rect 11974 4128 11980 4140
rect 10275 4100 11980 4128
rect 10275 4097 10287 4100
rect 10229 4091 10287 4097
rect 11974 4088 11980 4100
rect 12032 4088 12038 4140
rect 14001 4131 14059 4137
rect 14001 4097 14013 4131
rect 14047 4128 14059 4131
rect 14108 4128 14136 4168
rect 14384 4140 14412 4168
rect 19613 4165 19625 4199
rect 19659 4196 19671 4199
rect 23750 4196 23756 4208
rect 19659 4168 23756 4196
rect 19659 4165 19671 4168
rect 19613 4159 19671 4165
rect 14274 4128 14280 4140
rect 14047 4100 14136 4128
rect 14235 4100 14280 4128
rect 14047 4097 14059 4100
rect 14001 4091 14059 4097
rect 14274 4088 14280 4100
rect 14332 4088 14338 4140
rect 14366 4088 14372 4140
rect 14424 4088 14430 4140
rect 14458 4088 14464 4140
rect 14516 4128 14522 4140
rect 18322 4128 18328 4140
rect 14516 4100 18328 4128
rect 14516 4088 14522 4100
rect 18322 4088 18328 4100
rect 18380 4088 18386 4140
rect 4203 4032 5120 4060
rect 4203 4029 4215 4032
rect 4157 4023 4215 4029
rect 4172 3924 4200 4023
rect 10502 4020 10508 4072
rect 10560 4060 10566 4072
rect 14093 4063 14151 4069
rect 10560 4032 13952 4060
rect 10560 4020 10566 4032
rect 9490 3992 9496 4004
rect 9451 3964 9496 3992
rect 9490 3952 9496 3964
rect 9548 3952 9554 4004
rect 3528 3896 4200 3924
rect 4246 3884 4252 3936
rect 4304 3924 4310 3936
rect 4801 3927 4859 3933
rect 4801 3924 4813 3927
rect 4304 3896 4813 3924
rect 4304 3884 4310 3896
rect 4801 3893 4813 3896
rect 4847 3924 4859 3927
rect 7466 3924 7472 3936
rect 4847 3896 7472 3924
rect 4847 3893 4859 3896
rect 4801 3887 4859 3893
rect 7466 3884 7472 3896
rect 7524 3884 7530 3936
rect 10778 3884 10784 3936
rect 10836 3924 10842 3936
rect 13817 3927 13875 3933
rect 13817 3924 13829 3927
rect 10836 3896 13829 3924
rect 10836 3884 10842 3896
rect 13817 3893 13829 3896
rect 13863 3893 13875 3927
rect 13924 3924 13952 4032
rect 14093 4029 14105 4063
rect 14139 4060 14151 4063
rect 15562 4060 15568 4072
rect 14139 4032 15568 4060
rect 14139 4029 14151 4032
rect 14093 4023 14151 4029
rect 15562 4020 15568 4032
rect 15620 4020 15626 4072
rect 17494 4060 17500 4072
rect 16546 4032 17500 4060
rect 14182 3992 14188 4004
rect 14143 3964 14188 3992
rect 14182 3952 14188 3964
rect 14240 3952 14246 4004
rect 16546 3992 16574 4032
rect 17494 4020 17500 4032
rect 17552 4060 17558 4072
rect 18049 4063 18107 4069
rect 18049 4060 18061 4063
rect 17552 4032 18061 4060
rect 17552 4020 17558 4032
rect 18049 4029 18061 4032
rect 18095 4029 18107 4063
rect 18049 4023 18107 4029
rect 14292 3964 16574 3992
rect 19061 3995 19119 4001
rect 14292 3924 14320 3964
rect 19061 3961 19073 3995
rect 19107 3992 19119 3995
rect 19628 3992 19656 4159
rect 23750 4156 23756 4168
rect 23808 4156 23814 4208
rect 27614 4196 27620 4208
rect 27575 4168 27620 4196
rect 27614 4156 27620 4168
rect 27672 4156 27678 4208
rect 20254 4128 20260 4140
rect 20215 4100 20260 4128
rect 20254 4088 20260 4100
rect 20312 4088 20318 4140
rect 20438 4128 20444 4140
rect 20399 4100 20444 4128
rect 20438 4088 20444 4100
rect 20496 4088 20502 4140
rect 23474 4128 23480 4140
rect 23435 4100 23480 4128
rect 23474 4088 23480 4100
rect 23532 4088 23538 4140
rect 27982 4088 27988 4140
rect 28040 4128 28046 4140
rect 28077 4131 28135 4137
rect 28077 4128 28089 4131
rect 28040 4100 28089 4128
rect 28040 4088 28046 4100
rect 28077 4097 28089 4100
rect 28123 4097 28135 4131
rect 28077 4091 28135 4097
rect 28353 4131 28411 4137
rect 28353 4097 28365 4131
rect 28399 4128 28411 4131
rect 30834 4128 30840 4140
rect 28399 4100 30840 4128
rect 28399 4097 28411 4100
rect 28353 4091 28411 4097
rect 30834 4088 30840 4100
rect 30892 4088 30898 4140
rect 19107 3964 19656 3992
rect 19107 3961 19119 3964
rect 19061 3955 19119 3961
rect 13924 3896 14320 3924
rect 13817 3887 13875 3893
rect 14366 3884 14372 3936
rect 14424 3924 14430 3936
rect 14918 3924 14924 3936
rect 14424 3896 14924 3924
rect 14424 3884 14430 3896
rect 14918 3884 14924 3896
rect 14976 3884 14982 3936
rect 19702 3924 19708 3936
rect 19663 3896 19708 3924
rect 19702 3884 19708 3896
rect 19760 3884 19766 3936
rect 20254 3924 20260 3936
rect 20215 3896 20260 3924
rect 20254 3884 20260 3896
rect 20312 3884 20318 3936
rect 23661 3927 23719 3933
rect 23661 3893 23673 3927
rect 23707 3924 23719 3927
rect 24302 3924 24308 3936
rect 23707 3896 24308 3924
rect 23707 3893 23719 3896
rect 23661 3887 23719 3893
rect 24302 3884 24308 3896
rect 24360 3884 24366 3936
rect 27433 3927 27491 3933
rect 27433 3893 27445 3927
rect 27479 3924 27491 3927
rect 28534 3924 28540 3936
rect 27479 3896 28540 3924
rect 27479 3893 27491 3896
rect 27433 3887 27491 3893
rect 28534 3884 28540 3896
rect 28592 3884 28598 3936
rect 1104 3834 38824 3856
rect 1104 3782 5674 3834
rect 5726 3782 5738 3834
rect 5790 3782 5802 3834
rect 5854 3782 5866 3834
rect 5918 3782 5930 3834
rect 5982 3782 15122 3834
rect 15174 3782 15186 3834
rect 15238 3782 15250 3834
rect 15302 3782 15314 3834
rect 15366 3782 15378 3834
rect 15430 3782 24570 3834
rect 24622 3782 24634 3834
rect 24686 3782 24698 3834
rect 24750 3782 24762 3834
rect 24814 3782 24826 3834
rect 24878 3782 34018 3834
rect 34070 3782 34082 3834
rect 34134 3782 34146 3834
rect 34198 3782 34210 3834
rect 34262 3782 34274 3834
rect 34326 3782 38824 3834
rect 1104 3760 38824 3782
rect 11517 3723 11575 3729
rect 11517 3689 11529 3723
rect 11563 3720 11575 3723
rect 12066 3720 12072 3732
rect 11563 3692 12072 3720
rect 11563 3689 11575 3692
rect 11517 3683 11575 3689
rect 12066 3680 12072 3692
rect 12124 3680 12130 3732
rect 14182 3680 14188 3732
rect 14240 3720 14246 3732
rect 15105 3723 15163 3729
rect 15105 3720 15117 3723
rect 14240 3692 15117 3720
rect 14240 3680 14246 3692
rect 15105 3689 15117 3692
rect 15151 3689 15163 3723
rect 16758 3720 16764 3732
rect 16719 3692 16764 3720
rect 15105 3683 15163 3689
rect 16758 3680 16764 3692
rect 16816 3680 16822 3732
rect 20714 3680 20720 3732
rect 20772 3720 20778 3732
rect 21361 3723 21419 3729
rect 21361 3720 21373 3723
rect 20772 3692 21373 3720
rect 20772 3680 20778 3692
rect 21361 3689 21373 3692
rect 21407 3689 21419 3723
rect 21361 3683 21419 3689
rect 31754 3680 31760 3732
rect 31812 3720 31818 3732
rect 32401 3723 32459 3729
rect 32401 3720 32413 3723
rect 31812 3692 32413 3720
rect 31812 3680 31818 3692
rect 32401 3689 32413 3692
rect 32447 3689 32459 3723
rect 36814 3720 36820 3732
rect 36775 3692 36820 3720
rect 32401 3683 32459 3689
rect 36814 3680 36820 3692
rect 36872 3680 36878 3732
rect 11974 3652 11980 3664
rect 11935 3624 11980 3652
rect 11974 3612 11980 3624
rect 12032 3612 12038 3664
rect 12989 3655 13047 3661
rect 12989 3652 13001 3655
rect 12176 3624 13001 3652
rect 10502 3584 10508 3596
rect 10463 3556 10508 3584
rect 10502 3544 10508 3556
rect 10560 3544 10566 3596
rect 1673 3519 1731 3525
rect 1673 3485 1685 3519
rect 1719 3516 1731 3519
rect 2866 3516 2872 3528
rect 1719 3488 2728 3516
rect 2827 3488 2872 3516
rect 1719 3485 1731 3488
rect 1673 3479 1731 3485
rect 1486 3380 1492 3392
rect 1447 3352 1492 3380
rect 1486 3340 1492 3352
rect 1544 3340 1550 3392
rect 2700 3389 2728 3488
rect 2866 3476 2872 3488
rect 2924 3476 2930 3528
rect 10778 3516 10784 3528
rect 10739 3488 10784 3516
rect 10778 3476 10784 3488
rect 10836 3476 10842 3528
rect 12176 3525 12204 3624
rect 12989 3621 13001 3624
rect 13035 3652 13047 3655
rect 14366 3652 14372 3664
rect 13035 3624 14372 3652
rect 13035 3621 13047 3624
rect 12989 3615 13047 3621
rect 14366 3612 14372 3624
rect 14424 3612 14430 3664
rect 21177 3655 21235 3661
rect 21177 3652 21189 3655
rect 16408 3624 21189 3652
rect 14458 3584 14464 3596
rect 12544 3556 14464 3584
rect 12161 3519 12219 3525
rect 12161 3485 12173 3519
rect 12207 3485 12219 3519
rect 12434 3516 12440 3528
rect 12395 3488 12440 3516
rect 12161 3479 12219 3485
rect 12434 3476 12440 3488
rect 12492 3476 12498 3528
rect 12345 3451 12403 3457
rect 12345 3417 12357 3451
rect 12391 3448 12403 3451
rect 12544 3448 12572 3556
rect 14458 3544 14464 3556
rect 14516 3544 14522 3596
rect 14642 3544 14648 3596
rect 14700 3584 14706 3596
rect 16408 3584 16436 3624
rect 21177 3621 21189 3624
rect 21223 3621 21235 3655
rect 21177 3615 21235 3621
rect 31294 3612 31300 3664
rect 31352 3652 31358 3664
rect 31389 3655 31447 3661
rect 31389 3652 31401 3655
rect 31352 3624 31401 3652
rect 31352 3612 31358 3624
rect 31389 3621 31401 3624
rect 31435 3652 31447 3655
rect 32217 3655 32275 3661
rect 32217 3652 32229 3655
rect 31435 3624 32229 3652
rect 31435 3621 31447 3624
rect 31389 3615 31447 3621
rect 32217 3621 32229 3624
rect 32263 3621 32275 3655
rect 36633 3655 36691 3661
rect 36633 3652 36645 3655
rect 32217 3615 32275 3621
rect 32508 3624 36645 3652
rect 20254 3584 20260 3596
rect 14700 3556 16436 3584
rect 16500 3556 20260 3584
rect 14700 3544 14706 3556
rect 14366 3516 14372 3528
rect 14327 3488 14372 3516
rect 14366 3476 14372 3488
rect 14424 3476 14430 3528
rect 14553 3519 14611 3525
rect 14553 3485 14565 3519
rect 14599 3485 14611 3519
rect 14553 3479 14611 3485
rect 14737 3519 14795 3525
rect 14737 3485 14749 3519
rect 14783 3485 14795 3519
rect 14737 3479 14795 3485
rect 14829 3519 14887 3525
rect 14829 3485 14841 3519
rect 14875 3516 14887 3519
rect 16500 3516 16528 3556
rect 20254 3544 20260 3556
rect 20312 3544 20318 3596
rect 21545 3587 21603 3593
rect 21545 3553 21557 3587
rect 21591 3584 21603 3587
rect 22922 3584 22928 3596
rect 21591 3556 22928 3584
rect 21591 3553 21603 3556
rect 21545 3547 21603 3553
rect 22922 3544 22928 3556
rect 22980 3544 22986 3596
rect 24394 3544 24400 3596
rect 24452 3584 24458 3596
rect 26878 3584 26884 3596
rect 24452 3556 26884 3584
rect 24452 3544 24458 3556
rect 26878 3544 26884 3556
rect 26936 3544 26942 3596
rect 30193 3587 30251 3593
rect 30193 3553 30205 3587
rect 30239 3584 30251 3587
rect 31481 3587 31539 3593
rect 31481 3584 31493 3587
rect 30239 3556 31493 3584
rect 30239 3553 30251 3556
rect 30193 3547 30251 3553
rect 31404 3528 31432 3556
rect 31481 3553 31493 3556
rect 31527 3553 31539 3587
rect 31481 3547 31539 3553
rect 31570 3544 31576 3596
rect 31628 3584 31634 3596
rect 32508 3584 32536 3624
rect 36633 3621 36645 3624
rect 36679 3621 36691 3655
rect 36633 3615 36691 3621
rect 31628 3556 32536 3584
rect 32585 3587 32643 3593
rect 31628 3544 31634 3556
rect 32585 3553 32597 3587
rect 32631 3584 32643 3587
rect 33686 3584 33692 3596
rect 32631 3556 33692 3584
rect 32631 3553 32643 3556
rect 32585 3547 32643 3553
rect 33686 3544 33692 3556
rect 33744 3544 33750 3596
rect 14875 3488 16528 3516
rect 16577 3519 16635 3525
rect 14875 3485 14887 3488
rect 14829 3479 14887 3485
rect 16577 3485 16589 3519
rect 16623 3485 16635 3519
rect 16577 3479 16635 3485
rect 16669 3519 16727 3525
rect 16669 3485 16681 3519
rect 16715 3516 16727 3519
rect 19242 3516 19248 3528
rect 16715 3488 19248 3516
rect 16715 3485 16727 3488
rect 16669 3479 16727 3485
rect 12391 3420 12572 3448
rect 12391 3417 12403 3420
rect 12345 3411 12403 3417
rect 14182 3408 14188 3460
rect 14240 3448 14246 3460
rect 14568 3448 14596 3479
rect 14240 3420 14596 3448
rect 14240 3408 14246 3420
rect 2685 3383 2743 3389
rect 2685 3349 2697 3383
rect 2731 3349 2743 3383
rect 2685 3343 2743 3349
rect 14550 3340 14556 3392
rect 14608 3380 14614 3392
rect 14752 3380 14780 3479
rect 16393 3383 16451 3389
rect 16393 3380 16405 3383
rect 14608 3352 16405 3380
rect 14608 3340 14614 3352
rect 16393 3349 16405 3352
rect 16439 3349 16451 3383
rect 16592 3380 16620 3479
rect 19242 3476 19248 3488
rect 19300 3476 19306 3528
rect 21358 3516 21364 3528
rect 21319 3488 21364 3516
rect 21358 3476 21364 3488
rect 21416 3476 21422 3528
rect 27157 3519 27215 3525
rect 27157 3485 27169 3519
rect 27203 3516 27215 3519
rect 27338 3516 27344 3528
rect 27203 3488 27344 3516
rect 27203 3485 27215 3488
rect 27157 3479 27215 3485
rect 27338 3476 27344 3488
rect 27396 3476 27402 3528
rect 27982 3516 27988 3528
rect 27943 3488 27988 3516
rect 27982 3476 27988 3488
rect 28040 3516 28046 3528
rect 28445 3519 28503 3525
rect 28445 3516 28457 3519
rect 28040 3488 28457 3516
rect 28040 3476 28046 3488
rect 28445 3485 28457 3488
rect 28491 3485 28503 3519
rect 28445 3479 28503 3485
rect 28534 3476 28540 3528
rect 28592 3516 28598 3528
rect 31297 3519 31355 3525
rect 31297 3516 31309 3519
rect 28592 3488 31309 3516
rect 28592 3476 28598 3488
rect 31297 3485 31309 3488
rect 31343 3485 31355 3519
rect 31297 3479 31355 3485
rect 31386 3476 31392 3528
rect 31444 3476 31450 3528
rect 31757 3519 31815 3525
rect 31757 3485 31769 3519
rect 31803 3516 31815 3519
rect 31846 3516 31852 3528
rect 31803 3488 31852 3516
rect 31803 3485 31815 3488
rect 31757 3479 31815 3485
rect 31846 3476 31852 3488
rect 31904 3476 31910 3528
rect 32398 3516 32404 3528
rect 32359 3488 32404 3516
rect 32398 3476 32404 3488
rect 32456 3476 32462 3528
rect 36817 3519 36875 3525
rect 36817 3485 36829 3519
rect 36863 3485 36875 3519
rect 36817 3479 36875 3485
rect 36909 3519 36967 3525
rect 36909 3485 36921 3519
rect 36955 3516 36967 3519
rect 37918 3516 37924 3528
rect 36955 3488 37924 3516
rect 36955 3485 36967 3488
rect 36909 3479 36967 3485
rect 16850 3448 16856 3460
rect 16811 3420 16856 3448
rect 16850 3408 16856 3420
rect 16908 3408 16914 3460
rect 21637 3451 21695 3457
rect 21637 3417 21649 3451
rect 21683 3448 21695 3451
rect 22462 3448 22468 3460
rect 21683 3420 22468 3448
rect 21683 3417 21695 3420
rect 21637 3411 21695 3417
rect 22462 3408 22468 3420
rect 22520 3408 22526 3460
rect 28994 3408 29000 3460
rect 29052 3448 29058 3460
rect 29825 3451 29883 3457
rect 29825 3448 29837 3451
rect 29052 3420 29837 3448
rect 29052 3408 29058 3420
rect 29825 3417 29837 3420
rect 29871 3417 29883 3451
rect 30006 3448 30012 3460
rect 29967 3420 30012 3448
rect 29825 3411 29883 3417
rect 30006 3408 30012 3420
rect 30064 3408 30070 3460
rect 32677 3451 32735 3457
rect 32677 3417 32689 3451
rect 32723 3448 32735 3451
rect 33226 3448 33232 3460
rect 32723 3420 33232 3448
rect 32723 3417 32735 3420
rect 32677 3411 32735 3417
rect 33226 3408 33232 3420
rect 33284 3408 33290 3460
rect 16666 3380 16672 3392
rect 16592 3352 16672 3380
rect 16393 3343 16451 3349
rect 16666 3340 16672 3352
rect 16724 3340 16730 3392
rect 23474 3380 23480 3392
rect 23435 3352 23480 3380
rect 23474 3340 23480 3352
rect 23532 3340 23538 3392
rect 31018 3380 31024 3392
rect 30979 3352 31024 3380
rect 31018 3340 31024 3352
rect 31076 3340 31082 3392
rect 36832 3380 36860 3479
rect 37918 3476 37924 3488
rect 37976 3476 37982 3528
rect 37093 3451 37151 3457
rect 37093 3417 37105 3451
rect 37139 3448 37151 3451
rect 37642 3448 37648 3460
rect 37139 3420 37648 3448
rect 37139 3417 37151 3420
rect 37093 3411 37151 3417
rect 37642 3408 37648 3420
rect 37700 3408 37706 3460
rect 37274 3380 37280 3392
rect 36832 3352 37280 3380
rect 37274 3340 37280 3352
rect 37332 3340 37338 3392
rect 38102 3380 38108 3392
rect 38063 3352 38108 3380
rect 38102 3340 38108 3352
rect 38160 3340 38166 3392
rect 1104 3290 38824 3312
rect 1104 3238 10398 3290
rect 10450 3238 10462 3290
rect 10514 3238 10526 3290
rect 10578 3238 10590 3290
rect 10642 3238 10654 3290
rect 10706 3238 19846 3290
rect 19898 3238 19910 3290
rect 19962 3238 19974 3290
rect 20026 3238 20038 3290
rect 20090 3238 20102 3290
rect 20154 3238 29294 3290
rect 29346 3238 29358 3290
rect 29410 3238 29422 3290
rect 29474 3238 29486 3290
rect 29538 3238 29550 3290
rect 29602 3238 38824 3290
rect 1104 3216 38824 3238
rect 2130 3176 2136 3188
rect 2091 3148 2136 3176
rect 2130 3136 2136 3148
rect 2188 3136 2194 3188
rect 4985 3179 5043 3185
rect 4985 3145 4997 3179
rect 5031 3176 5043 3179
rect 5534 3176 5540 3188
rect 5031 3148 5540 3176
rect 5031 3145 5043 3148
rect 4985 3139 5043 3145
rect 5534 3136 5540 3148
rect 5592 3136 5598 3188
rect 12434 3136 12440 3188
rect 12492 3176 12498 3188
rect 14461 3179 14519 3185
rect 14461 3176 14473 3179
rect 12492 3148 14473 3176
rect 12492 3136 12498 3148
rect 14461 3145 14473 3148
rect 14507 3145 14519 3179
rect 37918 3176 37924 3188
rect 37879 3148 37924 3176
rect 14461 3139 14519 3145
rect 37918 3136 37924 3148
rect 37976 3136 37982 3188
rect 14185 3111 14243 3117
rect 14185 3077 14197 3111
rect 14231 3108 14243 3111
rect 14366 3108 14372 3120
rect 14231 3080 14372 3108
rect 14231 3077 14243 3080
rect 14185 3071 14243 3077
rect 14366 3068 14372 3080
rect 14424 3068 14430 3120
rect 14550 3108 14556 3120
rect 14511 3080 14556 3108
rect 14550 3068 14556 3080
rect 14608 3068 14614 3120
rect 14918 3068 14924 3120
rect 14976 3108 14982 3120
rect 31018 3108 31024 3120
rect 14976 3080 31024 3108
rect 14976 3068 14982 3080
rect 31018 3068 31024 3080
rect 31076 3068 31082 3120
rect 31570 3108 31576 3120
rect 31531 3080 31576 3108
rect 31570 3068 31576 3080
rect 31628 3068 31634 3120
rect 2869 3043 2927 3049
rect 2869 3009 2881 3043
rect 2915 3040 2927 3043
rect 23477 3043 23535 3049
rect 2915 3012 3464 3040
rect 2915 3009 2927 3012
rect 2869 3003 2927 3009
rect 3436 2913 3464 3012
rect 23477 3009 23489 3043
rect 23523 3040 23535 3043
rect 23566 3040 23572 3052
rect 23523 3012 23572 3040
rect 23523 3009 23535 3012
rect 23477 3003 23535 3009
rect 23566 3000 23572 3012
rect 23624 3000 23630 3052
rect 24302 3040 24308 3052
rect 24263 3012 24308 3040
rect 24302 3000 24308 3012
rect 24360 3000 24366 3052
rect 24394 3000 24400 3052
rect 24452 3040 24458 3052
rect 24581 3043 24639 3049
rect 24581 3040 24593 3043
rect 24452 3012 24593 3040
rect 24452 3000 24458 3012
rect 24581 3009 24593 3012
rect 24627 3009 24639 3043
rect 31294 3040 31300 3052
rect 31255 3012 31300 3040
rect 24581 3003 24639 3009
rect 31294 3000 31300 3012
rect 31352 3000 31358 3052
rect 31386 3000 31392 3052
rect 31444 3040 31450 3052
rect 38102 3040 38108 3052
rect 31444 3012 31489 3040
rect 38015 3012 38108 3040
rect 31444 3000 31450 3012
rect 38102 3000 38108 3012
rect 38160 3040 38166 3052
rect 39114 3040 39120 3052
rect 38160 3012 39120 3040
rect 38160 3000 38166 3012
rect 39114 3000 39120 3012
rect 39172 3000 39178 3052
rect 14369 2975 14427 2981
rect 14369 2941 14381 2975
rect 14415 2972 14427 2975
rect 14642 2972 14648 2984
rect 14415 2944 14648 2972
rect 14415 2941 14427 2944
rect 14369 2935 14427 2941
rect 14642 2932 14648 2944
rect 14700 2932 14706 2984
rect 17586 2972 17592 2984
rect 16546 2944 17592 2972
rect 3421 2907 3479 2913
rect 3421 2873 3433 2907
rect 3467 2904 3479 2907
rect 16546 2904 16574 2944
rect 17586 2932 17592 2944
rect 17644 2932 17650 2984
rect 36725 2975 36783 2981
rect 36725 2941 36737 2975
rect 36771 2972 36783 2975
rect 38010 2972 38016 2984
rect 36771 2944 38016 2972
rect 36771 2941 36783 2944
rect 36725 2935 36783 2941
rect 38010 2932 38016 2944
rect 38068 2932 38074 2984
rect 3467 2876 16574 2904
rect 3467 2873 3479 2876
rect 3421 2867 3479 2873
rect 27522 2864 27528 2916
rect 27580 2904 27586 2916
rect 31297 2907 31355 2913
rect 31297 2904 31309 2907
rect 27580 2876 31309 2904
rect 27580 2864 27586 2876
rect 31297 2873 31309 2876
rect 31343 2873 31355 2907
rect 31297 2867 31355 2873
rect 2222 2796 2228 2848
rect 2280 2836 2286 2848
rect 2685 2839 2743 2845
rect 2685 2836 2697 2839
rect 2280 2808 2697 2836
rect 2280 2796 2286 2808
rect 2685 2805 2697 2808
rect 2731 2805 2743 2839
rect 12802 2836 12808 2848
rect 12763 2808 12808 2836
rect 2685 2799 2743 2805
rect 12802 2796 12808 2808
rect 12860 2796 12866 2848
rect 13725 2839 13783 2845
rect 13725 2805 13737 2839
rect 13771 2836 13783 2839
rect 13998 2836 14004 2848
rect 13771 2808 14004 2836
rect 13771 2805 13783 2808
rect 13725 2799 13783 2805
rect 13998 2796 14004 2808
rect 14056 2796 14062 2848
rect 14182 2796 14188 2848
rect 14240 2836 14246 2848
rect 14277 2839 14335 2845
rect 14277 2836 14289 2839
rect 14240 2808 14289 2836
rect 14240 2796 14246 2808
rect 14277 2805 14289 2808
rect 14323 2805 14335 2839
rect 17586 2836 17592 2848
rect 17547 2808 17592 2836
rect 14277 2799 14335 2805
rect 17586 2796 17592 2808
rect 17644 2796 17650 2848
rect 19981 2839 20039 2845
rect 19981 2805 19993 2839
rect 20027 2836 20039 2839
rect 20254 2836 20260 2848
rect 20027 2808 20260 2836
rect 20027 2805 20039 2808
rect 19981 2799 20039 2805
rect 20254 2796 20260 2808
rect 20312 2796 20318 2848
rect 28350 2836 28356 2848
rect 28311 2808 28356 2836
rect 28350 2796 28356 2808
rect 28408 2796 28414 2848
rect 31938 2796 31944 2848
rect 31996 2836 32002 2848
rect 32125 2839 32183 2845
rect 32125 2836 32137 2839
rect 31996 2808 32137 2836
rect 31996 2796 32002 2808
rect 32125 2805 32137 2808
rect 32171 2805 32183 2839
rect 34514 2836 34520 2848
rect 34475 2808 34520 2836
rect 32125 2799 32183 2805
rect 34514 2796 34520 2808
rect 34572 2796 34578 2848
rect 36722 2796 36728 2848
rect 36780 2836 36786 2848
rect 37277 2839 37335 2845
rect 37277 2836 37289 2839
rect 36780 2808 37289 2836
rect 36780 2796 36786 2808
rect 37277 2805 37289 2808
rect 37323 2836 37335 2839
rect 37458 2836 37464 2848
rect 37323 2808 37464 2836
rect 37323 2805 37335 2808
rect 37277 2799 37335 2805
rect 37458 2796 37464 2808
rect 37516 2796 37522 2848
rect 1104 2746 38824 2768
rect 1104 2694 5674 2746
rect 5726 2694 5738 2746
rect 5790 2694 5802 2746
rect 5854 2694 5866 2746
rect 5918 2694 5930 2746
rect 5982 2694 15122 2746
rect 15174 2694 15186 2746
rect 15238 2694 15250 2746
rect 15302 2694 15314 2746
rect 15366 2694 15378 2746
rect 15430 2694 24570 2746
rect 24622 2694 24634 2746
rect 24686 2694 24698 2746
rect 24750 2694 24762 2746
rect 24814 2694 24826 2746
rect 24878 2694 34018 2746
rect 34070 2694 34082 2746
rect 34134 2694 34146 2746
rect 34198 2694 34210 2746
rect 34262 2694 34274 2746
rect 34326 2694 38824 2746
rect 1104 2672 38824 2694
rect 13081 2635 13139 2641
rect 13081 2601 13093 2635
rect 13127 2632 13139 2635
rect 14182 2632 14188 2644
rect 13127 2604 14188 2632
rect 13127 2601 13139 2604
rect 13081 2595 13139 2601
rect 14182 2592 14188 2604
rect 14240 2592 14246 2644
rect 14277 2635 14335 2641
rect 14277 2601 14289 2635
rect 14323 2632 14335 2635
rect 14366 2632 14372 2644
rect 14323 2604 14372 2632
rect 14323 2601 14335 2604
rect 14277 2595 14335 2601
rect 14366 2592 14372 2604
rect 14424 2592 14430 2644
rect 16666 2632 16672 2644
rect 16627 2604 16672 2632
rect 16666 2592 16672 2604
rect 16724 2592 16730 2644
rect 16850 2592 16856 2644
rect 16908 2632 16914 2644
rect 17681 2635 17739 2641
rect 17681 2632 17693 2635
rect 16908 2604 17693 2632
rect 16908 2592 16914 2604
rect 17681 2601 17693 2604
rect 17727 2601 17739 2635
rect 19242 2632 19248 2644
rect 19203 2604 19248 2632
rect 17681 2595 17739 2601
rect 19242 2592 19248 2604
rect 19300 2592 19306 2644
rect 20257 2635 20315 2641
rect 20257 2601 20269 2635
rect 20303 2632 20315 2635
rect 20714 2632 20720 2644
rect 20303 2604 20720 2632
rect 20303 2601 20315 2604
rect 20257 2595 20315 2601
rect 20714 2592 20720 2604
rect 20772 2592 20778 2644
rect 21358 2592 21364 2644
rect 21416 2632 21422 2644
rect 21821 2635 21879 2641
rect 21821 2632 21833 2635
rect 21416 2604 21833 2632
rect 21416 2592 21422 2604
rect 21821 2601 21833 2604
rect 21867 2601 21879 2635
rect 22462 2632 22468 2644
rect 22423 2604 22468 2632
rect 21821 2595 21879 2601
rect 22462 2592 22468 2604
rect 22520 2592 22526 2644
rect 22922 2592 22928 2644
rect 22980 2632 22986 2644
rect 23661 2635 23719 2641
rect 23661 2632 23673 2635
rect 22980 2604 23673 2632
rect 22980 2592 22986 2604
rect 23661 2601 23673 2604
rect 23707 2601 23719 2635
rect 23661 2595 23719 2601
rect 28629 2635 28687 2641
rect 28629 2601 28641 2635
rect 28675 2632 28687 2635
rect 28994 2632 29000 2644
rect 28675 2604 29000 2632
rect 28675 2601 28687 2604
rect 28629 2595 28687 2601
rect 28994 2592 29000 2604
rect 29052 2592 29058 2644
rect 29825 2635 29883 2641
rect 29825 2601 29837 2635
rect 29871 2632 29883 2635
rect 30006 2632 30012 2644
rect 29871 2604 30012 2632
rect 29871 2601 29883 2604
rect 29825 2595 29883 2601
rect 30006 2592 30012 2604
rect 30064 2592 30070 2644
rect 31021 2635 31079 2641
rect 31021 2601 31033 2635
rect 31067 2632 31079 2635
rect 31754 2632 31760 2644
rect 31067 2604 31760 2632
rect 31067 2601 31079 2604
rect 31021 2595 31079 2601
rect 31754 2592 31760 2604
rect 31812 2592 31818 2644
rect 32309 2635 32367 2641
rect 32309 2601 32321 2635
rect 32355 2632 32367 2635
rect 32398 2632 32404 2644
rect 32355 2604 32404 2632
rect 32355 2601 32367 2604
rect 32309 2595 32367 2601
rect 32398 2592 32404 2604
rect 32456 2592 32462 2644
rect 33226 2632 33232 2644
rect 33187 2604 33232 2632
rect 33226 2592 33232 2604
rect 33284 2592 33290 2644
rect 33686 2592 33692 2644
rect 33744 2632 33750 2644
rect 34701 2635 34759 2641
rect 34701 2632 34713 2635
rect 33744 2604 34713 2632
rect 33744 2592 33750 2604
rect 34701 2601 34713 2604
rect 34747 2601 34759 2635
rect 34701 2595 34759 2601
rect 35805 2635 35863 2641
rect 35805 2601 35817 2635
rect 35851 2632 35863 2635
rect 36814 2632 36820 2644
rect 35851 2604 36820 2632
rect 35851 2601 35863 2604
rect 35805 2595 35863 2601
rect 36814 2592 36820 2604
rect 36872 2592 36878 2644
rect 37274 2632 37280 2644
rect 37235 2604 37280 2632
rect 37274 2592 37280 2604
rect 37332 2592 37338 2644
rect 37642 2592 37648 2644
rect 37700 2632 37706 2644
rect 37921 2635 37979 2641
rect 37921 2632 37933 2635
rect 37700 2604 37933 2632
rect 37700 2592 37706 2604
rect 37921 2601 37933 2604
rect 37967 2601 37979 2635
rect 37921 2595 37979 2601
rect 3973 2567 4031 2573
rect 3973 2533 3985 2567
rect 4019 2564 4031 2567
rect 14826 2564 14832 2576
rect 4019 2536 14832 2564
rect 4019 2533 4031 2536
rect 3973 2527 4031 2533
rect 14826 2524 14832 2536
rect 14884 2524 14890 2576
rect 15473 2567 15531 2573
rect 15473 2533 15485 2567
rect 15519 2564 15531 2567
rect 16758 2564 16764 2576
rect 15519 2536 16764 2564
rect 15519 2533 15531 2536
rect 15473 2527 15531 2533
rect 16758 2524 16764 2536
rect 16816 2524 16822 2576
rect 2130 2456 2136 2508
rect 2188 2496 2194 2508
rect 2188 2468 2452 2496
rect 2188 2456 2194 2468
rect 1673 2431 1731 2437
rect 1673 2397 1685 2431
rect 1719 2428 1731 2431
rect 2222 2428 2228 2440
rect 1719 2400 2228 2428
rect 1719 2397 1731 2400
rect 1673 2391 1731 2397
rect 2222 2388 2228 2400
rect 2280 2388 2286 2440
rect 2424 2437 2452 2468
rect 4430 2456 4436 2508
rect 4488 2496 4494 2508
rect 27982 2496 27988 2508
rect 4488 2468 25176 2496
rect 4488 2456 4494 2468
rect 2409 2431 2467 2437
rect 2409 2397 2421 2431
rect 2455 2397 2467 2431
rect 3789 2431 3847 2437
rect 3789 2428 3801 2431
rect 2409 2391 2467 2397
rect 3252 2400 3801 2428
rect 3252 2304 3280 2400
rect 3789 2397 3801 2400
rect 3835 2397 3847 2431
rect 3789 2391 3847 2397
rect 4801 2431 4859 2437
rect 4801 2397 4813 2431
rect 4847 2428 4859 2431
rect 5534 2428 5540 2440
rect 4847 2400 5540 2428
rect 4847 2397 4859 2400
rect 4801 2391 4859 2397
rect 5534 2388 5540 2400
rect 5592 2388 5598 2440
rect 5813 2431 5871 2437
rect 5813 2397 5825 2431
rect 5859 2428 5871 2431
rect 6270 2428 6276 2440
rect 5859 2400 6276 2428
rect 5859 2397 5871 2400
rect 5813 2391 5871 2397
rect 6270 2388 6276 2400
rect 6328 2388 6334 2440
rect 7190 2428 7196 2440
rect 7151 2400 7196 2428
rect 7190 2388 7196 2400
rect 7248 2388 7254 2440
rect 8386 2428 8392 2440
rect 8347 2400 8392 2428
rect 8386 2388 8392 2400
rect 8444 2388 8450 2440
rect 9585 2431 9643 2437
rect 9585 2397 9597 2431
rect 9631 2428 9643 2431
rect 11977 2431 12035 2437
rect 9631 2400 10180 2428
rect 9631 2397 9643 2400
rect 9585 2391 9643 2397
rect 10152 2369 10180 2400
rect 11977 2397 11989 2431
rect 12023 2428 12035 2431
rect 12434 2428 12440 2440
rect 12023 2400 12440 2428
rect 12023 2397 12035 2400
rect 11977 2391 12035 2397
rect 12434 2388 12440 2400
rect 12492 2388 12498 2440
rect 12802 2388 12808 2440
rect 12860 2428 12866 2440
rect 12897 2431 12955 2437
rect 12897 2428 12909 2431
rect 12860 2400 12909 2428
rect 12860 2388 12866 2400
rect 12897 2397 12909 2400
rect 12943 2397 12955 2431
rect 12897 2391 12955 2397
rect 13998 2388 14004 2440
rect 14056 2428 14062 2440
rect 14093 2431 14151 2437
rect 14093 2428 14105 2431
rect 14056 2400 14105 2428
rect 14056 2388 14062 2400
rect 14093 2397 14105 2400
rect 14139 2397 14151 2431
rect 14093 2391 14151 2397
rect 14829 2431 14887 2437
rect 14829 2397 14841 2431
rect 14875 2428 14887 2431
rect 15194 2428 15200 2440
rect 14875 2400 15200 2428
rect 14875 2397 14887 2400
rect 14829 2391 14887 2397
rect 15194 2388 15200 2400
rect 15252 2428 15258 2440
rect 15289 2431 15347 2437
rect 15289 2428 15301 2431
rect 15252 2400 15301 2428
rect 15252 2388 15258 2400
rect 15289 2397 15301 2400
rect 15335 2397 15347 2431
rect 15289 2391 15347 2397
rect 16117 2431 16175 2437
rect 16117 2397 16129 2431
rect 16163 2428 16175 2431
rect 16390 2428 16396 2440
rect 16163 2400 16396 2428
rect 16163 2397 16175 2400
rect 16117 2391 16175 2397
rect 16390 2388 16396 2400
rect 16448 2428 16454 2440
rect 16853 2431 16911 2437
rect 16853 2428 16865 2431
rect 16448 2400 16865 2428
rect 16448 2388 16454 2400
rect 16853 2397 16865 2400
rect 16899 2397 16911 2431
rect 16853 2391 16911 2397
rect 17586 2388 17592 2440
rect 17644 2428 17650 2440
rect 17865 2431 17923 2437
rect 17865 2428 17877 2431
rect 17644 2400 17877 2428
rect 17644 2388 17650 2400
rect 17865 2397 17877 2400
rect 17911 2397 17923 2431
rect 17865 2391 17923 2397
rect 18782 2388 18788 2440
rect 18840 2428 18846 2440
rect 19429 2431 19487 2437
rect 19429 2428 19441 2431
rect 18840 2400 19441 2428
rect 18840 2388 18846 2400
rect 19429 2397 19441 2400
rect 19475 2397 19487 2431
rect 19429 2391 19487 2397
rect 20073 2431 20131 2437
rect 20073 2397 20085 2431
rect 20119 2428 20131 2431
rect 20254 2428 20260 2440
rect 20119 2400 20260 2428
rect 20119 2397 20131 2400
rect 20073 2391 20131 2397
rect 20254 2388 20260 2400
rect 20312 2388 20318 2440
rect 22005 2431 22063 2437
rect 22005 2428 22017 2431
rect 21192 2400 22017 2428
rect 10137 2363 10195 2369
rect 10137 2329 10149 2363
rect 10183 2360 10195 2363
rect 19702 2360 19708 2372
rect 10183 2332 19708 2360
rect 10183 2329 10195 2332
rect 10137 2323 10195 2329
rect 19702 2320 19708 2332
rect 19760 2320 19766 2372
rect 21192 2304 21220 2400
rect 22005 2397 22017 2400
rect 22051 2397 22063 2431
rect 22005 2391 22063 2397
rect 22370 2388 22376 2440
rect 22428 2428 22434 2440
rect 22649 2431 22707 2437
rect 22649 2428 22661 2431
rect 22428 2400 22661 2428
rect 22428 2388 22434 2400
rect 22649 2397 22661 2400
rect 22695 2428 22707 2431
rect 23109 2431 23167 2437
rect 23109 2428 23121 2431
rect 22695 2400 23121 2428
rect 22695 2397 22707 2400
rect 22649 2391 22707 2397
rect 23109 2397 23121 2400
rect 23155 2397 23167 2431
rect 23109 2391 23167 2397
rect 23566 2388 23572 2440
rect 23624 2428 23630 2440
rect 25148 2437 25176 2468
rect 26206 2468 27988 2496
rect 23845 2431 23903 2437
rect 23845 2428 23857 2431
rect 23624 2400 23857 2428
rect 23624 2388 23630 2400
rect 23845 2397 23857 2400
rect 23891 2397 23903 2431
rect 23845 2391 23903 2397
rect 25133 2431 25191 2437
rect 25133 2397 25145 2431
rect 25179 2428 25191 2431
rect 25593 2431 25651 2437
rect 25593 2428 25605 2431
rect 25179 2400 25605 2428
rect 25179 2397 25191 2400
rect 25133 2391 25191 2397
rect 25593 2397 25605 2400
rect 25639 2428 25651 2431
rect 26206 2428 26234 2468
rect 27982 2456 27988 2468
rect 28040 2456 28046 2508
rect 27522 2428 27528 2440
rect 25639 2400 26234 2428
rect 27483 2400 27528 2428
rect 25639 2397 25651 2400
rect 25593 2391 25651 2397
rect 27522 2388 27528 2400
rect 27580 2388 27586 2440
rect 28350 2388 28356 2440
rect 28408 2428 28414 2440
rect 28445 2431 28503 2437
rect 28445 2428 28457 2431
rect 28408 2400 28457 2428
rect 28408 2388 28414 2400
rect 28445 2397 28457 2400
rect 28491 2397 28503 2431
rect 29638 2428 29644 2440
rect 29599 2400 29644 2428
rect 28445 2391 28503 2397
rect 29638 2388 29644 2400
rect 29696 2428 29702 2440
rect 30285 2431 30343 2437
rect 30285 2428 30297 2431
rect 29696 2400 30297 2428
rect 29696 2388 29702 2400
rect 30285 2397 30297 2400
rect 30331 2397 30343 2431
rect 30285 2391 30343 2397
rect 30742 2388 30748 2440
rect 30800 2428 30806 2440
rect 30837 2431 30895 2437
rect 30837 2428 30849 2431
rect 30800 2400 30849 2428
rect 30800 2388 30806 2400
rect 30837 2397 30849 2400
rect 30883 2428 30895 2431
rect 31481 2431 31539 2437
rect 31481 2428 31493 2431
rect 30883 2400 31493 2428
rect 30883 2397 30895 2400
rect 30837 2391 30895 2397
rect 31481 2397 31493 2400
rect 31527 2397 31539 2431
rect 31481 2391 31539 2397
rect 31938 2388 31944 2440
rect 31996 2428 32002 2440
rect 32125 2431 32183 2437
rect 32125 2428 32137 2431
rect 31996 2400 32137 2428
rect 31996 2388 32002 2400
rect 32125 2397 32137 2400
rect 32171 2397 32183 2431
rect 32125 2391 32183 2397
rect 33134 2388 33140 2440
rect 33192 2428 33198 2440
rect 33413 2431 33471 2437
rect 33413 2428 33425 2431
rect 33192 2400 33425 2428
rect 33192 2388 33198 2400
rect 33413 2397 33425 2400
rect 33459 2428 33471 2431
rect 33873 2431 33931 2437
rect 33873 2428 33885 2431
rect 33459 2400 33885 2428
rect 33459 2397 33471 2400
rect 33413 2391 33471 2397
rect 33873 2397 33885 2400
rect 33919 2397 33931 2431
rect 33873 2391 33931 2397
rect 34514 2388 34520 2440
rect 34572 2428 34578 2440
rect 34885 2431 34943 2437
rect 34885 2428 34897 2431
rect 34572 2400 34897 2428
rect 34572 2388 34578 2400
rect 34885 2397 34897 2400
rect 34931 2397 34943 2431
rect 34885 2391 34943 2397
rect 35526 2388 35532 2440
rect 35584 2428 35590 2440
rect 35621 2431 35679 2437
rect 35621 2428 35633 2431
rect 35584 2400 35633 2428
rect 35584 2388 35590 2400
rect 35621 2397 35633 2400
rect 35667 2428 35679 2431
rect 36265 2431 36323 2437
rect 36265 2428 36277 2431
rect 35667 2400 36277 2428
rect 35667 2397 35679 2400
rect 35621 2391 35679 2397
rect 36265 2397 36277 2400
rect 36311 2397 36323 2431
rect 37458 2428 37464 2440
rect 37419 2400 37464 2428
rect 36265 2391 36323 2397
rect 37458 2388 37464 2400
rect 37516 2388 37522 2440
rect 38010 2388 38016 2440
rect 38068 2428 38074 2440
rect 38105 2431 38163 2437
rect 38105 2428 38117 2431
rect 38068 2400 38117 2428
rect 38068 2388 38074 2400
rect 38105 2397 38117 2400
rect 38151 2397 38163 2431
rect 38105 2391 38163 2397
rect 1486 2292 1492 2304
rect 1447 2264 1492 2292
rect 1486 2252 1492 2264
rect 1544 2252 1550 2304
rect 2038 2252 2044 2304
rect 2096 2292 2102 2304
rect 2225 2295 2283 2301
rect 2225 2292 2237 2295
rect 2096 2264 2237 2292
rect 2096 2252 2102 2264
rect 2225 2261 2237 2264
rect 2271 2261 2283 2295
rect 3234 2292 3240 2304
rect 3195 2264 3240 2292
rect 2225 2255 2283 2261
rect 3234 2252 3240 2264
rect 3292 2252 3298 2304
rect 4430 2252 4436 2304
rect 4488 2292 4494 2304
rect 4617 2295 4675 2301
rect 4617 2292 4629 2295
rect 4488 2264 4629 2292
rect 4488 2252 4494 2264
rect 4617 2261 4629 2264
rect 4663 2261 4675 2295
rect 5626 2292 5632 2304
rect 5587 2264 5632 2292
rect 4617 2255 4675 2261
rect 5626 2252 5632 2264
rect 5684 2252 5690 2304
rect 6822 2252 6828 2304
rect 6880 2292 6886 2304
rect 7009 2295 7067 2301
rect 7009 2292 7021 2295
rect 6880 2264 7021 2292
rect 6880 2252 6886 2264
rect 7009 2261 7021 2264
rect 7055 2261 7067 2295
rect 7009 2255 7067 2261
rect 8018 2252 8024 2304
rect 8076 2292 8082 2304
rect 8205 2295 8263 2301
rect 8205 2292 8217 2295
rect 8076 2264 8217 2292
rect 8076 2252 8082 2264
rect 8205 2261 8217 2264
rect 8251 2261 8263 2295
rect 8205 2255 8263 2261
rect 9214 2252 9220 2304
rect 9272 2292 9278 2304
rect 9401 2295 9459 2301
rect 9401 2292 9413 2295
rect 9272 2264 9413 2292
rect 9272 2252 9278 2264
rect 9401 2261 9413 2264
rect 9447 2261 9459 2295
rect 9401 2255 9459 2261
rect 11606 2252 11612 2304
rect 11664 2292 11670 2304
rect 11793 2295 11851 2301
rect 11793 2292 11805 2295
rect 11664 2264 11805 2292
rect 11664 2252 11670 2264
rect 11793 2261 11805 2264
rect 11839 2261 11851 2295
rect 11793 2255 11851 2261
rect 18693 2295 18751 2301
rect 18693 2261 18705 2295
rect 18739 2292 18751 2295
rect 18782 2292 18788 2304
rect 18739 2264 18788 2292
rect 18739 2261 18751 2264
rect 18693 2255 18751 2261
rect 18782 2252 18788 2264
rect 18840 2252 18846 2304
rect 21174 2292 21180 2304
rect 21135 2264 21180 2292
rect 21174 2252 21180 2264
rect 21232 2252 21238 2304
rect 24762 2252 24768 2304
rect 24820 2292 24826 2304
rect 24949 2295 25007 2301
rect 24949 2292 24961 2295
rect 24820 2264 24961 2292
rect 24820 2252 24826 2264
rect 24949 2261 24961 2264
rect 24995 2261 25007 2295
rect 24949 2255 25007 2261
rect 27154 2252 27160 2304
rect 27212 2292 27218 2304
rect 27341 2295 27399 2301
rect 27341 2292 27353 2295
rect 27212 2264 27353 2292
rect 27212 2252 27218 2264
rect 27341 2261 27353 2264
rect 27387 2261 27399 2295
rect 27341 2255 27399 2261
rect 1104 2202 38824 2224
rect 1104 2150 10398 2202
rect 10450 2150 10462 2202
rect 10514 2150 10526 2202
rect 10578 2150 10590 2202
rect 10642 2150 10654 2202
rect 10706 2150 19846 2202
rect 19898 2150 19910 2202
rect 19962 2150 19974 2202
rect 20026 2150 20038 2202
rect 20090 2150 20102 2202
rect 20154 2150 29294 2202
rect 29346 2150 29358 2202
rect 29410 2150 29422 2202
rect 29474 2150 29486 2202
rect 29538 2150 29550 2202
rect 29602 2150 38824 2202
rect 1104 2128 38824 2150
<< via1 >>
rect 10398 33702 10450 33754
rect 10462 33702 10514 33754
rect 10526 33702 10578 33754
rect 10590 33702 10642 33754
rect 10654 33702 10706 33754
rect 19846 33702 19898 33754
rect 19910 33702 19962 33754
rect 19974 33702 20026 33754
rect 20038 33702 20090 33754
rect 20102 33702 20154 33754
rect 29294 33702 29346 33754
rect 29358 33702 29410 33754
rect 29422 33702 29474 33754
rect 29486 33702 29538 33754
rect 29550 33702 29602 33754
rect 8576 33532 8628 33584
rect 9128 33532 9180 33584
rect 14096 33464 14148 33516
rect 20260 33464 20312 33516
rect 25780 33507 25832 33516
rect 25780 33473 25789 33507
rect 25789 33473 25823 33507
rect 25823 33473 25832 33507
rect 25780 33464 25832 33473
rect 31760 33464 31812 33516
rect 37096 33464 37148 33516
rect 1492 33303 1544 33312
rect 1492 33269 1501 33303
rect 1501 33269 1535 33303
rect 1535 33269 1544 33303
rect 1492 33260 1544 33269
rect 9404 33260 9456 33312
rect 5674 33158 5726 33210
rect 5738 33158 5790 33210
rect 5802 33158 5854 33210
rect 5866 33158 5918 33210
rect 5930 33158 5982 33210
rect 15122 33158 15174 33210
rect 15186 33158 15238 33210
rect 15250 33158 15302 33210
rect 15314 33158 15366 33210
rect 15378 33158 15430 33210
rect 24570 33158 24622 33210
rect 24634 33158 24686 33210
rect 24698 33158 24750 33210
rect 24762 33158 24814 33210
rect 24826 33158 24878 33210
rect 34018 33158 34070 33210
rect 34082 33158 34134 33210
rect 34146 33158 34198 33210
rect 34210 33158 34262 33210
rect 34274 33158 34326 33210
rect 1400 33056 1452 33108
rect 9128 33099 9180 33108
rect 9128 33065 9137 33099
rect 9137 33065 9171 33099
rect 9171 33065 9180 33099
rect 9128 33056 9180 33065
rect 9036 32920 9088 32972
rect 12532 32852 12584 32904
rect 2228 32759 2280 32768
rect 2228 32725 2237 32759
rect 2237 32725 2271 32759
rect 2271 32725 2280 32759
rect 2228 32716 2280 32725
rect 10398 32614 10450 32666
rect 10462 32614 10514 32666
rect 10526 32614 10578 32666
rect 10590 32614 10642 32666
rect 10654 32614 10706 32666
rect 19846 32614 19898 32666
rect 19910 32614 19962 32666
rect 19974 32614 20026 32666
rect 20038 32614 20090 32666
rect 20102 32614 20154 32666
rect 29294 32614 29346 32666
rect 29358 32614 29410 32666
rect 29422 32614 29474 32666
rect 29486 32614 29538 32666
rect 29550 32614 29602 32666
rect 2228 32512 2280 32564
rect 12900 32512 12952 32564
rect 3332 32419 3384 32428
rect 3332 32385 3341 32419
rect 3341 32385 3375 32419
rect 3375 32385 3384 32419
rect 3332 32376 3384 32385
rect 3976 32308 4028 32360
rect 9036 32444 9088 32496
rect 17224 32444 17276 32496
rect 6644 32376 6696 32428
rect 11796 32419 11848 32428
rect 11796 32385 11830 32419
rect 11830 32385 11848 32419
rect 11796 32376 11848 32385
rect 16396 32376 16448 32428
rect 1768 32172 1820 32224
rect 4988 32172 5040 32224
rect 8024 32172 8076 32224
rect 10876 32215 10928 32224
rect 10876 32181 10885 32215
rect 10885 32181 10919 32215
rect 10919 32181 10928 32215
rect 10876 32172 10928 32181
rect 12900 32215 12952 32224
rect 12900 32181 12909 32215
rect 12909 32181 12943 32215
rect 12943 32181 12952 32215
rect 12900 32172 12952 32181
rect 18328 32172 18380 32224
rect 22376 32172 22428 32224
rect 5674 32070 5726 32122
rect 5738 32070 5790 32122
rect 5802 32070 5854 32122
rect 5866 32070 5918 32122
rect 5930 32070 5982 32122
rect 15122 32070 15174 32122
rect 15186 32070 15238 32122
rect 15250 32070 15302 32122
rect 15314 32070 15366 32122
rect 15378 32070 15430 32122
rect 24570 32070 24622 32122
rect 24634 32070 24686 32122
rect 24698 32070 24750 32122
rect 24762 32070 24814 32122
rect 24826 32070 24878 32122
rect 34018 32070 34070 32122
rect 34082 32070 34134 32122
rect 34146 32070 34198 32122
rect 34210 32070 34262 32122
rect 34274 32070 34326 32122
rect 3332 31968 3384 32020
rect 6644 32011 6696 32020
rect 6644 31977 6653 32011
rect 6653 31977 6687 32011
rect 6687 31977 6696 32011
rect 6644 31968 6696 31977
rect 18788 31968 18840 32020
rect 8024 31900 8076 31952
rect 11520 31943 11572 31952
rect 11520 31909 11529 31943
rect 11529 31909 11563 31943
rect 11563 31909 11572 31943
rect 11520 31900 11572 31909
rect 16396 31943 16448 31952
rect 16396 31909 16405 31943
rect 16405 31909 16439 31943
rect 16439 31909 16448 31943
rect 16396 31900 16448 31909
rect 18328 31943 18380 31952
rect 18328 31909 18337 31943
rect 18337 31909 18371 31943
rect 18371 31909 18380 31943
rect 18328 31900 18380 31909
rect 12532 31875 12584 31884
rect 12532 31841 12541 31875
rect 12541 31841 12575 31875
rect 12575 31841 12584 31875
rect 12532 31832 12584 31841
rect 2688 31807 2740 31816
rect 2688 31773 2697 31807
rect 2697 31773 2731 31807
rect 2731 31773 2740 31807
rect 2688 31764 2740 31773
rect 6460 31807 6512 31816
rect 6460 31773 6469 31807
rect 6469 31773 6503 31807
rect 6503 31773 6512 31807
rect 6460 31764 6512 31773
rect 9128 31807 9180 31816
rect 9128 31773 9137 31807
rect 9137 31773 9171 31807
rect 9171 31773 9180 31807
rect 9128 31764 9180 31773
rect 12256 31807 12308 31816
rect 12256 31773 12265 31807
rect 12265 31773 12299 31807
rect 12299 31773 12308 31807
rect 12256 31764 12308 31773
rect 16212 31807 16264 31816
rect 16212 31773 16221 31807
rect 16221 31773 16255 31807
rect 16255 31773 16264 31807
rect 16212 31764 16264 31773
rect 17224 31764 17276 31816
rect 17592 31807 17644 31816
rect 17592 31773 17601 31807
rect 17601 31773 17635 31807
rect 17635 31773 17644 31807
rect 17592 31764 17644 31773
rect 20720 31807 20772 31816
rect 20720 31773 20729 31807
rect 20729 31773 20763 31807
rect 20763 31773 20772 31807
rect 20720 31764 20772 31773
rect 23480 31968 23532 32020
rect 22376 31943 22428 31952
rect 22376 31909 22385 31943
rect 22385 31909 22419 31943
rect 22419 31909 22428 31943
rect 22376 31900 22428 31909
rect 25412 31968 25464 32020
rect 29000 32011 29052 32020
rect 29000 31977 29009 32011
rect 29009 31977 29043 32011
rect 29043 31977 29052 32011
rect 29000 31968 29052 31977
rect 22100 31764 22152 31816
rect 25044 31807 25096 31816
rect 25044 31773 25053 31807
rect 25053 31773 25087 31807
rect 25087 31773 25096 31807
rect 25044 31764 25096 31773
rect 25320 31807 25372 31816
rect 25320 31773 25329 31807
rect 25329 31773 25363 31807
rect 25363 31773 25372 31807
rect 25320 31764 25372 31773
rect 28264 31807 28316 31816
rect 28264 31773 28273 31807
rect 28273 31773 28307 31807
rect 28307 31773 28316 31807
rect 28264 31764 28316 31773
rect 28172 31696 28224 31748
rect 1492 31671 1544 31680
rect 1492 31637 1501 31671
rect 1501 31637 1535 31671
rect 1535 31637 1544 31671
rect 1492 31628 1544 31637
rect 8760 31628 8812 31680
rect 10398 31526 10450 31578
rect 10462 31526 10514 31578
rect 10526 31526 10578 31578
rect 10590 31526 10642 31578
rect 10654 31526 10706 31578
rect 19846 31526 19898 31578
rect 19910 31526 19962 31578
rect 19974 31526 20026 31578
rect 20038 31526 20090 31578
rect 20102 31526 20154 31578
rect 29294 31526 29346 31578
rect 29358 31526 29410 31578
rect 29422 31526 29474 31578
rect 29486 31526 29538 31578
rect 29550 31526 29602 31578
rect 2688 31467 2740 31476
rect 2688 31433 2697 31467
rect 2697 31433 2731 31467
rect 2731 31433 2740 31467
rect 2688 31424 2740 31433
rect 6460 31424 6512 31476
rect 8024 31467 8076 31476
rect 8024 31433 8033 31467
rect 8033 31433 8067 31467
rect 8067 31433 8076 31467
rect 8024 31424 8076 31433
rect 12256 31424 12308 31476
rect 16212 31424 16264 31476
rect 17592 31424 17644 31476
rect 20720 31424 20772 31476
rect 22100 31424 22152 31476
rect 29000 31424 29052 31476
rect 3424 31288 3476 31340
rect 6552 31331 6604 31340
rect 6552 31297 6561 31331
rect 6561 31297 6595 31331
rect 6595 31297 6604 31331
rect 6552 31288 6604 31297
rect 8760 31331 8812 31340
rect 8760 31297 8769 31331
rect 8769 31297 8803 31331
rect 8803 31297 8812 31331
rect 8760 31288 8812 31297
rect 9036 31331 9088 31340
rect 9036 31297 9045 31331
rect 9045 31297 9079 31331
rect 9079 31297 9088 31331
rect 9036 31288 9088 31297
rect 11704 31331 11756 31340
rect 11704 31297 11713 31331
rect 11713 31297 11747 31331
rect 11747 31297 11756 31331
rect 11704 31288 11756 31297
rect 15844 31331 15896 31340
rect 15844 31297 15853 31331
rect 15853 31297 15887 31331
rect 15887 31297 15896 31331
rect 15844 31288 15896 31297
rect 21180 31288 21232 31340
rect 21364 31288 21416 31340
rect 29552 31288 29604 31340
rect 3148 31220 3200 31272
rect 6920 31220 6972 31272
rect 13176 31220 13228 31272
rect 15660 31263 15712 31272
rect 15660 31229 15669 31263
rect 15669 31229 15703 31263
rect 15703 31229 15712 31263
rect 15660 31220 15712 31229
rect 19524 31220 19576 31272
rect 28172 31220 28224 31272
rect 5674 30982 5726 31034
rect 5738 30982 5790 31034
rect 5802 30982 5854 31034
rect 5866 30982 5918 31034
rect 5930 30982 5982 31034
rect 15122 30982 15174 31034
rect 15186 30982 15238 31034
rect 15250 30982 15302 31034
rect 15314 30982 15366 31034
rect 15378 30982 15430 31034
rect 24570 30982 24622 31034
rect 24634 30982 24686 31034
rect 24698 30982 24750 31034
rect 24762 30982 24814 31034
rect 24826 30982 24878 31034
rect 34018 30982 34070 31034
rect 34082 30982 34134 31034
rect 34146 30982 34198 31034
rect 34210 30982 34262 31034
rect 34274 30982 34326 31034
rect 4988 30923 5040 30932
rect 4988 30889 4997 30923
rect 4997 30889 5031 30923
rect 5031 30889 5040 30923
rect 4988 30880 5040 30889
rect 9128 30880 9180 30932
rect 15660 30880 15712 30932
rect 21364 30923 21416 30932
rect 21364 30889 21373 30923
rect 21373 30889 21407 30923
rect 21407 30889 21416 30923
rect 21364 30880 21416 30889
rect 25044 30880 25096 30932
rect 25320 30880 25372 30932
rect 28264 30880 28316 30932
rect 29552 30923 29604 30932
rect 29552 30889 29561 30923
rect 29561 30889 29595 30923
rect 29595 30889 29604 30923
rect 29552 30880 29604 30889
rect 3976 30787 4028 30796
rect 3976 30753 3985 30787
rect 3985 30753 4019 30787
rect 4019 30753 4028 30787
rect 3976 30744 4028 30753
rect 6920 30744 6972 30796
rect 12716 30744 12768 30796
rect 13176 30744 13228 30796
rect 1676 30719 1728 30728
rect 1676 30685 1685 30719
rect 1685 30685 1719 30719
rect 1719 30685 1728 30719
rect 1676 30676 1728 30685
rect 4252 30719 4304 30728
rect 4252 30685 4261 30719
rect 4261 30685 4295 30719
rect 4295 30685 4304 30719
rect 4252 30676 4304 30685
rect 6552 30676 6604 30728
rect 9864 30676 9916 30728
rect 20812 30676 20864 30728
rect 21180 30719 21232 30728
rect 11796 30608 11848 30660
rect 21180 30685 21189 30719
rect 21189 30685 21223 30719
rect 21223 30685 21232 30719
rect 21180 30676 21232 30685
rect 23940 30744 23992 30796
rect 24492 30676 24544 30728
rect 25228 30719 25280 30728
rect 25228 30685 25237 30719
rect 25237 30685 25271 30719
rect 25271 30685 25280 30719
rect 25228 30676 25280 30685
rect 28816 30719 28868 30728
rect 28816 30685 28825 30719
rect 28825 30685 28859 30719
rect 28859 30685 28868 30719
rect 28816 30676 28868 30685
rect 29736 30719 29788 30728
rect 29736 30685 29745 30719
rect 29745 30685 29779 30719
rect 29779 30685 29788 30719
rect 29736 30676 29788 30685
rect 1492 30583 1544 30592
rect 1492 30549 1501 30583
rect 1501 30549 1535 30583
rect 1535 30549 1544 30583
rect 1492 30540 1544 30549
rect 9864 30583 9916 30592
rect 9864 30549 9873 30583
rect 9873 30549 9907 30583
rect 9907 30549 9916 30583
rect 9864 30540 9916 30549
rect 10398 30438 10450 30490
rect 10462 30438 10514 30490
rect 10526 30438 10578 30490
rect 10590 30438 10642 30490
rect 10654 30438 10706 30490
rect 19846 30438 19898 30490
rect 19910 30438 19962 30490
rect 19974 30438 20026 30490
rect 20038 30438 20090 30490
rect 20102 30438 20154 30490
rect 29294 30438 29346 30490
rect 29358 30438 29410 30490
rect 29422 30438 29474 30490
rect 29486 30438 29538 30490
rect 29550 30438 29602 30490
rect 4252 30379 4304 30388
rect 4252 30345 4261 30379
rect 4261 30345 4295 30379
rect 4295 30345 4304 30379
rect 4252 30336 4304 30345
rect 11704 30336 11756 30388
rect 3424 30243 3476 30252
rect 3424 30209 3433 30243
rect 3433 30209 3467 30243
rect 3467 30209 3476 30243
rect 3424 30200 3476 30209
rect 12440 30200 12492 30252
rect 24400 30200 24452 30252
rect 4160 30132 4212 30184
rect 13820 30132 13872 30184
rect 24492 30175 24544 30184
rect 24492 30141 24501 30175
rect 24501 30141 24535 30175
rect 24535 30141 24544 30175
rect 24492 30132 24544 30141
rect 12440 30039 12492 30048
rect 12440 30005 12449 30039
rect 12449 30005 12483 30039
rect 12483 30005 12492 30039
rect 12440 29996 12492 30005
rect 25412 29996 25464 30048
rect 5674 29894 5726 29946
rect 5738 29894 5790 29946
rect 5802 29894 5854 29946
rect 5866 29894 5918 29946
rect 5930 29894 5982 29946
rect 15122 29894 15174 29946
rect 15186 29894 15238 29946
rect 15250 29894 15302 29946
rect 15314 29894 15366 29946
rect 15378 29894 15430 29946
rect 24570 29894 24622 29946
rect 24634 29894 24686 29946
rect 24698 29894 24750 29946
rect 24762 29894 24814 29946
rect 24826 29894 24878 29946
rect 34018 29894 34070 29946
rect 34082 29894 34134 29946
rect 34146 29894 34198 29946
rect 34210 29894 34262 29946
rect 34274 29894 34326 29946
rect 1676 29792 1728 29844
rect 11520 29792 11572 29844
rect 25228 29792 25280 29844
rect 28816 29792 28868 29844
rect 23940 29656 23992 29708
rect 24768 29699 24820 29708
rect 24768 29665 24777 29699
rect 24777 29665 24811 29699
rect 24811 29665 24820 29699
rect 24768 29656 24820 29665
rect 2964 29588 3016 29640
rect 12532 29631 12584 29640
rect 12532 29597 12541 29631
rect 12541 29597 12575 29631
rect 12575 29597 12584 29631
rect 12532 29588 12584 29597
rect 12624 29588 12676 29640
rect 24124 29588 24176 29640
rect 24768 29520 24820 29572
rect 28908 29588 28960 29640
rect 4160 29452 4212 29504
rect 4620 29452 4672 29504
rect 31392 29520 31444 29572
rect 32680 29452 32732 29504
rect 10398 29350 10450 29402
rect 10462 29350 10514 29402
rect 10526 29350 10578 29402
rect 10590 29350 10642 29402
rect 10654 29350 10706 29402
rect 19846 29350 19898 29402
rect 19910 29350 19962 29402
rect 19974 29350 20026 29402
rect 20038 29350 20090 29402
rect 20102 29350 20154 29402
rect 29294 29350 29346 29402
rect 29358 29350 29410 29402
rect 29422 29350 29474 29402
rect 29486 29350 29538 29402
rect 29550 29350 29602 29402
rect 12532 29248 12584 29300
rect 24400 29248 24452 29300
rect 29736 29248 29788 29300
rect 31392 29291 31444 29300
rect 31392 29257 31401 29291
rect 31401 29257 31435 29291
rect 31435 29257 31444 29291
rect 31392 29248 31444 29257
rect 32680 29291 32732 29300
rect 32680 29257 32689 29291
rect 32689 29257 32723 29291
rect 32723 29257 32732 29291
rect 32680 29248 32732 29257
rect 34796 29248 34848 29300
rect 11796 29155 11848 29164
rect 11796 29121 11805 29155
rect 11805 29121 11839 29155
rect 11839 29121 11848 29155
rect 11796 29112 11848 29121
rect 12992 29155 13044 29164
rect 12992 29121 13001 29155
rect 13001 29121 13035 29155
rect 13035 29121 13044 29155
rect 12992 29112 13044 29121
rect 15844 29155 15896 29164
rect 15844 29121 15853 29155
rect 15853 29121 15887 29155
rect 15887 29121 15896 29155
rect 15844 29112 15896 29121
rect 17500 29155 17552 29164
rect 17500 29121 17509 29155
rect 17509 29121 17543 29155
rect 17543 29121 17552 29155
rect 17500 29112 17552 29121
rect 24952 29155 25004 29164
rect 24952 29121 24961 29155
rect 24961 29121 24995 29155
rect 24995 29121 25004 29155
rect 24952 29112 25004 29121
rect 28908 29155 28960 29164
rect 28908 29121 28917 29155
rect 28917 29121 28951 29155
rect 28951 29121 28960 29155
rect 28908 29112 28960 29121
rect 31300 29155 31352 29164
rect 31300 29121 31309 29155
rect 31309 29121 31343 29155
rect 31343 29121 31352 29155
rect 31300 29112 31352 29121
rect 32312 29112 32364 29164
rect 12440 29044 12492 29096
rect 13820 29044 13872 29096
rect 17224 29087 17276 29096
rect 17224 29053 17233 29087
rect 17233 29053 17267 29087
rect 17267 29053 17276 29087
rect 17224 29044 17276 29053
rect 31208 29044 31260 29096
rect 1492 29019 1544 29028
rect 1492 28985 1501 29019
rect 1501 28985 1535 29019
rect 1535 28985 1544 29019
rect 1492 28976 1544 28985
rect 2044 28976 2096 29028
rect 2964 29019 3016 29028
rect 2964 28985 2973 29019
rect 2973 28985 3007 29019
rect 3007 28985 3016 29019
rect 2964 28976 3016 28985
rect 16672 28976 16724 29028
rect 18328 28976 18380 29028
rect 19432 28976 19484 29028
rect 13452 28951 13504 28960
rect 13452 28917 13461 28951
rect 13461 28917 13495 28951
rect 13495 28917 13504 28951
rect 13452 28908 13504 28917
rect 5674 28806 5726 28858
rect 5738 28806 5790 28858
rect 5802 28806 5854 28858
rect 5866 28806 5918 28858
rect 5930 28806 5982 28858
rect 15122 28806 15174 28858
rect 15186 28806 15238 28858
rect 15250 28806 15302 28858
rect 15314 28806 15366 28858
rect 15378 28806 15430 28858
rect 24570 28806 24622 28858
rect 24634 28806 24686 28858
rect 24698 28806 24750 28858
rect 24762 28806 24814 28858
rect 24826 28806 24878 28858
rect 34018 28806 34070 28858
rect 34082 28806 34134 28858
rect 34146 28806 34198 28858
rect 34210 28806 34262 28858
rect 34274 28806 34326 28858
rect 12992 28704 13044 28756
rect 17500 28704 17552 28756
rect 34796 28747 34848 28756
rect 34796 28713 34805 28747
rect 34805 28713 34839 28747
rect 34839 28713 34848 28747
rect 34796 28704 34848 28713
rect 17224 28636 17276 28688
rect 9128 28543 9180 28552
rect 9128 28509 9137 28543
rect 9137 28509 9171 28543
rect 9171 28509 9180 28543
rect 9128 28500 9180 28509
rect 12256 28543 12308 28552
rect 12256 28509 12265 28543
rect 12265 28509 12299 28543
rect 12299 28509 12308 28543
rect 12256 28500 12308 28509
rect 12440 28568 12492 28620
rect 13452 28568 13504 28620
rect 13820 28568 13872 28620
rect 21180 28568 21232 28620
rect 14004 28500 14056 28552
rect 14096 28543 14148 28552
rect 14096 28509 14105 28543
rect 14105 28509 14139 28543
rect 14139 28509 14148 28543
rect 16672 28543 16724 28552
rect 14096 28500 14148 28509
rect 16672 28509 16681 28543
rect 16681 28509 16715 28543
rect 16715 28509 16724 28543
rect 16672 28500 16724 28509
rect 20720 28543 20772 28552
rect 8392 28364 8444 28416
rect 12624 28364 12676 28416
rect 20720 28509 20729 28543
rect 20729 28509 20763 28543
rect 20763 28509 20772 28543
rect 20720 28500 20772 28509
rect 21272 28432 21324 28484
rect 31300 28432 31352 28484
rect 31576 28475 31628 28484
rect 31576 28441 31585 28475
rect 31585 28441 31619 28475
rect 31619 28441 31628 28475
rect 31576 28432 31628 28441
rect 32312 28407 32364 28416
rect 32312 28373 32321 28407
rect 32321 28373 32355 28407
rect 32355 28373 32364 28407
rect 32312 28364 32364 28373
rect 10398 28262 10450 28314
rect 10462 28262 10514 28314
rect 10526 28262 10578 28314
rect 10590 28262 10642 28314
rect 10654 28262 10706 28314
rect 19846 28262 19898 28314
rect 19910 28262 19962 28314
rect 19974 28262 20026 28314
rect 20038 28262 20090 28314
rect 20102 28262 20154 28314
rect 29294 28262 29346 28314
rect 29358 28262 29410 28314
rect 29422 28262 29474 28314
rect 29486 28262 29538 28314
rect 29550 28262 29602 28314
rect 24952 28203 25004 28212
rect 24952 28169 24961 28203
rect 24961 28169 24995 28203
rect 24995 28169 25004 28203
rect 24952 28160 25004 28169
rect 29000 28160 29052 28212
rect 32312 28092 32364 28144
rect 8392 28067 8444 28076
rect 1492 27863 1544 27872
rect 1492 27829 1501 27863
rect 1501 27829 1535 27863
rect 1535 27829 1544 27863
rect 1492 27820 1544 27829
rect 8392 28033 8401 28067
rect 8401 28033 8435 28067
rect 8435 28033 8444 28067
rect 8392 28024 8444 28033
rect 20996 28067 21048 28076
rect 20996 28033 21005 28067
rect 21005 28033 21039 28067
rect 21039 28033 21048 28067
rect 20996 28024 21048 28033
rect 21272 28067 21324 28076
rect 21272 28033 21281 28067
rect 21281 28033 21315 28067
rect 21315 28033 21324 28067
rect 21272 28024 21324 28033
rect 8116 27999 8168 28008
rect 8116 27965 8125 27999
rect 8125 27965 8159 27999
rect 8159 27965 8168 27999
rect 8116 27956 8168 27965
rect 24124 28024 24176 28076
rect 28172 28067 28224 28076
rect 28172 28033 28181 28067
rect 28181 28033 28215 28067
rect 28215 28033 28224 28067
rect 28172 28024 28224 28033
rect 28448 28067 28500 28076
rect 28448 28033 28457 28067
rect 28457 28033 28491 28067
rect 28491 28033 28500 28067
rect 28448 28024 28500 28033
rect 31852 28024 31904 28076
rect 23480 27956 23532 28008
rect 12256 27888 12308 27940
rect 19340 27888 19392 27940
rect 19432 27888 19484 27940
rect 31208 27956 31260 28008
rect 34520 27956 34572 28008
rect 34796 27956 34848 28008
rect 2320 27820 2372 27872
rect 8392 27820 8444 27872
rect 13452 27863 13504 27872
rect 13452 27829 13461 27863
rect 13461 27829 13495 27863
rect 13495 27829 13504 27863
rect 13452 27820 13504 27829
rect 19708 27863 19760 27872
rect 19708 27829 19717 27863
rect 19717 27829 19751 27863
rect 19751 27829 19760 27863
rect 19708 27820 19760 27829
rect 24308 27820 24360 27872
rect 34980 27820 35032 27872
rect 35900 27820 35952 27872
rect 5674 27718 5726 27770
rect 5738 27718 5790 27770
rect 5802 27718 5854 27770
rect 5866 27718 5918 27770
rect 5930 27718 5982 27770
rect 15122 27718 15174 27770
rect 15186 27718 15238 27770
rect 15250 27718 15302 27770
rect 15314 27718 15366 27770
rect 15378 27718 15430 27770
rect 24570 27718 24622 27770
rect 24634 27718 24686 27770
rect 24698 27718 24750 27770
rect 24762 27718 24814 27770
rect 24826 27718 24878 27770
rect 34018 27718 34070 27770
rect 34082 27718 34134 27770
rect 34146 27718 34198 27770
rect 34210 27718 34262 27770
rect 34274 27718 34326 27770
rect 3056 27548 3108 27600
rect 9128 27616 9180 27668
rect 20996 27659 21048 27668
rect 20996 27625 21005 27659
rect 21005 27625 21039 27659
rect 21039 27625 21048 27659
rect 20996 27616 21048 27625
rect 8392 27548 8444 27600
rect 23480 27548 23532 27600
rect 31392 27548 31444 27600
rect 2872 27412 2924 27464
rect 5080 27455 5132 27464
rect 5080 27421 5089 27455
rect 5089 27421 5123 27455
rect 5123 27421 5132 27455
rect 5080 27412 5132 27421
rect 5540 27412 5592 27464
rect 6736 27455 6788 27464
rect 6736 27421 6745 27455
rect 6745 27421 6779 27455
rect 6779 27421 6788 27455
rect 6736 27412 6788 27421
rect 6920 27455 6972 27464
rect 6920 27421 6929 27455
rect 6929 27421 6963 27455
rect 6963 27421 6972 27455
rect 24124 27480 24176 27532
rect 6920 27412 6972 27421
rect 9220 27412 9272 27464
rect 5724 27344 5776 27396
rect 7380 27344 7432 27396
rect 8116 27344 8168 27396
rect 3240 27276 3292 27328
rect 6552 27319 6604 27328
rect 6552 27285 6561 27319
rect 6561 27285 6595 27319
rect 6595 27285 6604 27319
rect 6552 27276 6604 27285
rect 9864 27319 9916 27328
rect 9864 27285 9873 27319
rect 9873 27285 9907 27319
rect 9907 27285 9916 27319
rect 9864 27276 9916 27285
rect 19340 27276 19392 27328
rect 28540 27455 28592 27464
rect 28540 27421 28549 27455
rect 28549 27421 28583 27455
rect 28583 27421 28592 27455
rect 28540 27412 28592 27421
rect 34980 27455 35032 27464
rect 34980 27421 34989 27455
rect 34989 27421 35023 27455
rect 35023 27421 35032 27455
rect 34980 27412 35032 27421
rect 35624 27455 35676 27464
rect 35624 27421 35633 27455
rect 35633 27421 35667 27455
rect 35667 27421 35676 27455
rect 35624 27412 35676 27421
rect 36728 27455 36780 27464
rect 20720 27344 20772 27396
rect 24952 27387 25004 27396
rect 24952 27353 24961 27387
rect 24961 27353 24995 27387
rect 24995 27353 25004 27387
rect 24952 27344 25004 27353
rect 36728 27421 36737 27455
rect 36737 27421 36771 27455
rect 36771 27421 36780 27455
rect 36728 27412 36780 27421
rect 28724 27276 28776 27328
rect 10398 27174 10450 27226
rect 10462 27174 10514 27226
rect 10526 27174 10578 27226
rect 10590 27174 10642 27226
rect 10654 27174 10706 27226
rect 19846 27174 19898 27226
rect 19910 27174 19962 27226
rect 19974 27174 20026 27226
rect 20038 27174 20090 27226
rect 20102 27174 20154 27226
rect 29294 27174 29346 27226
rect 29358 27174 29410 27226
rect 29422 27174 29474 27226
rect 29486 27174 29538 27226
rect 29550 27174 29602 27226
rect 3056 27072 3108 27124
rect 5540 27115 5592 27124
rect 5540 27081 5549 27115
rect 5549 27081 5583 27115
rect 5583 27081 5592 27115
rect 5540 27072 5592 27081
rect 24124 27115 24176 27124
rect 24124 27081 24133 27115
rect 24133 27081 24167 27115
rect 24167 27081 24176 27115
rect 24124 27072 24176 27081
rect 28448 27072 28500 27124
rect 3976 27004 4028 27056
rect 6736 27004 6788 27056
rect 3240 26979 3292 26988
rect 3240 26945 3249 26979
rect 3249 26945 3283 26979
rect 3283 26945 3292 26979
rect 3240 26936 3292 26945
rect 5080 26936 5132 26988
rect 5632 26936 5684 26988
rect 6552 26936 6604 26988
rect 7840 26979 7892 26988
rect 7840 26945 7849 26979
rect 7849 26945 7883 26979
rect 7883 26945 7892 26979
rect 7840 26936 7892 26945
rect 23572 26936 23624 26988
rect 28724 26979 28776 26988
rect 28724 26945 28733 26979
rect 28733 26945 28767 26979
rect 28767 26945 28776 26979
rect 28724 26936 28776 26945
rect 30656 26936 30708 26988
rect 31300 26979 31352 26988
rect 31300 26945 31309 26979
rect 31309 26945 31343 26979
rect 31343 26945 31352 26979
rect 31300 26936 31352 26945
rect 31852 26936 31904 26988
rect 32956 26979 33008 26988
rect 32956 26945 32965 26979
rect 32965 26945 32999 26979
rect 32999 26945 33008 26979
rect 32956 26936 33008 26945
rect 35900 26979 35952 26988
rect 35900 26945 35909 26979
rect 35909 26945 35943 26979
rect 35943 26945 35952 26979
rect 36728 26979 36780 26988
rect 35900 26936 35952 26945
rect 36728 26945 36737 26979
rect 36737 26945 36771 26979
rect 36771 26945 36780 26979
rect 36728 26936 36780 26945
rect 33784 26868 33836 26920
rect 35624 26911 35676 26920
rect 35624 26877 35633 26911
rect 35633 26877 35667 26911
rect 35667 26877 35676 26911
rect 35624 26868 35676 26877
rect 7656 26775 7708 26784
rect 7656 26741 7665 26775
rect 7665 26741 7699 26775
rect 7699 26741 7708 26775
rect 7656 26732 7708 26741
rect 9864 26732 9916 26784
rect 14924 26732 14976 26784
rect 19524 26732 19576 26784
rect 20720 26732 20772 26784
rect 21272 26732 21324 26784
rect 31668 26732 31720 26784
rect 33876 26732 33928 26784
rect 5674 26630 5726 26682
rect 5738 26630 5790 26682
rect 5802 26630 5854 26682
rect 5866 26630 5918 26682
rect 5930 26630 5982 26682
rect 15122 26630 15174 26682
rect 15186 26630 15238 26682
rect 15250 26630 15302 26682
rect 15314 26630 15366 26682
rect 15378 26630 15430 26682
rect 24570 26630 24622 26682
rect 24634 26630 24686 26682
rect 24698 26630 24750 26682
rect 24762 26630 24814 26682
rect 24826 26630 24878 26682
rect 34018 26630 34070 26682
rect 34082 26630 34134 26682
rect 34146 26630 34198 26682
rect 34210 26630 34262 26682
rect 34274 26630 34326 26682
rect 2872 26571 2924 26580
rect 2872 26537 2881 26571
rect 2881 26537 2915 26571
rect 2915 26537 2924 26571
rect 2872 26528 2924 26537
rect 8392 26571 8444 26580
rect 8392 26537 8401 26571
rect 8401 26537 8435 26571
rect 8435 26537 8444 26571
rect 8392 26528 8444 26537
rect 14004 26528 14056 26580
rect 32956 26528 33008 26580
rect 7380 26435 7432 26444
rect 7380 26401 7389 26435
rect 7389 26401 7423 26435
rect 7423 26401 7432 26435
rect 7380 26392 7432 26401
rect 14924 26435 14976 26444
rect 14924 26401 14933 26435
rect 14933 26401 14967 26435
rect 14967 26401 14976 26435
rect 14924 26392 14976 26401
rect 2412 26367 2464 26376
rect 2412 26333 2421 26367
rect 2421 26333 2455 26367
rect 2455 26333 2464 26367
rect 2412 26324 2464 26333
rect 2964 26324 3016 26376
rect 3148 26367 3200 26376
rect 3148 26333 3157 26367
rect 3157 26333 3191 26367
rect 3191 26333 3200 26367
rect 3148 26324 3200 26333
rect 3884 26324 3936 26376
rect 7656 26367 7708 26376
rect 7656 26333 7665 26367
rect 7665 26333 7699 26367
rect 7699 26333 7708 26367
rect 7656 26324 7708 26333
rect 12348 26367 12400 26376
rect 12348 26333 12357 26367
rect 12357 26333 12391 26367
rect 12391 26333 12400 26367
rect 12348 26324 12400 26333
rect 15016 26324 15068 26376
rect 15568 26324 15620 26376
rect 16028 26367 16080 26376
rect 16028 26333 16037 26367
rect 16037 26333 16071 26367
rect 16071 26333 16080 26367
rect 16028 26324 16080 26333
rect 21824 26324 21876 26376
rect 24860 26367 24912 26376
rect 24860 26333 24869 26367
rect 24869 26333 24903 26367
rect 24903 26333 24912 26367
rect 24860 26324 24912 26333
rect 31668 26367 31720 26376
rect 31668 26333 31677 26367
rect 31677 26333 31711 26367
rect 31711 26333 31720 26367
rect 31668 26324 31720 26333
rect 3976 26256 4028 26308
rect 19616 26299 19668 26308
rect 19616 26265 19625 26299
rect 19625 26265 19659 26299
rect 19659 26265 19668 26299
rect 19616 26256 19668 26265
rect 1492 26231 1544 26240
rect 1492 26197 1501 26231
rect 1501 26197 1535 26231
rect 1535 26197 1544 26231
rect 1492 26188 1544 26197
rect 12164 26231 12216 26240
rect 12164 26197 12173 26231
rect 12173 26197 12207 26231
rect 12207 26197 12216 26231
rect 12164 26188 12216 26197
rect 15752 26188 15804 26240
rect 17040 26188 17092 26240
rect 25044 26231 25096 26240
rect 25044 26197 25053 26231
rect 25053 26197 25087 26231
rect 25087 26197 25096 26231
rect 25044 26188 25096 26197
rect 10398 26086 10450 26138
rect 10462 26086 10514 26138
rect 10526 26086 10578 26138
rect 10590 26086 10642 26138
rect 10654 26086 10706 26138
rect 19846 26086 19898 26138
rect 19910 26086 19962 26138
rect 19974 26086 20026 26138
rect 20038 26086 20090 26138
rect 20102 26086 20154 26138
rect 29294 26086 29346 26138
rect 29358 26086 29410 26138
rect 29422 26086 29474 26138
rect 29486 26086 29538 26138
rect 29550 26086 29602 26138
rect 7840 25984 7892 26036
rect 16028 25984 16080 26036
rect 24860 25984 24912 26036
rect 9220 25848 9272 25900
rect 12164 25848 12216 25900
rect 15752 25891 15804 25900
rect 15752 25857 15761 25891
rect 15761 25857 15795 25891
rect 15795 25857 15804 25891
rect 15752 25848 15804 25857
rect 25044 25891 25096 25900
rect 25044 25857 25053 25891
rect 25053 25857 25087 25891
rect 25087 25857 25096 25891
rect 25044 25848 25096 25857
rect 25964 25891 26016 25900
rect 25964 25857 25973 25891
rect 25973 25857 26007 25891
rect 26007 25857 26016 25891
rect 25964 25848 26016 25857
rect 28448 25891 28500 25900
rect 28448 25857 28457 25891
rect 28457 25857 28491 25891
rect 28491 25857 28500 25891
rect 28448 25848 28500 25857
rect 7380 25823 7432 25832
rect 7380 25789 7389 25823
rect 7389 25789 7423 25823
rect 7423 25789 7432 25823
rect 7380 25780 7432 25789
rect 11704 25823 11756 25832
rect 11704 25789 11713 25823
rect 11713 25789 11747 25823
rect 11747 25789 11756 25823
rect 11704 25780 11756 25789
rect 25320 25823 25372 25832
rect 25320 25789 25329 25823
rect 25329 25789 25363 25823
rect 25363 25789 25372 25823
rect 25320 25780 25372 25789
rect 2412 25644 2464 25696
rect 4344 25644 4396 25696
rect 12440 25644 12492 25696
rect 17040 25644 17092 25696
rect 22836 25644 22888 25696
rect 30656 25780 30708 25832
rect 27712 25712 27764 25764
rect 27804 25644 27856 25696
rect 5674 25542 5726 25594
rect 5738 25542 5790 25594
rect 5802 25542 5854 25594
rect 5866 25542 5918 25594
rect 5930 25542 5982 25594
rect 15122 25542 15174 25594
rect 15186 25542 15238 25594
rect 15250 25542 15302 25594
rect 15314 25542 15366 25594
rect 15378 25542 15430 25594
rect 24570 25542 24622 25594
rect 24634 25542 24686 25594
rect 24698 25542 24750 25594
rect 24762 25542 24814 25594
rect 24826 25542 24878 25594
rect 34018 25542 34070 25594
rect 34082 25542 34134 25594
rect 34146 25542 34198 25594
rect 34210 25542 34262 25594
rect 34274 25542 34326 25594
rect 12348 25440 12400 25492
rect 21824 25440 21876 25492
rect 12716 25304 12768 25356
rect 15568 25347 15620 25356
rect 15568 25313 15577 25347
rect 15577 25313 15611 25347
rect 15611 25313 15620 25347
rect 15568 25304 15620 25313
rect 21824 25347 21876 25356
rect 21824 25313 21833 25347
rect 21833 25313 21867 25347
rect 21867 25313 21876 25347
rect 21824 25304 21876 25313
rect 15016 25236 15068 25288
rect 15844 25279 15896 25288
rect 15844 25245 15853 25279
rect 15853 25245 15887 25279
rect 15887 25245 15896 25279
rect 15844 25236 15896 25245
rect 1492 25143 1544 25152
rect 1492 25109 1501 25143
rect 1501 25109 1535 25143
rect 1535 25109 1544 25143
rect 1492 25100 1544 25109
rect 2228 25143 2280 25152
rect 2228 25109 2237 25143
rect 2237 25109 2271 25143
rect 2271 25109 2280 25143
rect 2228 25100 2280 25109
rect 17040 25100 17092 25152
rect 19708 25100 19760 25152
rect 20536 25236 20588 25288
rect 20996 25279 21048 25288
rect 20996 25245 21005 25279
rect 21005 25245 21039 25279
rect 21039 25245 21048 25279
rect 22100 25279 22152 25288
rect 20996 25236 21048 25245
rect 22100 25245 22109 25279
rect 22109 25245 22143 25279
rect 22143 25245 22152 25279
rect 22100 25236 22152 25245
rect 25320 25236 25372 25288
rect 27804 25279 27856 25288
rect 25964 25168 26016 25220
rect 27804 25245 27813 25279
rect 27813 25245 27847 25279
rect 27847 25245 27856 25279
rect 27804 25236 27856 25245
rect 27712 25168 27764 25220
rect 21824 25100 21876 25152
rect 22836 25143 22888 25152
rect 22836 25109 22845 25143
rect 22845 25109 22879 25143
rect 22879 25109 22888 25143
rect 22836 25100 22888 25109
rect 28724 25100 28776 25152
rect 10398 24998 10450 25050
rect 10462 24998 10514 25050
rect 10526 24998 10578 25050
rect 10590 24998 10642 25050
rect 10654 24998 10706 25050
rect 19846 24998 19898 25050
rect 19910 24998 19962 25050
rect 19974 24998 20026 25050
rect 20038 24998 20090 25050
rect 20102 24998 20154 25050
rect 29294 24998 29346 25050
rect 29358 24998 29410 25050
rect 29422 24998 29474 25050
rect 29486 24998 29538 25050
rect 29550 24998 29602 25050
rect 2228 24896 2280 24948
rect 13268 24896 13320 24948
rect 15844 24896 15896 24948
rect 28448 24896 28500 24948
rect 2320 24760 2372 24812
rect 12716 24556 12768 24608
rect 13544 24556 13596 24608
rect 15016 24760 15068 24812
rect 19616 24760 19668 24812
rect 21824 24803 21876 24812
rect 21824 24769 21833 24803
rect 21833 24769 21867 24803
rect 21867 24769 21876 24803
rect 21824 24760 21876 24769
rect 25964 24760 26016 24812
rect 28632 24760 28684 24812
rect 32956 24803 33008 24812
rect 32956 24769 32965 24803
rect 32965 24769 32999 24803
rect 32999 24769 33008 24803
rect 32956 24760 33008 24769
rect 20996 24624 21048 24676
rect 31208 24692 31260 24744
rect 32864 24692 32916 24744
rect 30564 24624 30616 24676
rect 15660 24556 15712 24608
rect 22100 24556 22152 24608
rect 33140 24599 33192 24608
rect 33140 24565 33149 24599
rect 33149 24565 33183 24599
rect 33183 24565 33192 24599
rect 33140 24556 33192 24565
rect 33784 24599 33836 24608
rect 33784 24565 33793 24599
rect 33793 24565 33827 24599
rect 33827 24565 33836 24599
rect 33784 24556 33836 24565
rect 5674 24454 5726 24506
rect 5738 24454 5790 24506
rect 5802 24454 5854 24506
rect 5866 24454 5918 24506
rect 5930 24454 5982 24506
rect 15122 24454 15174 24506
rect 15186 24454 15238 24506
rect 15250 24454 15302 24506
rect 15314 24454 15366 24506
rect 15378 24454 15430 24506
rect 24570 24454 24622 24506
rect 24634 24454 24686 24506
rect 24698 24454 24750 24506
rect 24762 24454 24814 24506
rect 24826 24454 24878 24506
rect 34018 24454 34070 24506
rect 34082 24454 34134 24506
rect 34146 24454 34198 24506
rect 34210 24454 34262 24506
rect 34274 24454 34326 24506
rect 3976 24191 4028 24200
rect 3976 24157 3985 24191
rect 3985 24157 4019 24191
rect 4019 24157 4028 24191
rect 3976 24148 4028 24157
rect 4160 24191 4212 24200
rect 4160 24157 4169 24191
rect 4169 24157 4203 24191
rect 4203 24157 4212 24191
rect 4620 24191 4672 24200
rect 4160 24148 4212 24157
rect 4620 24157 4629 24191
rect 4629 24157 4663 24191
rect 4663 24157 4672 24191
rect 4620 24148 4672 24157
rect 19708 24216 19760 24268
rect 8944 24191 8996 24200
rect 8944 24157 8953 24191
rect 8953 24157 8987 24191
rect 8987 24157 8996 24191
rect 8944 24148 8996 24157
rect 9220 24191 9272 24200
rect 9220 24157 9229 24191
rect 9229 24157 9263 24191
rect 9263 24157 9272 24191
rect 9220 24148 9272 24157
rect 19524 24148 19576 24200
rect 20996 24216 21048 24268
rect 28540 24216 28592 24268
rect 31300 24216 31352 24268
rect 28632 24191 28684 24200
rect 28632 24157 28641 24191
rect 28641 24157 28675 24191
rect 28675 24157 28684 24191
rect 28632 24148 28684 24157
rect 32864 24191 32916 24200
rect 28540 24080 28592 24132
rect 32864 24157 32873 24191
rect 32873 24157 32907 24191
rect 32907 24157 32916 24191
rect 32864 24148 32916 24157
rect 33140 24191 33192 24200
rect 33140 24157 33149 24191
rect 33149 24157 33183 24191
rect 33183 24157 33192 24191
rect 33140 24148 33192 24157
rect 33876 24148 33928 24200
rect 3608 24012 3660 24064
rect 20628 24012 20680 24064
rect 28816 24055 28868 24064
rect 28816 24021 28825 24055
rect 28825 24021 28859 24055
rect 28859 24021 28868 24055
rect 28816 24012 28868 24021
rect 30564 24012 30616 24064
rect 31208 24055 31260 24064
rect 31208 24021 31217 24055
rect 31217 24021 31251 24055
rect 31251 24021 31260 24055
rect 31208 24012 31260 24021
rect 10398 23910 10450 23962
rect 10462 23910 10514 23962
rect 10526 23910 10578 23962
rect 10590 23910 10642 23962
rect 10654 23910 10706 23962
rect 19846 23910 19898 23962
rect 19910 23910 19962 23962
rect 19974 23910 20026 23962
rect 20038 23910 20090 23962
rect 20102 23910 20154 23962
rect 29294 23910 29346 23962
rect 29358 23910 29410 23962
rect 29422 23910 29474 23962
rect 29486 23910 29538 23962
rect 29550 23910 29602 23962
rect 8024 23851 8076 23860
rect 8024 23817 8033 23851
rect 8033 23817 8067 23851
rect 8067 23817 8076 23851
rect 8024 23808 8076 23817
rect 8392 23808 8444 23860
rect 25872 23808 25924 23860
rect 28540 23808 28592 23860
rect 28724 23851 28776 23860
rect 28724 23817 28733 23851
rect 28733 23817 28767 23851
rect 28767 23817 28776 23851
rect 28724 23808 28776 23817
rect 32956 23851 33008 23860
rect 1860 23672 1912 23724
rect 3608 23715 3660 23724
rect 3608 23681 3617 23715
rect 3617 23681 3651 23715
rect 3651 23681 3660 23715
rect 3608 23672 3660 23681
rect 9496 23740 9548 23792
rect 13544 23740 13596 23792
rect 32956 23817 32965 23851
rect 32965 23817 32999 23851
rect 32999 23817 33008 23851
rect 32956 23808 33008 23817
rect 33876 23808 33928 23860
rect 36728 23808 36780 23860
rect 9864 23672 9916 23724
rect 13268 23715 13320 23724
rect 13268 23681 13277 23715
rect 13277 23681 13311 23715
rect 13311 23681 13320 23715
rect 13268 23672 13320 23681
rect 13912 23672 13964 23724
rect 16856 23715 16908 23724
rect 16856 23681 16865 23715
rect 16865 23681 16899 23715
rect 16899 23681 16908 23715
rect 16856 23672 16908 23681
rect 20628 23715 20680 23724
rect 20628 23681 20637 23715
rect 20637 23681 20671 23715
rect 20671 23681 20680 23715
rect 20628 23672 20680 23681
rect 20904 23715 20956 23724
rect 20904 23681 20913 23715
rect 20913 23681 20947 23715
rect 20947 23681 20956 23715
rect 20904 23672 20956 23681
rect 21732 23672 21784 23724
rect 33784 23740 33836 23792
rect 28816 23672 28868 23724
rect 31300 23715 31352 23724
rect 31300 23681 31309 23715
rect 31309 23681 31343 23715
rect 31343 23681 31352 23715
rect 31300 23672 31352 23681
rect 31852 23672 31904 23724
rect 35900 23715 35952 23724
rect 35900 23681 35909 23715
rect 35909 23681 35943 23715
rect 35943 23681 35952 23715
rect 36728 23715 36780 23724
rect 35900 23672 35952 23681
rect 36728 23681 36737 23715
rect 36737 23681 36771 23715
rect 36771 23681 36780 23715
rect 36728 23672 36780 23681
rect 9496 23647 9548 23656
rect 9496 23613 9505 23647
rect 9505 23613 9539 23647
rect 9539 23613 9548 23647
rect 27712 23647 27764 23656
rect 9496 23604 9548 23613
rect 27712 23613 27721 23647
rect 27721 23613 27755 23647
rect 27755 23613 27764 23647
rect 27712 23604 27764 23613
rect 32036 23604 32088 23656
rect 1492 23511 1544 23520
rect 1492 23477 1501 23511
rect 1501 23477 1535 23511
rect 1535 23477 1544 23511
rect 1492 23468 1544 23477
rect 2872 23511 2924 23520
rect 2872 23477 2881 23511
rect 2881 23477 2915 23511
rect 2915 23477 2924 23511
rect 2872 23468 2924 23477
rect 9956 23511 10008 23520
rect 9956 23477 9965 23511
rect 9965 23477 9999 23511
rect 9999 23477 10008 23511
rect 9956 23468 10008 23477
rect 12256 23468 12308 23520
rect 13912 23511 13964 23520
rect 13912 23477 13921 23511
rect 13921 23477 13955 23511
rect 13955 23477 13964 23511
rect 13912 23468 13964 23477
rect 16672 23511 16724 23520
rect 16672 23477 16681 23511
rect 16681 23477 16715 23511
rect 16715 23477 16724 23511
rect 16672 23468 16724 23477
rect 20996 23468 21048 23520
rect 22836 23468 22888 23520
rect 31300 23468 31352 23520
rect 34612 23647 34664 23656
rect 34612 23613 34621 23647
rect 34621 23613 34655 23647
rect 34655 23613 34664 23647
rect 34612 23604 34664 23613
rect 35532 23468 35584 23520
rect 5674 23366 5726 23418
rect 5738 23366 5790 23418
rect 5802 23366 5854 23418
rect 5866 23366 5918 23418
rect 5930 23366 5982 23418
rect 15122 23366 15174 23418
rect 15186 23366 15238 23418
rect 15250 23366 15302 23418
rect 15314 23366 15366 23418
rect 15378 23366 15430 23418
rect 24570 23366 24622 23418
rect 24634 23366 24686 23418
rect 24698 23366 24750 23418
rect 24762 23366 24814 23418
rect 24826 23366 24878 23418
rect 34018 23366 34070 23418
rect 34082 23366 34134 23418
rect 34146 23366 34198 23418
rect 34210 23366 34262 23418
rect 34274 23366 34326 23418
rect 9864 23307 9916 23316
rect 9864 23273 9873 23307
rect 9873 23273 9907 23307
rect 9907 23273 9916 23307
rect 9864 23264 9916 23273
rect 15568 23264 15620 23316
rect 35900 23264 35952 23316
rect 6920 23128 6972 23180
rect 8944 23128 8996 23180
rect 5448 23060 5500 23112
rect 9036 23103 9088 23112
rect 9036 23069 9045 23103
rect 9045 23069 9079 23103
rect 9079 23069 9088 23103
rect 9036 23060 9088 23069
rect 9588 23128 9640 23180
rect 31852 23128 31904 23180
rect 11704 23060 11756 23112
rect 16672 23060 16724 23112
rect 30932 23103 30984 23112
rect 30932 23069 30941 23103
rect 30941 23069 30975 23103
rect 30975 23069 30984 23103
rect 30932 23060 30984 23069
rect 35532 23103 35584 23112
rect 35532 23069 35541 23103
rect 35541 23069 35575 23103
rect 35575 23069 35584 23103
rect 35532 23060 35584 23069
rect 9956 22992 10008 23044
rect 6000 22924 6052 22976
rect 17040 22967 17092 22976
rect 17040 22933 17049 22967
rect 17049 22933 17083 22967
rect 17083 22933 17092 22967
rect 17040 22924 17092 22933
rect 10398 22822 10450 22874
rect 10462 22822 10514 22874
rect 10526 22822 10578 22874
rect 10590 22822 10642 22874
rect 10654 22822 10706 22874
rect 19846 22822 19898 22874
rect 19910 22822 19962 22874
rect 19974 22822 20026 22874
rect 20038 22822 20090 22874
rect 20102 22822 20154 22874
rect 29294 22822 29346 22874
rect 29358 22822 29410 22874
rect 29422 22822 29474 22874
rect 29486 22822 29538 22874
rect 29550 22822 29602 22874
rect 3884 22763 3936 22772
rect 3884 22729 3893 22763
rect 3893 22729 3927 22763
rect 3927 22729 3936 22763
rect 3884 22720 3936 22729
rect 9496 22720 9548 22772
rect 16856 22720 16908 22772
rect 4620 22584 4672 22636
rect 5448 22584 5500 22636
rect 10140 22627 10192 22636
rect 10140 22593 10149 22627
rect 10149 22593 10183 22627
rect 10183 22593 10192 22627
rect 10140 22584 10192 22593
rect 14740 22584 14792 22636
rect 15016 22584 15068 22636
rect 20812 22584 20864 22636
rect 25688 22627 25740 22636
rect 25688 22593 25697 22627
rect 25697 22593 25731 22627
rect 25731 22593 25740 22627
rect 25688 22584 25740 22593
rect 7380 22516 7432 22568
rect 13820 22516 13872 22568
rect 3884 22448 3936 22500
rect 13544 22448 13596 22500
rect 1400 22423 1452 22432
rect 1400 22389 1409 22423
rect 1409 22389 1443 22423
rect 1443 22389 1452 22423
rect 1400 22380 1452 22389
rect 3056 22380 3108 22432
rect 6920 22380 6972 22432
rect 12992 22380 13044 22432
rect 26240 22380 26292 22432
rect 5674 22278 5726 22330
rect 5738 22278 5790 22330
rect 5802 22278 5854 22330
rect 5866 22278 5918 22330
rect 5930 22278 5982 22330
rect 15122 22278 15174 22330
rect 15186 22278 15238 22330
rect 15250 22278 15302 22330
rect 15314 22278 15366 22330
rect 15378 22278 15430 22330
rect 24570 22278 24622 22330
rect 24634 22278 24686 22330
rect 24698 22278 24750 22330
rect 24762 22278 24814 22330
rect 24826 22278 24878 22330
rect 34018 22278 34070 22330
rect 34082 22278 34134 22330
rect 34146 22278 34198 22330
rect 34210 22278 34262 22330
rect 34274 22278 34326 22330
rect 10140 22176 10192 22228
rect 11704 22176 11756 22228
rect 14740 22083 14792 22092
rect 14740 22049 14749 22083
rect 14749 22049 14783 22083
rect 14783 22049 14792 22083
rect 14740 22040 14792 22049
rect 23480 22040 23532 22092
rect 24400 22083 24452 22092
rect 24400 22049 24409 22083
rect 24409 22049 24443 22083
rect 24443 22049 24452 22083
rect 24400 22040 24452 22049
rect 6000 21972 6052 22024
rect 6920 22015 6972 22024
rect 6920 21981 6929 22015
rect 6929 21981 6963 22015
rect 6963 21981 6972 22015
rect 6920 21972 6972 21981
rect 10048 21972 10100 22024
rect 12992 22015 13044 22024
rect 12992 21981 13001 22015
rect 13001 21981 13035 22015
rect 13035 21981 13044 22015
rect 12992 21972 13044 21981
rect 23664 22015 23716 22024
rect 12072 21904 12124 21956
rect 14832 21904 14884 21956
rect 23664 21981 23673 22015
rect 23673 21981 23707 22015
rect 23707 21981 23716 22015
rect 23664 21972 23716 21981
rect 6000 21879 6052 21888
rect 6000 21845 6009 21879
rect 6009 21845 6043 21879
rect 6043 21845 6052 21879
rect 6000 21836 6052 21845
rect 7012 21836 7064 21888
rect 12164 21836 12216 21888
rect 12348 21836 12400 21888
rect 25872 21972 25924 22024
rect 26240 22015 26292 22024
rect 26240 21981 26249 22015
rect 26249 21981 26283 22015
rect 26283 21981 26292 22015
rect 26240 21972 26292 21981
rect 27068 22015 27120 22024
rect 27068 21981 27077 22015
rect 27077 21981 27111 22015
rect 27111 21981 27120 22015
rect 27068 21972 27120 21981
rect 33876 21972 33928 22024
rect 25412 21879 25464 21888
rect 25412 21845 25421 21879
rect 25421 21845 25455 21879
rect 25455 21845 25464 21879
rect 25412 21836 25464 21845
rect 10398 21734 10450 21786
rect 10462 21734 10514 21786
rect 10526 21734 10578 21786
rect 10590 21734 10642 21786
rect 10654 21734 10706 21786
rect 19846 21734 19898 21786
rect 19910 21734 19962 21786
rect 19974 21734 20026 21786
rect 20038 21734 20090 21786
rect 20102 21734 20154 21786
rect 29294 21734 29346 21786
rect 29358 21734 29410 21786
rect 29422 21734 29474 21786
rect 29486 21734 29538 21786
rect 29550 21734 29602 21786
rect 19340 21632 19392 21684
rect 23480 21632 23532 21684
rect 23664 21675 23716 21684
rect 23664 21641 23673 21675
rect 23673 21641 23707 21675
rect 23707 21641 23716 21675
rect 23664 21632 23716 21641
rect 25688 21632 25740 21684
rect 3056 21539 3108 21548
rect 3056 21505 3065 21539
rect 3065 21505 3099 21539
rect 3099 21505 3108 21539
rect 3056 21496 3108 21505
rect 18788 21539 18840 21548
rect 18788 21505 18797 21539
rect 18797 21505 18831 21539
rect 18831 21505 18840 21539
rect 18788 21496 18840 21505
rect 19248 21496 19300 21548
rect 19708 21496 19760 21548
rect 20352 21496 20404 21548
rect 23480 21539 23532 21548
rect 23480 21505 23489 21539
rect 23489 21505 23523 21539
rect 23523 21505 23532 21539
rect 23480 21496 23532 21505
rect 25136 21539 25188 21548
rect 25136 21505 25145 21539
rect 25145 21505 25179 21539
rect 25179 21505 25188 21539
rect 25136 21496 25188 21505
rect 30932 21496 30984 21548
rect 34520 21539 34572 21548
rect 34520 21505 34529 21539
rect 34529 21505 34563 21539
rect 34563 21505 34572 21539
rect 34520 21496 34572 21505
rect 23388 21428 23440 21480
rect 34428 21428 34480 21480
rect 2964 21292 3016 21344
rect 20260 21292 20312 21344
rect 35992 21292 36044 21344
rect 5674 21190 5726 21242
rect 5738 21190 5790 21242
rect 5802 21190 5854 21242
rect 5866 21190 5918 21242
rect 5930 21190 5982 21242
rect 15122 21190 15174 21242
rect 15186 21190 15238 21242
rect 15250 21190 15302 21242
rect 15314 21190 15366 21242
rect 15378 21190 15430 21242
rect 24570 21190 24622 21242
rect 24634 21190 24686 21242
rect 24698 21190 24750 21242
rect 24762 21190 24814 21242
rect 24826 21190 24878 21242
rect 34018 21190 34070 21242
rect 34082 21190 34134 21242
rect 34146 21190 34198 21242
rect 34210 21190 34262 21242
rect 34274 21190 34326 21242
rect 1768 20884 1820 20936
rect 2964 20927 3016 20936
rect 2964 20893 2973 20927
rect 2973 20893 3007 20927
rect 3007 20893 3016 20927
rect 2964 20884 3016 20893
rect 3884 20884 3936 20936
rect 6000 20927 6052 20936
rect 6000 20893 6009 20927
rect 6009 20893 6043 20927
rect 6043 20893 6052 20927
rect 6000 20884 6052 20893
rect 6644 20884 6696 20936
rect 7012 20927 7064 20936
rect 7012 20893 7021 20927
rect 7021 20893 7055 20927
rect 7055 20893 7064 20927
rect 7012 20884 7064 20893
rect 20904 21088 20956 21140
rect 20260 20927 20312 20936
rect 20260 20893 20269 20927
rect 20269 20893 20303 20927
rect 20303 20893 20312 20927
rect 20260 20884 20312 20893
rect 29736 20927 29788 20936
rect 29736 20893 29745 20927
rect 29745 20893 29779 20927
rect 29779 20893 29788 20927
rect 29736 20884 29788 20893
rect 30472 20884 30524 20936
rect 35992 20927 36044 20936
rect 35992 20893 36001 20927
rect 36001 20893 36035 20927
rect 36035 20893 36044 20927
rect 35992 20884 36044 20893
rect 25412 20816 25464 20868
rect 1492 20791 1544 20800
rect 1492 20757 1501 20791
rect 1501 20757 1535 20791
rect 1535 20757 1544 20791
rect 1492 20748 1544 20757
rect 2228 20791 2280 20800
rect 2228 20757 2237 20791
rect 2237 20757 2271 20791
rect 2271 20757 2280 20791
rect 2228 20748 2280 20757
rect 6736 20748 6788 20800
rect 19248 20791 19300 20800
rect 19248 20757 19257 20791
rect 19257 20757 19291 20791
rect 19291 20757 19300 20791
rect 19248 20748 19300 20757
rect 20996 20791 21048 20800
rect 20996 20757 21005 20791
rect 21005 20757 21039 20791
rect 21039 20757 21048 20791
rect 20996 20748 21048 20757
rect 29920 20791 29972 20800
rect 29920 20757 29929 20791
rect 29929 20757 29963 20791
rect 29963 20757 29972 20791
rect 29920 20748 29972 20757
rect 30380 20791 30432 20800
rect 30380 20757 30389 20791
rect 30389 20757 30423 20791
rect 30423 20757 30432 20791
rect 30380 20748 30432 20757
rect 36912 20748 36964 20800
rect 10398 20646 10450 20698
rect 10462 20646 10514 20698
rect 10526 20646 10578 20698
rect 10590 20646 10642 20698
rect 10654 20646 10706 20698
rect 19846 20646 19898 20698
rect 19910 20646 19962 20698
rect 19974 20646 20026 20698
rect 20038 20646 20090 20698
rect 20102 20646 20154 20698
rect 29294 20646 29346 20698
rect 29358 20646 29410 20698
rect 29422 20646 29474 20698
rect 29486 20646 29538 20698
rect 29550 20646 29602 20698
rect 1768 20587 1820 20596
rect 1768 20553 1777 20587
rect 1777 20553 1811 20587
rect 1811 20553 1820 20587
rect 1768 20544 1820 20553
rect 2780 20544 2832 20596
rect 19708 20544 19760 20596
rect 29736 20544 29788 20596
rect 19248 20476 19300 20528
rect 22928 20476 22980 20528
rect 19616 20451 19668 20460
rect 19616 20417 19625 20451
rect 19625 20417 19659 20451
rect 19659 20417 19668 20451
rect 19616 20408 19668 20417
rect 27528 20408 27580 20460
rect 31300 20408 31352 20460
rect 33232 20408 33284 20460
rect 34336 20408 34388 20460
rect 17224 20383 17276 20392
rect 17224 20349 17233 20383
rect 17233 20349 17267 20383
rect 17267 20349 17276 20383
rect 17224 20340 17276 20349
rect 23388 20340 23440 20392
rect 30472 20340 30524 20392
rect 31208 20272 31260 20324
rect 9588 20247 9640 20256
rect 9588 20213 9597 20247
rect 9597 20213 9631 20247
rect 9631 20213 9640 20247
rect 9588 20204 9640 20213
rect 33876 20204 33928 20256
rect 35992 20204 36044 20256
rect 5674 20102 5726 20154
rect 5738 20102 5790 20154
rect 5802 20102 5854 20154
rect 5866 20102 5918 20154
rect 5930 20102 5982 20154
rect 15122 20102 15174 20154
rect 15186 20102 15238 20154
rect 15250 20102 15302 20154
rect 15314 20102 15366 20154
rect 15378 20102 15430 20154
rect 24570 20102 24622 20154
rect 24634 20102 24686 20154
rect 24698 20102 24750 20154
rect 24762 20102 24814 20154
rect 24826 20102 24878 20154
rect 34018 20102 34070 20154
rect 34082 20102 34134 20154
rect 34146 20102 34198 20154
rect 34210 20102 34262 20154
rect 34274 20102 34326 20154
rect 6644 20043 6696 20052
rect 6644 20009 6653 20043
rect 6653 20009 6687 20043
rect 6687 20009 6696 20043
rect 6644 20000 6696 20009
rect 14832 20043 14884 20052
rect 14832 20009 14841 20043
rect 14841 20009 14875 20043
rect 14875 20009 14884 20043
rect 14832 20000 14884 20009
rect 17040 20000 17092 20052
rect 15568 19864 15620 19916
rect 6276 19796 6328 19848
rect 9680 19796 9732 19848
rect 20536 19864 20588 19916
rect 17040 19796 17092 19848
rect 11704 19728 11756 19780
rect 14556 19728 14608 19780
rect 1492 19703 1544 19712
rect 1492 19669 1501 19703
rect 1501 19669 1535 19703
rect 1535 19669 1544 19703
rect 1492 19660 1544 19669
rect 20352 19728 20404 19780
rect 28908 19796 28960 19848
rect 29920 19839 29972 19848
rect 29920 19805 29929 19839
rect 29929 19805 29963 19839
rect 29963 19805 29972 19839
rect 29920 19796 29972 19805
rect 33876 19839 33928 19848
rect 33876 19805 33885 19839
rect 33885 19805 33919 19839
rect 33919 19805 33928 19839
rect 33876 19796 33928 19805
rect 35992 19839 36044 19848
rect 35992 19805 36001 19839
rect 36001 19805 36035 19839
rect 36035 19805 36044 19839
rect 35992 19796 36044 19805
rect 25044 19728 25096 19780
rect 27528 19728 27580 19780
rect 35900 19728 35952 19780
rect 22008 19660 22060 19712
rect 30472 19660 30524 19712
rect 34704 19660 34756 19712
rect 37464 19660 37516 19712
rect 10398 19558 10450 19610
rect 10462 19558 10514 19610
rect 10526 19558 10578 19610
rect 10590 19558 10642 19610
rect 10654 19558 10706 19610
rect 19846 19558 19898 19610
rect 19910 19558 19962 19610
rect 19974 19558 20026 19610
rect 20038 19558 20090 19610
rect 20102 19558 20154 19610
rect 29294 19558 29346 19610
rect 29358 19558 29410 19610
rect 29422 19558 29474 19610
rect 29486 19558 29538 19610
rect 29550 19558 29602 19610
rect 11704 19456 11756 19508
rect 17040 19499 17092 19508
rect 4620 19320 4672 19372
rect 7104 19363 7156 19372
rect 7104 19329 7113 19363
rect 7113 19329 7147 19363
rect 7147 19329 7156 19363
rect 7104 19320 7156 19329
rect 9404 19320 9456 19372
rect 17040 19465 17049 19499
rect 17049 19465 17083 19499
rect 17083 19465 17092 19499
rect 17040 19456 17092 19465
rect 28908 19456 28960 19508
rect 30472 19456 30524 19508
rect 37464 19456 37516 19508
rect 11336 19320 11388 19372
rect 14832 19320 14884 19372
rect 22008 19363 22060 19372
rect 22008 19329 22017 19363
rect 22017 19329 22051 19363
rect 22051 19329 22060 19363
rect 22008 19320 22060 19329
rect 25964 19363 26016 19372
rect 4160 19252 4212 19304
rect 17224 19252 17276 19304
rect 25964 19329 25973 19363
rect 25973 19329 26007 19363
rect 26007 19329 26016 19363
rect 25964 19320 26016 19329
rect 28908 19320 28960 19372
rect 30380 19320 30432 19372
rect 34704 19363 34756 19372
rect 34704 19329 34713 19363
rect 34713 19329 34747 19363
rect 34747 19329 34756 19363
rect 34704 19320 34756 19329
rect 35900 19320 35952 19372
rect 36636 19320 36688 19372
rect 26240 19184 26292 19236
rect 3976 19116 4028 19168
rect 7012 19116 7064 19168
rect 21640 19116 21692 19168
rect 5674 19014 5726 19066
rect 5738 19014 5790 19066
rect 5802 19014 5854 19066
rect 5866 19014 5918 19066
rect 5930 19014 5982 19066
rect 15122 19014 15174 19066
rect 15186 19014 15238 19066
rect 15250 19014 15302 19066
rect 15314 19014 15366 19066
rect 15378 19014 15430 19066
rect 24570 19014 24622 19066
rect 24634 19014 24686 19066
rect 24698 19014 24750 19066
rect 24762 19014 24814 19066
rect 24826 19014 24878 19066
rect 34018 19014 34070 19066
rect 34082 19014 34134 19066
rect 34146 19014 34198 19066
rect 34210 19014 34262 19066
rect 34274 19014 34326 19066
rect 6736 18912 6788 18964
rect 10048 18955 10100 18964
rect 10048 18921 10057 18955
rect 10057 18921 10091 18955
rect 10091 18921 10100 18955
rect 10048 18912 10100 18921
rect 20904 18955 20956 18964
rect 20904 18921 20913 18955
rect 20913 18921 20947 18955
rect 20947 18921 20956 18955
rect 20904 18912 20956 18921
rect 29828 18912 29880 18964
rect 30472 18912 30524 18964
rect 9496 18776 9548 18828
rect 23388 18776 23440 18828
rect 3976 18751 4028 18760
rect 3976 18717 3985 18751
rect 3985 18717 4019 18751
rect 4019 18717 4028 18751
rect 3976 18708 4028 18717
rect 6276 18708 6328 18760
rect 7012 18708 7064 18760
rect 9864 18751 9916 18760
rect 9864 18717 9873 18751
rect 9873 18717 9907 18751
rect 9907 18717 9916 18751
rect 9864 18708 9916 18717
rect 21640 18751 21692 18760
rect 21640 18717 21649 18751
rect 21649 18717 21683 18751
rect 21683 18717 21692 18751
rect 21640 18708 21692 18717
rect 11152 18640 11204 18692
rect 11336 18640 11388 18692
rect 20628 18640 20680 18692
rect 24492 18708 24544 18760
rect 25412 18708 25464 18760
rect 36636 18751 36688 18760
rect 36636 18717 36645 18751
rect 36645 18717 36679 18751
rect 36679 18717 36688 18751
rect 36636 18708 36688 18717
rect 36912 18751 36964 18760
rect 36912 18717 36921 18751
rect 36921 18717 36955 18751
rect 36955 18717 36964 18751
rect 36912 18708 36964 18717
rect 25964 18640 26016 18692
rect 3608 18572 3660 18624
rect 12256 18572 12308 18624
rect 25228 18572 25280 18624
rect 37464 18572 37516 18624
rect 10398 18470 10450 18522
rect 10462 18470 10514 18522
rect 10526 18470 10578 18522
rect 10590 18470 10642 18522
rect 10654 18470 10706 18522
rect 19846 18470 19898 18522
rect 19910 18470 19962 18522
rect 19974 18470 20026 18522
rect 20038 18470 20090 18522
rect 20102 18470 20154 18522
rect 29294 18470 29346 18522
rect 29358 18470 29410 18522
rect 29422 18470 29474 18522
rect 29486 18470 29538 18522
rect 29550 18470 29602 18522
rect 7104 18368 7156 18420
rect 12900 18368 12952 18420
rect 25412 18411 25464 18420
rect 25412 18377 25421 18411
rect 25421 18377 25455 18411
rect 25455 18377 25464 18411
rect 25412 18368 25464 18377
rect 8300 18300 8352 18352
rect 9588 18300 9640 18352
rect 11152 18300 11204 18352
rect 1952 18232 2004 18284
rect 3608 18275 3660 18284
rect 3608 18241 3617 18275
rect 3617 18241 3651 18275
rect 3651 18241 3660 18275
rect 3608 18232 3660 18241
rect 3884 18275 3936 18284
rect 3884 18241 3893 18275
rect 3893 18241 3927 18275
rect 3927 18241 3936 18275
rect 3884 18232 3936 18241
rect 4620 18164 4672 18216
rect 14372 18275 14424 18284
rect 14372 18241 14381 18275
rect 14381 18241 14415 18275
rect 14415 18241 14424 18275
rect 14372 18232 14424 18241
rect 14556 18275 14608 18284
rect 14556 18241 14565 18275
rect 14565 18241 14599 18275
rect 14599 18241 14608 18275
rect 25228 18275 25280 18284
rect 14556 18232 14608 18241
rect 25228 18241 25237 18275
rect 25237 18241 25271 18275
rect 25271 18241 25280 18275
rect 25228 18232 25280 18241
rect 7288 18207 7340 18216
rect 7288 18173 7297 18207
rect 7297 18173 7331 18207
rect 7331 18173 7340 18207
rect 7288 18164 7340 18173
rect 9128 18164 9180 18216
rect 10876 18164 10928 18216
rect 12900 18164 12952 18216
rect 13268 18164 13320 18216
rect 1492 18071 1544 18080
rect 1492 18037 1501 18071
rect 1501 18037 1535 18071
rect 1535 18037 1544 18071
rect 1492 18028 1544 18037
rect 1952 18028 2004 18080
rect 2228 18028 2280 18080
rect 14280 18071 14332 18080
rect 14280 18037 14289 18071
rect 14289 18037 14323 18071
rect 14323 18037 14332 18071
rect 14280 18028 14332 18037
rect 5674 17926 5726 17978
rect 5738 17926 5790 17978
rect 5802 17926 5854 17978
rect 5866 17926 5918 17978
rect 5930 17926 5982 17978
rect 15122 17926 15174 17978
rect 15186 17926 15238 17978
rect 15250 17926 15302 17978
rect 15314 17926 15366 17978
rect 15378 17926 15430 17978
rect 24570 17926 24622 17978
rect 24634 17926 24686 17978
rect 24698 17926 24750 17978
rect 24762 17926 24814 17978
rect 24826 17926 24878 17978
rect 34018 17926 34070 17978
rect 34082 17926 34134 17978
rect 34146 17926 34198 17978
rect 34210 17926 34262 17978
rect 34274 17926 34326 17978
rect 9864 17824 9916 17876
rect 14280 17824 14332 17876
rect 4620 17731 4672 17740
rect 4620 17697 4629 17731
rect 4629 17697 4663 17731
rect 4663 17697 4672 17731
rect 4620 17688 4672 17697
rect 3976 17552 4028 17604
rect 8208 17620 8260 17672
rect 14372 17620 14424 17672
rect 14740 17663 14792 17672
rect 14740 17629 14749 17663
rect 14749 17629 14783 17663
rect 14783 17629 14792 17663
rect 14740 17620 14792 17629
rect 15476 17620 15528 17672
rect 23572 17620 23624 17672
rect 24492 17620 24544 17672
rect 25044 17620 25096 17672
rect 26332 17620 26384 17672
rect 26976 17663 27028 17672
rect 26976 17629 26985 17663
rect 26985 17629 27019 17663
rect 27019 17629 27028 17663
rect 26976 17620 27028 17629
rect 10968 17552 11020 17604
rect 17960 17552 18012 17604
rect 19432 17552 19484 17604
rect 7288 17484 7340 17536
rect 8852 17484 8904 17536
rect 17776 17484 17828 17536
rect 22100 17484 22152 17536
rect 29092 17484 29144 17536
rect 10398 17382 10450 17434
rect 10462 17382 10514 17434
rect 10526 17382 10578 17434
rect 10590 17382 10642 17434
rect 10654 17382 10706 17434
rect 19846 17382 19898 17434
rect 19910 17382 19962 17434
rect 19974 17382 20026 17434
rect 20038 17382 20090 17434
rect 20102 17382 20154 17434
rect 29294 17382 29346 17434
rect 29358 17382 29410 17434
rect 29422 17382 29474 17434
rect 29486 17382 29538 17434
rect 29550 17382 29602 17434
rect 13452 17280 13504 17332
rect 17776 17323 17828 17332
rect 17776 17289 17785 17323
rect 17785 17289 17819 17323
rect 17819 17289 17828 17323
rect 17776 17280 17828 17289
rect 19616 17280 19668 17332
rect 25136 17280 25188 17332
rect 26976 17280 27028 17332
rect 30656 17280 30708 17332
rect 17960 17144 18012 17196
rect 19064 17144 19116 17196
rect 19800 17212 19852 17264
rect 22100 17255 22152 17264
rect 22100 17221 22109 17255
rect 22109 17221 22143 17255
rect 22143 17221 22152 17255
rect 22100 17212 22152 17221
rect 22284 17255 22336 17264
rect 22284 17221 22309 17255
rect 22309 17221 22336 17255
rect 22284 17212 22336 17221
rect 28908 17212 28960 17264
rect 29092 17187 29144 17196
rect 29092 17153 29101 17187
rect 29101 17153 29135 17187
rect 29135 17153 29144 17187
rect 29092 17144 29144 17153
rect 33232 17187 33284 17196
rect 33232 17153 33241 17187
rect 33241 17153 33275 17187
rect 33275 17153 33284 17187
rect 33232 17144 33284 17153
rect 35072 17144 35124 17196
rect 29828 17051 29880 17060
rect 29828 17017 29837 17051
rect 29837 17017 29871 17051
rect 29871 17017 29880 17051
rect 29828 17008 29880 17017
rect 30748 17008 30800 17060
rect 1492 16983 1544 16992
rect 1492 16949 1501 16983
rect 1501 16949 1535 16983
rect 1535 16949 1544 16983
rect 1492 16940 1544 16949
rect 17776 16983 17828 16992
rect 17776 16949 17785 16983
rect 17785 16949 17819 16983
rect 17819 16949 17828 16983
rect 17776 16940 17828 16949
rect 18788 16983 18840 16992
rect 18788 16949 18797 16983
rect 18797 16949 18831 16983
rect 18831 16949 18840 16983
rect 18788 16940 18840 16949
rect 21456 16940 21508 16992
rect 33416 16983 33468 16992
rect 33416 16949 33425 16983
rect 33425 16949 33459 16983
rect 33459 16949 33468 16983
rect 33416 16940 33468 16949
rect 36728 16940 36780 16992
rect 5674 16838 5726 16890
rect 5738 16838 5790 16890
rect 5802 16838 5854 16890
rect 5866 16838 5918 16890
rect 5930 16838 5982 16890
rect 15122 16838 15174 16890
rect 15186 16838 15238 16890
rect 15250 16838 15302 16890
rect 15314 16838 15366 16890
rect 15378 16838 15430 16890
rect 24570 16838 24622 16890
rect 24634 16838 24686 16890
rect 24698 16838 24750 16890
rect 24762 16838 24814 16890
rect 24826 16838 24878 16890
rect 34018 16838 34070 16890
rect 34082 16838 34134 16890
rect 34146 16838 34198 16890
rect 34210 16838 34262 16890
rect 34274 16838 34326 16890
rect 4160 16736 4212 16788
rect 9036 16736 9088 16788
rect 9680 16736 9732 16788
rect 23480 16736 23532 16788
rect 35072 16779 35124 16788
rect 35072 16745 35081 16779
rect 35081 16745 35115 16779
rect 35115 16745 35124 16779
rect 35072 16736 35124 16745
rect 1584 16668 1636 16720
rect 2228 16711 2280 16720
rect 2228 16677 2237 16711
rect 2237 16677 2271 16711
rect 2271 16677 2280 16711
rect 2228 16668 2280 16677
rect 2964 16575 3016 16584
rect 2964 16541 2973 16575
rect 2973 16541 3007 16575
rect 3007 16541 3016 16575
rect 2964 16532 3016 16541
rect 3976 16575 4028 16584
rect 3976 16541 3985 16575
rect 3985 16541 4019 16575
rect 4019 16541 4028 16575
rect 3976 16532 4028 16541
rect 4160 16575 4212 16584
rect 4160 16541 4169 16575
rect 4169 16541 4203 16575
rect 4203 16541 4212 16575
rect 4160 16532 4212 16541
rect 9404 16668 9456 16720
rect 9956 16668 10008 16720
rect 16120 16711 16172 16720
rect 16120 16677 16129 16711
rect 16129 16677 16163 16711
rect 16163 16677 16172 16711
rect 16120 16668 16172 16677
rect 6920 16600 6972 16652
rect 8208 16600 8260 16652
rect 11704 16600 11756 16652
rect 12072 16643 12124 16652
rect 12072 16609 12081 16643
rect 12081 16609 12115 16643
rect 12115 16609 12124 16643
rect 12072 16600 12124 16609
rect 19800 16643 19852 16652
rect 19800 16609 19809 16643
rect 19809 16609 19843 16643
rect 19843 16609 19852 16643
rect 19800 16600 19852 16609
rect 22284 16668 22336 16720
rect 21088 16643 21140 16652
rect 21088 16609 21097 16643
rect 21097 16609 21131 16643
rect 21131 16609 21140 16643
rect 21088 16600 21140 16609
rect 22836 16643 22888 16652
rect 22836 16609 22845 16643
rect 22845 16609 22879 16643
rect 22879 16609 22888 16643
rect 22836 16600 22888 16609
rect 37464 16668 37516 16720
rect 23480 16600 23532 16652
rect 33232 16600 33284 16652
rect 6276 16532 6328 16584
rect 9588 16532 9640 16584
rect 9956 16532 10008 16584
rect 10784 16532 10836 16584
rect 14556 16532 14608 16584
rect 6920 16464 6972 16516
rect 10968 16464 11020 16516
rect 14372 16464 14424 16516
rect 15844 16507 15896 16516
rect 15844 16473 15853 16507
rect 15853 16473 15887 16507
rect 15887 16473 15896 16507
rect 15844 16464 15896 16473
rect 21180 16464 21232 16516
rect 22100 16464 22152 16516
rect 22284 16464 22336 16516
rect 2780 16396 2832 16448
rect 7104 16439 7156 16448
rect 7104 16405 7113 16439
rect 7113 16405 7147 16439
rect 7147 16405 7156 16439
rect 7104 16396 7156 16405
rect 11336 16439 11388 16448
rect 11336 16405 11345 16439
rect 11345 16405 11379 16439
rect 11379 16405 11388 16439
rect 11336 16396 11388 16405
rect 12348 16439 12400 16448
rect 12348 16405 12357 16439
rect 12357 16405 12391 16439
rect 12391 16405 12400 16439
rect 12348 16396 12400 16405
rect 17776 16396 17828 16448
rect 21456 16439 21508 16448
rect 21456 16405 21465 16439
rect 21465 16405 21499 16439
rect 21499 16405 21508 16439
rect 21456 16396 21508 16405
rect 21824 16396 21876 16448
rect 23572 16532 23624 16584
rect 32128 16532 32180 16584
rect 33416 16532 33468 16584
rect 34612 16532 34664 16584
rect 35716 16575 35768 16584
rect 35716 16541 35725 16575
rect 35725 16541 35759 16575
rect 35759 16541 35768 16575
rect 35716 16532 35768 16541
rect 23664 16464 23716 16516
rect 33232 16396 33284 16448
rect 10398 16294 10450 16346
rect 10462 16294 10514 16346
rect 10526 16294 10578 16346
rect 10590 16294 10642 16346
rect 10654 16294 10706 16346
rect 19846 16294 19898 16346
rect 19910 16294 19962 16346
rect 19974 16294 20026 16346
rect 20038 16294 20090 16346
rect 20102 16294 20154 16346
rect 29294 16294 29346 16346
rect 29358 16294 29410 16346
rect 29422 16294 29474 16346
rect 29486 16294 29538 16346
rect 29550 16294 29602 16346
rect 2964 16235 3016 16244
rect 2964 16201 2973 16235
rect 2973 16201 3007 16235
rect 3007 16201 3016 16235
rect 2964 16192 3016 16201
rect 10784 16192 10836 16244
rect 11704 16192 11756 16244
rect 20628 16192 20680 16244
rect 25872 16235 25924 16244
rect 25872 16201 25881 16235
rect 25881 16201 25915 16235
rect 25915 16201 25924 16235
rect 25872 16192 25924 16201
rect 36452 16192 36504 16244
rect 36636 16192 36688 16244
rect 8300 16124 8352 16176
rect 11060 16124 11112 16176
rect 14832 16124 14884 16176
rect 26240 16124 26292 16176
rect 2780 16099 2832 16108
rect 2780 16065 2789 16099
rect 2789 16065 2823 16099
rect 2823 16065 2832 16099
rect 2780 16056 2832 16065
rect 9404 16056 9456 16108
rect 12348 16056 12400 16108
rect 25136 16056 25188 16108
rect 26332 16099 26384 16108
rect 10140 16031 10192 16040
rect 10140 15997 10149 16031
rect 10149 15997 10183 16031
rect 10183 15997 10192 16031
rect 10140 15988 10192 15997
rect 10324 16031 10376 16040
rect 10324 15997 10333 16031
rect 10333 15997 10367 16031
rect 10367 15997 10376 16031
rect 11704 16031 11756 16040
rect 10324 15988 10376 15997
rect 11704 15997 11713 16031
rect 11713 15997 11747 16031
rect 11747 15997 11756 16031
rect 11704 15988 11756 15997
rect 8852 15920 8904 15972
rect 11336 15920 11388 15972
rect 24492 15988 24544 16040
rect 26332 16065 26341 16099
rect 26341 16065 26375 16099
rect 26375 16065 26384 16099
rect 26332 16056 26384 16065
rect 34520 16056 34572 16108
rect 35716 16099 35768 16108
rect 35716 16065 35725 16099
rect 35725 16065 35759 16099
rect 35759 16065 35768 16099
rect 35716 16056 35768 16065
rect 12256 15963 12308 15972
rect 12256 15929 12265 15963
rect 12265 15929 12299 15963
rect 12299 15929 12308 15963
rect 12256 15920 12308 15929
rect 16120 15920 16172 15972
rect 24308 15920 24360 15972
rect 34612 15920 34664 15972
rect 9036 15852 9088 15904
rect 9496 15852 9548 15904
rect 30196 15852 30248 15904
rect 5674 15750 5726 15802
rect 5738 15750 5790 15802
rect 5802 15750 5854 15802
rect 5866 15750 5918 15802
rect 5930 15750 5982 15802
rect 15122 15750 15174 15802
rect 15186 15750 15238 15802
rect 15250 15750 15302 15802
rect 15314 15750 15366 15802
rect 15378 15750 15430 15802
rect 24570 15750 24622 15802
rect 24634 15750 24686 15802
rect 24698 15750 24750 15802
rect 24762 15750 24814 15802
rect 24826 15750 24878 15802
rect 34018 15750 34070 15802
rect 34082 15750 34134 15802
rect 34146 15750 34198 15802
rect 34210 15750 34262 15802
rect 34274 15750 34326 15802
rect 9680 15648 9732 15700
rect 24952 15648 25004 15700
rect 30748 15691 30800 15700
rect 30748 15657 30757 15691
rect 30757 15657 30791 15691
rect 30791 15657 30800 15691
rect 30748 15648 30800 15657
rect 37464 15691 37516 15700
rect 37464 15657 37473 15691
rect 37473 15657 37507 15691
rect 37507 15657 37516 15691
rect 37464 15648 37516 15657
rect 8392 15580 8444 15632
rect 9404 15580 9456 15632
rect 11704 15580 11756 15632
rect 15844 15580 15896 15632
rect 27068 15580 27120 15632
rect 26240 15512 26292 15564
rect 36452 15555 36504 15564
rect 36452 15521 36461 15555
rect 36461 15521 36495 15555
rect 36495 15521 36504 15555
rect 36452 15512 36504 15521
rect 12256 15444 12308 15496
rect 14372 15487 14424 15496
rect 14372 15453 14381 15487
rect 14381 15453 14415 15487
rect 14415 15453 14424 15487
rect 14372 15444 14424 15453
rect 14556 15487 14608 15496
rect 14556 15453 14565 15487
rect 14565 15453 14599 15487
rect 14599 15453 14608 15487
rect 14556 15444 14608 15453
rect 14832 15487 14884 15496
rect 14832 15453 14841 15487
rect 14841 15453 14875 15487
rect 14875 15453 14884 15487
rect 14832 15444 14884 15453
rect 15752 15444 15804 15496
rect 30012 15487 30064 15496
rect 30012 15453 30021 15487
rect 30021 15453 30055 15487
rect 30055 15453 30064 15487
rect 30012 15444 30064 15453
rect 36728 15487 36780 15496
rect 36728 15453 36737 15487
rect 36737 15453 36771 15487
rect 36771 15453 36780 15487
rect 36728 15444 36780 15453
rect 8852 15376 8904 15428
rect 11060 15376 11112 15428
rect 24492 15376 24544 15428
rect 26056 15376 26108 15428
rect 1492 15351 1544 15360
rect 1492 15317 1501 15351
rect 1501 15317 1535 15351
rect 1535 15317 1544 15351
rect 1492 15308 1544 15317
rect 9680 15351 9732 15360
rect 9680 15317 9689 15351
rect 9689 15317 9723 15351
rect 9723 15317 9732 15351
rect 9680 15308 9732 15317
rect 10398 15206 10450 15258
rect 10462 15206 10514 15258
rect 10526 15206 10578 15258
rect 10590 15206 10642 15258
rect 10654 15206 10706 15258
rect 19846 15206 19898 15258
rect 19910 15206 19962 15258
rect 19974 15206 20026 15258
rect 20038 15206 20090 15258
rect 20102 15206 20154 15258
rect 29294 15206 29346 15258
rect 29358 15206 29410 15258
rect 29422 15206 29474 15258
rect 29486 15206 29538 15258
rect 29550 15206 29602 15258
rect 18788 15147 18840 15156
rect 18788 15113 18797 15147
rect 18797 15113 18831 15147
rect 18831 15113 18840 15147
rect 18788 15104 18840 15113
rect 27712 15104 27764 15156
rect 30012 15147 30064 15156
rect 30012 15113 30021 15147
rect 30021 15113 30055 15147
rect 30055 15113 30064 15147
rect 30012 15104 30064 15113
rect 37464 15104 37516 15156
rect 13820 15036 13872 15088
rect 14556 15036 14608 15088
rect 11060 14968 11112 15020
rect 14832 14968 14884 15020
rect 10140 14943 10192 14952
rect 10140 14909 10149 14943
rect 10149 14909 10183 14943
rect 10183 14909 10192 14943
rect 10140 14900 10192 14909
rect 15752 14943 15804 14952
rect 15752 14909 15761 14943
rect 15761 14909 15795 14943
rect 15795 14909 15804 14943
rect 15752 14900 15804 14909
rect 16120 14968 16172 15020
rect 17684 14968 17736 15020
rect 26424 15036 26476 15088
rect 22008 14968 22060 15020
rect 23480 14968 23532 15020
rect 26056 15011 26108 15020
rect 17500 14943 17552 14952
rect 17500 14909 17509 14943
rect 17509 14909 17543 14943
rect 17543 14909 17552 14943
rect 17500 14900 17552 14909
rect 26056 14977 26065 15011
rect 26065 14977 26099 15011
rect 26099 14977 26108 15011
rect 26056 14968 26108 14977
rect 30196 15011 30248 15020
rect 30196 14977 30205 15011
rect 30205 14977 30239 15011
rect 30239 14977 30248 15011
rect 30196 14968 30248 14977
rect 31484 14968 31536 15020
rect 33692 14968 33744 15020
rect 26976 14943 27028 14952
rect 26976 14909 26985 14943
rect 26985 14909 27019 14943
rect 27019 14909 27028 14943
rect 26976 14900 27028 14909
rect 34520 14943 34572 14952
rect 24492 14832 24544 14884
rect 34520 14909 34529 14943
rect 34529 14909 34563 14943
rect 34563 14909 34572 14943
rect 34520 14900 34572 14909
rect 8852 14807 8904 14816
rect 8852 14773 8861 14807
rect 8861 14773 8895 14807
rect 8895 14773 8904 14807
rect 8852 14764 8904 14773
rect 5674 14662 5726 14714
rect 5738 14662 5790 14714
rect 5802 14662 5854 14714
rect 5866 14662 5918 14714
rect 5930 14662 5982 14714
rect 15122 14662 15174 14714
rect 15186 14662 15238 14714
rect 15250 14662 15302 14714
rect 15314 14662 15366 14714
rect 15378 14662 15430 14714
rect 24570 14662 24622 14714
rect 24634 14662 24686 14714
rect 24698 14662 24750 14714
rect 24762 14662 24814 14714
rect 24826 14662 24878 14714
rect 34018 14662 34070 14714
rect 34082 14662 34134 14714
rect 34146 14662 34198 14714
rect 34210 14662 34262 14714
rect 34274 14662 34326 14714
rect 27252 14560 27304 14612
rect 31300 14603 31352 14612
rect 31300 14569 31309 14603
rect 31309 14569 31343 14603
rect 31343 14569 31352 14603
rect 31300 14560 31352 14569
rect 31484 14603 31536 14612
rect 31484 14569 31493 14603
rect 31493 14569 31527 14603
rect 31527 14569 31536 14603
rect 31484 14560 31536 14569
rect 33692 14603 33744 14612
rect 33692 14569 33701 14603
rect 33701 14569 33735 14603
rect 33735 14569 33744 14603
rect 33692 14560 33744 14569
rect 15752 14492 15804 14544
rect 1676 14399 1728 14408
rect 1676 14365 1685 14399
rect 1685 14365 1719 14399
rect 1719 14365 1728 14399
rect 1676 14356 1728 14365
rect 3792 14356 3844 14408
rect 9036 14424 9088 14476
rect 10324 14424 10376 14476
rect 15844 14424 15896 14476
rect 17500 14424 17552 14476
rect 21824 14467 21876 14476
rect 21824 14433 21833 14467
rect 21833 14433 21867 14467
rect 21867 14433 21876 14467
rect 21824 14424 21876 14433
rect 22468 14424 22520 14476
rect 23664 14424 23716 14476
rect 30656 14424 30708 14476
rect 9680 14399 9732 14408
rect 6000 14288 6052 14340
rect 7748 14288 7800 14340
rect 1492 14263 1544 14272
rect 1492 14229 1501 14263
rect 1501 14229 1535 14263
rect 1535 14229 1544 14263
rect 1492 14220 1544 14229
rect 7196 14263 7248 14272
rect 7196 14229 7205 14263
rect 7205 14229 7239 14263
rect 7239 14229 7248 14263
rect 9680 14365 9689 14399
rect 9689 14365 9723 14399
rect 9723 14365 9732 14399
rect 9680 14356 9732 14365
rect 15476 14399 15528 14408
rect 15476 14365 15485 14399
rect 15485 14365 15519 14399
rect 15519 14365 15528 14399
rect 15476 14356 15528 14365
rect 17592 14356 17644 14408
rect 19340 14356 19392 14408
rect 22192 14356 22244 14408
rect 26976 14356 27028 14408
rect 26056 14288 26108 14340
rect 32496 14356 32548 14408
rect 7196 14220 7248 14229
rect 20720 14220 20772 14272
rect 21916 14220 21968 14272
rect 22836 14220 22888 14272
rect 32036 14220 32088 14272
rect 35348 14220 35400 14272
rect 10398 14118 10450 14170
rect 10462 14118 10514 14170
rect 10526 14118 10578 14170
rect 10590 14118 10642 14170
rect 10654 14118 10706 14170
rect 19846 14118 19898 14170
rect 19910 14118 19962 14170
rect 19974 14118 20026 14170
rect 20038 14118 20090 14170
rect 20102 14118 20154 14170
rect 29294 14118 29346 14170
rect 29358 14118 29410 14170
rect 29422 14118 29474 14170
rect 29486 14118 29538 14170
rect 29550 14118 29602 14170
rect 7748 14059 7800 14068
rect 7748 14025 7757 14059
rect 7757 14025 7791 14059
rect 7791 14025 7800 14059
rect 7748 14016 7800 14025
rect 9588 14016 9640 14068
rect 22008 14016 22060 14068
rect 22192 14059 22244 14068
rect 22192 14025 22201 14059
rect 22201 14025 22235 14059
rect 22235 14025 22244 14059
rect 22192 14016 22244 14025
rect 15476 13948 15528 14000
rect 18236 13948 18288 14000
rect 20904 13948 20956 14000
rect 21088 13948 21140 14000
rect 21824 13948 21876 14000
rect 22560 13948 22612 14000
rect 23664 14016 23716 14068
rect 32496 14059 32548 14068
rect 32496 14025 32505 14059
rect 32505 14025 32539 14059
rect 32539 14025 32548 14059
rect 32496 14016 32548 14025
rect 23572 13948 23624 14000
rect 26240 13948 26292 14000
rect 17592 13923 17644 13932
rect 17592 13889 17601 13923
rect 17601 13889 17635 13923
rect 17635 13889 17644 13923
rect 17592 13880 17644 13889
rect 20720 13880 20772 13932
rect 21824 13855 21876 13864
rect 21824 13821 21833 13855
rect 21833 13821 21867 13855
rect 21867 13821 21876 13855
rect 21824 13812 21876 13821
rect 18052 13744 18104 13796
rect 21180 13744 21232 13796
rect 21916 13676 21968 13728
rect 22284 13812 22336 13864
rect 26332 13855 26384 13864
rect 26332 13821 26341 13855
rect 26341 13821 26375 13855
rect 26375 13821 26384 13855
rect 26332 13812 26384 13821
rect 32036 13880 32088 13932
rect 30288 13812 30340 13864
rect 27252 13719 27304 13728
rect 27252 13685 27261 13719
rect 27261 13685 27295 13719
rect 27295 13685 27304 13719
rect 27252 13676 27304 13685
rect 27436 13719 27488 13728
rect 27436 13685 27445 13719
rect 27445 13685 27479 13719
rect 27479 13685 27488 13719
rect 27436 13676 27488 13685
rect 5674 13574 5726 13626
rect 5738 13574 5790 13626
rect 5802 13574 5854 13626
rect 5866 13574 5918 13626
rect 5930 13574 5982 13626
rect 15122 13574 15174 13626
rect 15186 13574 15238 13626
rect 15250 13574 15302 13626
rect 15314 13574 15366 13626
rect 15378 13574 15430 13626
rect 24570 13574 24622 13626
rect 24634 13574 24686 13626
rect 24698 13574 24750 13626
rect 24762 13574 24814 13626
rect 24826 13574 24878 13626
rect 34018 13574 34070 13626
rect 34082 13574 34134 13626
rect 34146 13574 34198 13626
rect 34210 13574 34262 13626
rect 34274 13574 34326 13626
rect 6000 13472 6052 13524
rect 8852 13472 8904 13524
rect 1860 13404 1912 13456
rect 7288 13268 7340 13320
rect 7380 13311 7432 13320
rect 7380 13277 7389 13311
rect 7389 13277 7423 13311
rect 7423 13277 7432 13311
rect 7380 13268 7432 13277
rect 9312 13311 9364 13320
rect 9312 13277 9321 13311
rect 9321 13277 9355 13311
rect 9355 13277 9364 13311
rect 9312 13268 9364 13277
rect 21180 13472 21232 13524
rect 21272 13515 21324 13524
rect 21272 13481 21281 13515
rect 21281 13481 21315 13515
rect 21315 13481 21324 13515
rect 21272 13472 21324 13481
rect 26332 13472 26384 13524
rect 13820 13404 13872 13456
rect 2044 13132 2096 13184
rect 8944 13132 8996 13184
rect 24308 13404 24360 13456
rect 26056 13404 26108 13456
rect 16488 13336 16540 13388
rect 14556 13268 14608 13320
rect 19616 13336 19668 13388
rect 17684 13268 17736 13320
rect 19524 13311 19576 13320
rect 19524 13277 19533 13311
rect 19533 13277 19567 13311
rect 19567 13277 19576 13311
rect 19524 13268 19576 13277
rect 20904 13243 20956 13252
rect 20904 13209 20913 13243
rect 20913 13209 20947 13243
rect 20947 13209 20956 13243
rect 21916 13268 21968 13320
rect 22192 13311 22244 13320
rect 22192 13277 22201 13311
rect 22201 13277 22235 13311
rect 22235 13277 22244 13311
rect 22192 13268 22244 13277
rect 22468 13311 22520 13320
rect 22468 13277 22477 13311
rect 22477 13277 22511 13311
rect 22511 13277 22520 13311
rect 22468 13268 22520 13277
rect 25136 13268 25188 13320
rect 20904 13200 20956 13209
rect 25044 13200 25096 13252
rect 18788 13132 18840 13184
rect 20996 13132 21048 13184
rect 21916 13132 21968 13184
rect 23756 13132 23808 13184
rect 10398 13030 10450 13082
rect 10462 13030 10514 13082
rect 10526 13030 10578 13082
rect 10590 13030 10642 13082
rect 10654 13030 10706 13082
rect 19846 13030 19898 13082
rect 19910 13030 19962 13082
rect 19974 13030 20026 13082
rect 20038 13030 20090 13082
rect 20102 13030 20154 13082
rect 29294 13030 29346 13082
rect 29358 13030 29410 13082
rect 29422 13030 29474 13082
rect 29486 13030 29538 13082
rect 29550 13030 29602 13082
rect 3332 12928 3384 12980
rect 9312 12928 9364 12980
rect 19524 12928 19576 12980
rect 21916 12971 21968 12980
rect 21916 12937 21925 12971
rect 21925 12937 21959 12971
rect 21959 12937 21968 12971
rect 21916 12928 21968 12937
rect 26240 12928 26292 12980
rect 27160 12971 27212 12980
rect 27160 12937 27185 12971
rect 27185 12937 27212 12971
rect 27160 12928 27212 12937
rect 30564 12928 30616 12980
rect 31116 12928 31168 12980
rect 18788 12860 18840 12912
rect 19064 12860 19116 12912
rect 3148 12792 3200 12844
rect 1492 12631 1544 12640
rect 1492 12597 1501 12631
rect 1501 12597 1535 12631
rect 1535 12597 1544 12631
rect 1492 12588 1544 12597
rect 3148 12588 3200 12640
rect 3608 12588 3660 12640
rect 14464 12792 14516 12844
rect 14004 12767 14056 12776
rect 14004 12733 14013 12767
rect 14013 12733 14047 12767
rect 14047 12733 14056 12767
rect 14004 12724 14056 12733
rect 14372 12724 14424 12776
rect 18052 12724 18104 12776
rect 14648 12656 14700 12708
rect 13268 12631 13320 12640
rect 13268 12597 13277 12631
rect 13277 12597 13311 12631
rect 13311 12597 13320 12631
rect 13268 12588 13320 12597
rect 13636 12588 13688 12640
rect 13820 12631 13872 12640
rect 13820 12597 13829 12631
rect 13829 12597 13863 12631
rect 13863 12597 13872 12631
rect 13820 12588 13872 12597
rect 14832 12631 14884 12640
rect 14832 12597 14841 12631
rect 14841 12597 14875 12631
rect 14875 12597 14884 12631
rect 14832 12588 14884 12597
rect 19340 12835 19392 12844
rect 19340 12801 19349 12835
rect 19349 12801 19383 12835
rect 19383 12801 19392 12835
rect 22192 12860 22244 12912
rect 19340 12792 19392 12801
rect 22008 12835 22060 12844
rect 22008 12801 22017 12835
rect 22017 12801 22051 12835
rect 22051 12801 22060 12835
rect 22008 12792 22060 12801
rect 23756 12835 23808 12844
rect 23756 12801 23765 12835
rect 23765 12801 23799 12835
rect 23799 12801 23808 12835
rect 23756 12792 23808 12801
rect 19432 12724 19484 12776
rect 25044 12656 25096 12708
rect 19616 12588 19668 12640
rect 22468 12588 22520 12640
rect 31300 12860 31352 12912
rect 30288 12792 30340 12844
rect 31668 12860 31720 12912
rect 31944 12860 31996 12912
rect 35348 12835 35400 12844
rect 35348 12801 35357 12835
rect 35357 12801 35391 12835
rect 35391 12801 35400 12835
rect 35348 12792 35400 12801
rect 26424 12588 26476 12640
rect 27344 12631 27396 12640
rect 27344 12597 27353 12631
rect 27353 12597 27387 12631
rect 27387 12597 27396 12631
rect 27344 12588 27396 12597
rect 31760 12588 31812 12640
rect 36084 12588 36136 12640
rect 36360 12631 36412 12640
rect 36360 12597 36369 12631
rect 36369 12597 36403 12631
rect 36403 12597 36412 12631
rect 36360 12588 36412 12597
rect 5674 12486 5726 12538
rect 5738 12486 5790 12538
rect 5802 12486 5854 12538
rect 5866 12486 5918 12538
rect 5930 12486 5982 12538
rect 15122 12486 15174 12538
rect 15186 12486 15238 12538
rect 15250 12486 15302 12538
rect 15314 12486 15366 12538
rect 15378 12486 15430 12538
rect 24570 12486 24622 12538
rect 24634 12486 24686 12538
rect 24698 12486 24750 12538
rect 24762 12486 24814 12538
rect 24826 12486 24878 12538
rect 34018 12486 34070 12538
rect 34082 12486 34134 12538
rect 34146 12486 34198 12538
rect 34210 12486 34262 12538
rect 34274 12486 34326 12538
rect 5540 12384 5592 12436
rect 8852 12384 8904 12436
rect 31944 12427 31996 12436
rect 31944 12393 31953 12427
rect 31953 12393 31987 12427
rect 31987 12393 31996 12427
rect 31944 12384 31996 12393
rect 3792 12291 3844 12300
rect 3792 12257 3801 12291
rect 3801 12257 3835 12291
rect 3835 12257 3844 12291
rect 3792 12248 3844 12257
rect 14004 12316 14056 12368
rect 7288 12248 7340 12300
rect 12716 12248 12768 12300
rect 13728 12248 13780 12300
rect 14372 12291 14424 12300
rect 14372 12257 14381 12291
rect 14381 12257 14415 12291
rect 14415 12257 14424 12291
rect 14372 12248 14424 12257
rect 14832 12316 14884 12368
rect 34796 12248 34848 12300
rect 35348 12248 35400 12300
rect 4160 12223 4212 12232
rect 4160 12189 4169 12223
rect 4169 12189 4203 12223
rect 4203 12189 4212 12223
rect 4160 12180 4212 12189
rect 2136 12044 2188 12096
rect 5172 12112 5224 12164
rect 3148 12087 3200 12096
rect 3148 12053 3157 12087
rect 3157 12053 3191 12087
rect 3191 12053 3200 12087
rect 3148 12044 3200 12053
rect 3424 12044 3476 12096
rect 9588 12180 9640 12232
rect 13268 12223 13320 12232
rect 13268 12189 13277 12223
rect 13277 12189 13311 12223
rect 13311 12189 13320 12223
rect 13268 12180 13320 12189
rect 13636 12180 13688 12232
rect 26240 12180 26292 12232
rect 27344 12223 27396 12232
rect 27344 12189 27353 12223
rect 27353 12189 27387 12223
rect 27387 12189 27396 12223
rect 27344 12180 27396 12189
rect 36084 12223 36136 12232
rect 36084 12189 36093 12223
rect 36093 12189 36127 12223
rect 36127 12189 36136 12223
rect 36084 12180 36136 12189
rect 14372 12112 14424 12164
rect 9220 12087 9272 12096
rect 9220 12053 9229 12087
rect 9229 12053 9263 12087
rect 9263 12053 9272 12087
rect 9220 12044 9272 12053
rect 13176 12044 13228 12096
rect 14464 12044 14516 12096
rect 16488 12112 16540 12164
rect 14648 12087 14700 12096
rect 14648 12053 14657 12087
rect 14657 12053 14691 12087
rect 14691 12053 14700 12087
rect 25228 12087 25280 12096
rect 14648 12044 14700 12053
rect 25228 12053 25237 12087
rect 25237 12053 25271 12087
rect 25271 12053 25280 12087
rect 31760 12112 31812 12164
rect 25228 12044 25280 12053
rect 27252 12044 27304 12096
rect 34520 12044 34572 12096
rect 35808 12044 35860 12096
rect 36360 12044 36412 12096
rect 10398 11942 10450 11994
rect 10462 11942 10514 11994
rect 10526 11942 10578 11994
rect 10590 11942 10642 11994
rect 10654 11942 10706 11994
rect 19846 11942 19898 11994
rect 19910 11942 19962 11994
rect 19974 11942 20026 11994
rect 20038 11942 20090 11994
rect 20102 11942 20154 11994
rect 29294 11942 29346 11994
rect 29358 11942 29410 11994
rect 29422 11942 29474 11994
rect 29486 11942 29538 11994
rect 29550 11942 29602 11994
rect 4160 11840 4212 11892
rect 5172 11840 5224 11892
rect 9128 11840 9180 11892
rect 12716 11883 12768 11892
rect 10048 11772 10100 11824
rect 3424 11747 3476 11756
rect 3424 11713 3433 11747
rect 3433 11713 3467 11747
rect 3467 11713 3476 11747
rect 3424 11704 3476 11713
rect 3608 11747 3660 11756
rect 3608 11713 3617 11747
rect 3617 11713 3651 11747
rect 3651 11713 3660 11747
rect 3608 11704 3660 11713
rect 9220 11704 9272 11756
rect 12716 11849 12725 11883
rect 12725 11849 12759 11883
rect 12759 11849 12768 11883
rect 12716 11840 12768 11849
rect 14464 11883 14516 11892
rect 14464 11849 14473 11883
rect 14473 11849 14507 11883
rect 14507 11849 14516 11883
rect 14464 11840 14516 11849
rect 14556 11883 14608 11892
rect 14556 11849 14565 11883
rect 14565 11849 14599 11883
rect 14599 11849 14608 11883
rect 14556 11840 14608 11849
rect 13176 11815 13228 11824
rect 13176 11781 13185 11815
rect 13185 11781 13219 11815
rect 13219 11781 13228 11815
rect 13176 11772 13228 11781
rect 25044 11772 25096 11824
rect 11796 11704 11848 11756
rect 13636 11704 13688 11756
rect 14372 11704 14424 11756
rect 14740 11704 14792 11756
rect 18052 11747 18104 11756
rect 18052 11713 18061 11747
rect 18061 11713 18095 11747
rect 18095 11713 18104 11747
rect 18052 11704 18104 11713
rect 18236 11747 18288 11756
rect 18236 11713 18245 11747
rect 18245 11713 18279 11747
rect 18279 11713 18288 11747
rect 18236 11704 18288 11713
rect 27252 11747 27304 11756
rect 27252 11713 27261 11747
rect 27261 11713 27295 11747
rect 27295 11713 27304 11747
rect 27252 11704 27304 11713
rect 28724 11747 28776 11756
rect 28724 11713 28733 11747
rect 28733 11713 28767 11747
rect 28767 11713 28776 11747
rect 28724 11704 28776 11713
rect 3332 11679 3384 11688
rect 3332 11645 3341 11679
rect 3341 11645 3375 11679
rect 3375 11645 3384 11679
rect 3332 11636 3384 11645
rect 10140 11636 10192 11688
rect 13820 11568 13872 11620
rect 16672 11568 16724 11620
rect 1492 11543 1544 11552
rect 1492 11509 1501 11543
rect 1501 11509 1535 11543
rect 1535 11509 1544 11543
rect 1492 11500 1544 11509
rect 2228 11543 2280 11552
rect 2228 11509 2237 11543
rect 2237 11509 2271 11543
rect 2271 11509 2280 11543
rect 2228 11500 2280 11509
rect 6276 11500 6328 11552
rect 9956 11500 10008 11552
rect 14280 11543 14332 11552
rect 14280 11509 14289 11543
rect 14289 11509 14323 11543
rect 14323 11509 14332 11543
rect 18052 11543 18104 11552
rect 14280 11500 14332 11509
rect 18052 11509 18061 11543
rect 18061 11509 18095 11543
rect 18095 11509 18104 11543
rect 18052 11500 18104 11509
rect 34520 11500 34572 11552
rect 5674 11398 5726 11450
rect 5738 11398 5790 11450
rect 5802 11398 5854 11450
rect 5866 11398 5918 11450
rect 5930 11398 5982 11450
rect 15122 11398 15174 11450
rect 15186 11398 15238 11450
rect 15250 11398 15302 11450
rect 15314 11398 15366 11450
rect 15378 11398 15430 11450
rect 24570 11398 24622 11450
rect 24634 11398 24686 11450
rect 24698 11398 24750 11450
rect 24762 11398 24814 11450
rect 24826 11398 24878 11450
rect 34018 11398 34070 11450
rect 34082 11398 34134 11450
rect 34146 11398 34198 11450
rect 34210 11398 34262 11450
rect 34274 11398 34326 11450
rect 10048 11339 10100 11348
rect 10048 11305 10057 11339
rect 10057 11305 10091 11339
rect 10091 11305 10100 11339
rect 10048 11296 10100 11305
rect 13636 11296 13688 11348
rect 14280 11296 14332 11348
rect 25228 11296 25280 11348
rect 28724 11296 28776 11348
rect 31760 11296 31812 11348
rect 2228 11228 2280 11280
rect 14556 11228 14608 11280
rect 14832 11228 14884 11280
rect 16672 11160 16724 11212
rect 10140 11135 10192 11144
rect 10140 11101 10149 11135
rect 10149 11101 10183 11135
rect 10183 11101 10192 11135
rect 10140 11092 10192 11101
rect 13268 11092 13320 11144
rect 14648 11092 14700 11144
rect 16028 11092 16080 11144
rect 16488 11135 16540 11144
rect 16488 11101 16497 11135
rect 16497 11101 16531 11135
rect 16531 11101 16540 11135
rect 16488 11092 16540 11101
rect 33692 11228 33744 11280
rect 31484 11160 31536 11212
rect 32220 11160 32272 11212
rect 23572 11024 23624 11076
rect 23756 11024 23808 11076
rect 24492 11024 24544 11076
rect 31484 11067 31536 11076
rect 31484 11033 31493 11067
rect 31493 11033 31527 11067
rect 31527 11033 31536 11067
rect 31484 11024 31536 11033
rect 32036 11024 32088 11076
rect 16672 10999 16724 11008
rect 16672 10965 16681 10999
rect 16681 10965 16715 10999
rect 16715 10965 16724 10999
rect 16672 10956 16724 10965
rect 31852 10999 31904 11008
rect 31852 10965 31861 10999
rect 31861 10965 31895 10999
rect 31895 10965 31904 10999
rect 31852 10956 31904 10965
rect 10398 10854 10450 10906
rect 10462 10854 10514 10906
rect 10526 10854 10578 10906
rect 10590 10854 10642 10906
rect 10654 10854 10706 10906
rect 19846 10854 19898 10906
rect 19910 10854 19962 10906
rect 19974 10854 20026 10906
rect 20038 10854 20090 10906
rect 20102 10854 20154 10906
rect 29294 10854 29346 10906
rect 29358 10854 29410 10906
rect 29422 10854 29474 10906
rect 29486 10854 29538 10906
rect 29550 10854 29602 10906
rect 3332 10752 3384 10804
rect 18052 10795 18104 10804
rect 7104 10727 7156 10736
rect 7104 10693 7131 10727
rect 7131 10693 7156 10727
rect 7104 10684 7156 10693
rect 18052 10761 18061 10795
rect 18061 10761 18095 10795
rect 18095 10761 18104 10795
rect 18052 10752 18104 10761
rect 22928 10795 22980 10804
rect 14556 10684 14608 10736
rect 16672 10684 16724 10736
rect 17868 10684 17920 10736
rect 19064 10684 19116 10736
rect 22928 10761 22937 10795
rect 22937 10761 22971 10795
rect 22971 10761 22980 10795
rect 22928 10752 22980 10761
rect 32036 10752 32088 10804
rect 35808 10795 35860 10804
rect 22468 10727 22520 10736
rect 22468 10693 22477 10727
rect 22477 10693 22511 10727
rect 22511 10693 22520 10727
rect 22468 10684 22520 10693
rect 35808 10761 35817 10795
rect 35817 10761 35851 10795
rect 35851 10761 35860 10795
rect 35808 10752 35860 10761
rect 18972 10616 19024 10668
rect 31852 10616 31904 10668
rect 33692 10659 33744 10668
rect 33692 10625 33701 10659
rect 33701 10625 33735 10659
rect 33735 10625 33744 10659
rect 33692 10616 33744 10625
rect 34796 10659 34848 10668
rect 34796 10625 34805 10659
rect 34805 10625 34839 10659
rect 34839 10625 34848 10659
rect 34796 10616 34848 10625
rect 4896 10412 4948 10464
rect 7380 10412 7432 10464
rect 17592 10412 17644 10464
rect 18972 10455 19024 10464
rect 18972 10421 18981 10455
rect 18981 10421 19015 10455
rect 19015 10421 19024 10455
rect 18972 10412 19024 10421
rect 35716 10412 35768 10464
rect 5674 10310 5726 10362
rect 5738 10310 5790 10362
rect 5802 10310 5854 10362
rect 5866 10310 5918 10362
rect 5930 10310 5982 10362
rect 15122 10310 15174 10362
rect 15186 10310 15238 10362
rect 15250 10310 15302 10362
rect 15314 10310 15366 10362
rect 15378 10310 15430 10362
rect 24570 10310 24622 10362
rect 24634 10310 24686 10362
rect 24698 10310 24750 10362
rect 24762 10310 24814 10362
rect 24826 10310 24878 10362
rect 34018 10310 34070 10362
rect 34082 10310 34134 10362
rect 34146 10310 34198 10362
rect 34210 10310 34262 10362
rect 34274 10310 34326 10362
rect 35808 10208 35860 10260
rect 16028 10115 16080 10124
rect 16028 10081 16037 10115
rect 16037 10081 16071 10115
rect 16071 10081 16080 10115
rect 16028 10072 16080 10081
rect 16672 10072 16724 10124
rect 34796 10072 34848 10124
rect 4896 10047 4948 10056
rect 4896 10013 4905 10047
rect 4905 10013 4939 10047
rect 4939 10013 4948 10047
rect 4896 10004 4948 10013
rect 27436 10047 27488 10056
rect 27436 10013 27445 10047
rect 27445 10013 27479 10047
rect 27479 10013 27488 10047
rect 27436 10004 27488 10013
rect 35716 10004 35768 10056
rect 20812 9936 20864 9988
rect 1492 9911 1544 9920
rect 1492 9877 1501 9911
rect 1501 9877 1535 9911
rect 1535 9877 1544 9911
rect 1492 9868 1544 9877
rect 4712 9911 4764 9920
rect 4712 9877 4721 9911
rect 4721 9877 4755 9911
rect 4755 9877 4764 9911
rect 4712 9868 4764 9877
rect 27436 9868 27488 9920
rect 10398 9766 10450 9818
rect 10462 9766 10514 9818
rect 10526 9766 10578 9818
rect 10590 9766 10642 9818
rect 10654 9766 10706 9818
rect 19846 9766 19898 9818
rect 19910 9766 19962 9818
rect 19974 9766 20026 9818
rect 20038 9766 20090 9818
rect 20102 9766 20154 9818
rect 29294 9766 29346 9818
rect 29358 9766 29410 9818
rect 29422 9766 29474 9818
rect 29486 9766 29538 9818
rect 29550 9766 29602 9818
rect 13268 9596 13320 9648
rect 18972 9596 19024 9648
rect 22468 9596 22520 9648
rect 22008 9528 22060 9580
rect 22928 9571 22980 9580
rect 22928 9537 22937 9571
rect 22937 9537 22971 9571
rect 22971 9537 22980 9571
rect 22928 9528 22980 9537
rect 24400 9571 24452 9580
rect 24400 9537 24409 9571
rect 24409 9537 24443 9571
rect 24443 9537 24452 9571
rect 24400 9528 24452 9537
rect 20260 9460 20312 9512
rect 26792 9460 26844 9512
rect 30656 9460 30708 9512
rect 1952 9392 2004 9444
rect 3700 9392 3752 9444
rect 6920 9435 6972 9444
rect 6920 9401 6929 9435
rect 6929 9401 6963 9435
rect 6963 9401 6972 9435
rect 6920 9392 6972 9401
rect 4988 9324 5040 9376
rect 6644 9324 6696 9376
rect 20628 9324 20680 9376
rect 30380 9392 30432 9444
rect 27160 9324 27212 9376
rect 30472 9324 30524 9376
rect 5674 9222 5726 9274
rect 5738 9222 5790 9274
rect 5802 9222 5854 9274
rect 5866 9222 5918 9274
rect 5930 9222 5982 9274
rect 15122 9222 15174 9274
rect 15186 9222 15238 9274
rect 15250 9222 15302 9274
rect 15314 9222 15366 9274
rect 15378 9222 15430 9274
rect 24570 9222 24622 9274
rect 24634 9222 24686 9274
rect 24698 9222 24750 9274
rect 24762 9222 24814 9274
rect 24826 9222 24878 9274
rect 34018 9222 34070 9274
rect 34082 9222 34134 9274
rect 34146 9222 34198 9274
rect 34210 9222 34262 9274
rect 34274 9222 34326 9274
rect 22008 9163 22060 9172
rect 2872 8984 2924 9036
rect 22008 9129 22017 9163
rect 22017 9129 22051 9163
rect 22051 9129 22060 9163
rect 22008 9120 22060 9129
rect 22468 9120 22520 9172
rect 24400 9120 24452 9172
rect 3700 9052 3752 9104
rect 2688 8891 2740 8900
rect 2688 8857 2697 8891
rect 2697 8857 2731 8891
rect 2731 8857 2740 8891
rect 2688 8848 2740 8857
rect 4988 8984 5040 9036
rect 21088 9027 21140 9036
rect 21088 8993 21097 9027
rect 21097 8993 21131 9027
rect 21131 8993 21140 9027
rect 21088 8984 21140 8993
rect 6644 8959 6696 8968
rect 6644 8925 6653 8959
rect 6653 8925 6687 8959
rect 6687 8925 6696 8959
rect 6644 8916 6696 8925
rect 17868 8916 17920 8968
rect 20812 8916 20864 8968
rect 13820 8848 13872 8900
rect 22284 8916 22336 8968
rect 22468 8984 22520 9036
rect 26792 9120 26844 9172
rect 31944 9120 31996 9172
rect 1492 8823 1544 8832
rect 1492 8789 1501 8823
rect 1501 8789 1535 8823
rect 1535 8789 1544 8823
rect 1492 8780 1544 8789
rect 2872 8823 2924 8832
rect 2872 8789 2897 8823
rect 2897 8789 2924 8823
rect 2872 8780 2924 8789
rect 3700 8780 3752 8832
rect 6184 8780 6236 8832
rect 7380 8823 7432 8832
rect 7380 8789 7389 8823
rect 7389 8789 7423 8823
rect 7423 8789 7432 8823
rect 7380 8780 7432 8789
rect 8852 8780 8904 8832
rect 20628 8780 20680 8832
rect 24768 8916 24820 8968
rect 31668 9052 31720 9104
rect 27436 9027 27488 9036
rect 27436 8993 27445 9027
rect 27445 8993 27479 9027
rect 27479 8993 27488 9027
rect 27436 8984 27488 8993
rect 27160 8959 27212 8968
rect 27160 8925 27169 8959
rect 27169 8925 27203 8959
rect 27203 8925 27212 8959
rect 27160 8916 27212 8925
rect 30656 8916 30708 8968
rect 24860 8848 24912 8900
rect 30472 8848 30524 8900
rect 28724 8780 28776 8832
rect 30748 8823 30800 8832
rect 30748 8789 30757 8823
rect 30757 8789 30791 8823
rect 30791 8789 30800 8823
rect 30748 8780 30800 8789
rect 10398 8678 10450 8730
rect 10462 8678 10514 8730
rect 10526 8678 10578 8730
rect 10590 8678 10642 8730
rect 10654 8678 10706 8730
rect 19846 8678 19898 8730
rect 19910 8678 19962 8730
rect 19974 8678 20026 8730
rect 20038 8678 20090 8730
rect 20102 8678 20154 8730
rect 29294 8678 29346 8730
rect 29358 8678 29410 8730
rect 29422 8678 29474 8730
rect 29486 8678 29538 8730
rect 29550 8678 29602 8730
rect 2688 8576 2740 8628
rect 4988 8619 5040 8628
rect 4988 8585 4997 8619
rect 4997 8585 5031 8619
rect 5031 8585 5040 8619
rect 4988 8576 5040 8585
rect 7012 8619 7064 8628
rect 7012 8585 7039 8619
rect 7039 8585 7064 8619
rect 7012 8576 7064 8585
rect 8852 8619 8904 8628
rect 2964 8508 3016 8560
rect 7104 8508 7156 8560
rect 7380 8508 7432 8560
rect 8852 8585 8861 8619
rect 8861 8585 8895 8619
rect 8895 8585 8904 8619
rect 8852 8576 8904 8585
rect 3700 8483 3752 8492
rect 3700 8449 3709 8483
rect 3709 8449 3743 8483
rect 3743 8449 3752 8483
rect 3700 8440 3752 8449
rect 4436 8347 4488 8356
rect 4436 8313 4445 8347
rect 4445 8313 4479 8347
rect 4479 8313 4488 8347
rect 4436 8304 4488 8313
rect 6920 8304 6972 8356
rect 7748 8304 7800 8356
rect 18972 8576 19024 8628
rect 13820 8508 13872 8560
rect 10140 8440 10192 8492
rect 13728 8440 13780 8492
rect 17776 8483 17828 8492
rect 17776 8449 17785 8483
rect 17785 8449 17819 8483
rect 17819 8449 17828 8483
rect 17776 8440 17828 8449
rect 30288 8576 30340 8628
rect 30472 8619 30524 8628
rect 30472 8585 30481 8619
rect 30481 8585 30515 8619
rect 30515 8585 30524 8619
rect 30472 8576 30524 8585
rect 34428 8576 34480 8628
rect 20628 8551 20680 8560
rect 20628 8517 20637 8551
rect 20637 8517 20671 8551
rect 20671 8517 20680 8551
rect 20628 8508 20680 8517
rect 20812 8551 20864 8560
rect 20812 8517 20821 8551
rect 20821 8517 20855 8551
rect 20855 8517 20864 8551
rect 20812 8508 20864 8517
rect 21088 8508 21140 8560
rect 23480 8508 23532 8560
rect 22284 8483 22336 8492
rect 17500 8415 17552 8424
rect 17500 8381 17509 8415
rect 17509 8381 17543 8415
rect 17543 8381 17552 8415
rect 17500 8372 17552 8381
rect 3240 8279 3292 8288
rect 3240 8245 3249 8279
rect 3249 8245 3283 8279
rect 3283 8245 3292 8279
rect 3240 8236 3292 8245
rect 4068 8236 4120 8288
rect 7564 8236 7616 8288
rect 22284 8449 22293 8483
rect 22293 8449 22327 8483
rect 22327 8449 22336 8483
rect 22284 8440 22336 8449
rect 22468 8440 22520 8492
rect 24768 8440 24820 8492
rect 20260 8372 20312 8424
rect 24860 8372 24912 8424
rect 23020 8347 23072 8356
rect 23020 8313 23029 8347
rect 23029 8313 23063 8347
rect 23063 8313 23072 8347
rect 23020 8304 23072 8313
rect 30380 8508 30432 8560
rect 30748 8440 30800 8492
rect 31668 8508 31720 8560
rect 27436 8372 27488 8424
rect 27620 8415 27672 8424
rect 27620 8381 27629 8415
rect 27629 8381 27663 8415
rect 27663 8381 27672 8415
rect 27620 8372 27672 8381
rect 28724 8372 28776 8424
rect 33140 8372 33192 8424
rect 30288 8304 30340 8356
rect 33784 8304 33836 8356
rect 13084 8279 13136 8288
rect 13084 8245 13093 8279
rect 13093 8245 13127 8279
rect 13127 8245 13136 8279
rect 13084 8236 13136 8245
rect 23756 8279 23808 8288
rect 23756 8245 23765 8279
rect 23765 8245 23799 8279
rect 23799 8245 23808 8279
rect 23756 8236 23808 8245
rect 30472 8236 30524 8288
rect 32036 8236 32088 8288
rect 5674 8134 5726 8186
rect 5738 8134 5790 8186
rect 5802 8134 5854 8186
rect 5866 8134 5918 8186
rect 5930 8134 5982 8186
rect 15122 8134 15174 8186
rect 15186 8134 15238 8186
rect 15250 8134 15302 8186
rect 15314 8134 15366 8186
rect 15378 8134 15430 8186
rect 24570 8134 24622 8186
rect 24634 8134 24686 8186
rect 24698 8134 24750 8186
rect 24762 8134 24814 8186
rect 24826 8134 24878 8186
rect 34018 8134 34070 8186
rect 34082 8134 34134 8186
rect 34146 8134 34198 8186
rect 34210 8134 34262 8186
rect 34274 8134 34326 8186
rect 7288 8032 7340 8084
rect 23480 8075 23532 8084
rect 23480 8041 23489 8075
rect 23489 8041 23523 8075
rect 23523 8041 23532 8075
rect 23480 8032 23532 8041
rect 31116 8075 31168 8084
rect 31116 8041 31125 8075
rect 31125 8041 31159 8075
rect 31159 8041 31168 8075
rect 31116 8032 31168 8041
rect 32036 8032 32088 8084
rect 32128 7964 32180 8016
rect 9036 7896 9088 7948
rect 11796 7939 11848 7948
rect 11796 7905 11805 7939
rect 11805 7905 11839 7939
rect 11839 7905 11848 7939
rect 11796 7896 11848 7905
rect 18236 7896 18288 7948
rect 3240 7828 3292 7880
rect 3792 7871 3844 7880
rect 3792 7837 3801 7871
rect 3801 7837 3835 7871
rect 3835 7837 3844 7871
rect 3792 7828 3844 7837
rect 4068 7871 4120 7880
rect 4068 7837 4077 7871
rect 4077 7837 4111 7871
rect 4111 7837 4120 7871
rect 4068 7828 4120 7837
rect 13728 7828 13780 7880
rect 27620 7828 27672 7880
rect 3148 7760 3200 7812
rect 3608 7692 3660 7744
rect 7380 7760 7432 7812
rect 9496 7760 9548 7812
rect 9956 7760 10008 7812
rect 12072 7803 12124 7812
rect 12072 7769 12081 7803
rect 12081 7769 12115 7803
rect 12115 7769 12124 7803
rect 12072 7760 12124 7769
rect 13084 7760 13136 7812
rect 6092 7692 6144 7744
rect 7104 7692 7156 7744
rect 7564 7735 7616 7744
rect 7564 7701 7573 7735
rect 7573 7701 7607 7735
rect 7607 7701 7616 7735
rect 7564 7692 7616 7701
rect 18052 7760 18104 7812
rect 14096 7692 14148 7744
rect 30104 7692 30156 7744
rect 33784 7871 33836 7880
rect 33784 7837 33793 7871
rect 33793 7837 33827 7871
rect 33827 7837 33836 7871
rect 33784 7828 33836 7837
rect 34428 7828 34480 7880
rect 35440 7828 35492 7880
rect 33968 7735 34020 7744
rect 33968 7701 33977 7735
rect 33977 7701 34011 7735
rect 34011 7701 34020 7735
rect 33968 7692 34020 7701
rect 36728 7735 36780 7744
rect 36728 7701 36737 7735
rect 36737 7701 36771 7735
rect 36771 7701 36780 7735
rect 36728 7692 36780 7701
rect 10398 7590 10450 7642
rect 10462 7590 10514 7642
rect 10526 7590 10578 7642
rect 10590 7590 10642 7642
rect 10654 7590 10706 7642
rect 19846 7590 19898 7642
rect 19910 7590 19962 7642
rect 19974 7590 20026 7642
rect 20038 7590 20090 7642
rect 20102 7590 20154 7642
rect 29294 7590 29346 7642
rect 29358 7590 29410 7642
rect 29422 7590 29474 7642
rect 29486 7590 29538 7642
rect 29550 7590 29602 7642
rect 7380 7531 7432 7540
rect 7380 7497 7389 7531
rect 7389 7497 7423 7531
rect 7423 7497 7432 7531
rect 7380 7488 7432 7497
rect 9956 7531 10008 7540
rect 9956 7497 9965 7531
rect 9965 7497 9999 7531
rect 9999 7497 10008 7531
rect 9956 7488 10008 7497
rect 11796 7488 11848 7540
rect 10140 7352 10192 7404
rect 30748 7488 30800 7540
rect 36452 7531 36504 7540
rect 36452 7497 36461 7531
rect 36461 7497 36495 7531
rect 36495 7497 36504 7531
rect 36452 7488 36504 7497
rect 36728 7488 36780 7540
rect 17408 7420 17460 7472
rect 23020 7420 23072 7472
rect 30380 7420 30432 7472
rect 14096 7352 14148 7404
rect 18236 7395 18288 7404
rect 18236 7361 18245 7395
rect 18245 7361 18279 7395
rect 18279 7361 18288 7395
rect 18236 7352 18288 7361
rect 33968 7352 34020 7404
rect 12164 7284 12216 7336
rect 12992 7327 13044 7336
rect 12992 7293 13001 7327
rect 13001 7293 13035 7327
rect 13035 7293 13044 7327
rect 12992 7284 13044 7293
rect 22008 7284 22060 7336
rect 35440 7327 35492 7336
rect 35440 7293 35449 7327
rect 35449 7293 35483 7327
rect 35483 7293 35492 7327
rect 35440 7284 35492 7293
rect 1492 7191 1544 7200
rect 1492 7157 1501 7191
rect 1501 7157 1535 7191
rect 1535 7157 1544 7191
rect 1492 7148 1544 7157
rect 7288 7148 7340 7200
rect 17960 7148 18012 7200
rect 18052 7191 18104 7200
rect 18052 7157 18061 7191
rect 18061 7157 18095 7191
rect 18095 7157 18104 7191
rect 30104 7191 30156 7200
rect 18052 7148 18104 7157
rect 30104 7157 30113 7191
rect 30113 7157 30147 7191
rect 30147 7157 30156 7191
rect 30104 7148 30156 7157
rect 32036 7148 32088 7200
rect 5674 7046 5726 7098
rect 5738 7046 5790 7098
rect 5802 7046 5854 7098
rect 5866 7046 5918 7098
rect 5930 7046 5982 7098
rect 15122 7046 15174 7098
rect 15186 7046 15238 7098
rect 15250 7046 15302 7098
rect 15314 7046 15366 7098
rect 15378 7046 15430 7098
rect 24570 7046 24622 7098
rect 24634 7046 24686 7098
rect 24698 7046 24750 7098
rect 24762 7046 24814 7098
rect 24826 7046 24878 7098
rect 34018 7046 34070 7098
rect 34082 7046 34134 7098
rect 34146 7046 34198 7098
rect 34210 7046 34262 7098
rect 34274 7046 34326 7098
rect 12992 6944 13044 6996
rect 30380 6944 30432 6996
rect 30840 6944 30892 6996
rect 31484 6944 31536 6996
rect 7564 6876 7616 6928
rect 17408 6876 17460 6928
rect 17500 6876 17552 6928
rect 19708 6876 19760 6928
rect 18052 6808 18104 6860
rect 6920 6783 6972 6792
rect 6920 6749 6929 6783
rect 6929 6749 6963 6783
rect 6963 6749 6972 6783
rect 6920 6740 6972 6749
rect 17960 6783 18012 6792
rect 17960 6749 17969 6783
rect 17969 6749 18003 6783
rect 18003 6749 18012 6783
rect 17960 6740 18012 6749
rect 19524 6783 19576 6792
rect 19524 6749 19533 6783
rect 19533 6749 19567 6783
rect 19567 6749 19576 6783
rect 19524 6740 19576 6749
rect 26516 6783 26568 6792
rect 26516 6749 26525 6783
rect 26525 6749 26559 6783
rect 26559 6749 26568 6783
rect 26516 6740 26568 6749
rect 26884 6740 26936 6792
rect 31668 6740 31720 6792
rect 32036 6783 32088 6792
rect 32036 6749 32045 6783
rect 32045 6749 32079 6783
rect 32079 6749 32088 6783
rect 32036 6740 32088 6749
rect 6644 6604 6696 6656
rect 17776 6647 17828 6656
rect 17776 6613 17785 6647
rect 17785 6613 17819 6647
rect 17819 6613 17828 6647
rect 17776 6604 17828 6613
rect 18328 6604 18380 6656
rect 30748 6604 30800 6656
rect 32404 6604 32456 6656
rect 34888 6647 34940 6656
rect 34888 6613 34897 6647
rect 34897 6613 34931 6647
rect 34931 6613 34940 6647
rect 34888 6604 34940 6613
rect 10398 6502 10450 6554
rect 10462 6502 10514 6554
rect 10526 6502 10578 6554
rect 10590 6502 10642 6554
rect 10654 6502 10706 6554
rect 19846 6502 19898 6554
rect 19910 6502 19962 6554
rect 19974 6502 20026 6554
rect 20038 6502 20090 6554
rect 20102 6502 20154 6554
rect 29294 6502 29346 6554
rect 29358 6502 29410 6554
rect 29422 6502 29474 6554
rect 29486 6502 29538 6554
rect 29550 6502 29602 6554
rect 31668 6400 31720 6452
rect 33140 6443 33192 6452
rect 33140 6409 33149 6443
rect 33149 6409 33183 6443
rect 33183 6409 33192 6443
rect 36452 6443 36504 6452
rect 33140 6400 33192 6409
rect 36452 6409 36461 6443
rect 36461 6409 36495 6443
rect 36495 6409 36504 6443
rect 36452 6400 36504 6409
rect 3792 6332 3844 6384
rect 1584 6264 1636 6316
rect 3608 6307 3660 6316
rect 3608 6273 3617 6307
rect 3617 6273 3651 6307
rect 3651 6273 3660 6307
rect 3608 6264 3660 6273
rect 18236 6332 18288 6384
rect 6184 6264 6236 6316
rect 32128 6307 32180 6316
rect 32128 6273 32137 6307
rect 32137 6273 32171 6307
rect 32171 6273 32180 6307
rect 32128 6264 32180 6273
rect 32404 6307 32456 6316
rect 32404 6273 32413 6307
rect 32413 6273 32447 6307
rect 32447 6273 32456 6307
rect 32404 6264 32456 6273
rect 34888 6264 34940 6316
rect 35440 6239 35492 6248
rect 35440 6205 35449 6239
rect 35449 6205 35483 6239
rect 35483 6205 35492 6239
rect 35440 6196 35492 6205
rect 20536 6128 20588 6180
rect 1492 6103 1544 6112
rect 1492 6069 1501 6103
rect 1501 6069 1535 6103
rect 1535 6069 1544 6103
rect 1492 6060 1544 6069
rect 3148 6060 3200 6112
rect 30840 6103 30892 6112
rect 30840 6069 30849 6103
rect 30849 6069 30883 6103
rect 30883 6069 30892 6103
rect 30840 6060 30892 6069
rect 5674 5958 5726 6010
rect 5738 5958 5790 6010
rect 5802 5958 5854 6010
rect 5866 5958 5918 6010
rect 5930 5958 5982 6010
rect 15122 5958 15174 6010
rect 15186 5958 15238 6010
rect 15250 5958 15302 6010
rect 15314 5958 15366 6010
rect 15378 5958 15430 6010
rect 24570 5958 24622 6010
rect 24634 5958 24686 6010
rect 24698 5958 24750 6010
rect 24762 5958 24814 6010
rect 24826 5958 24878 6010
rect 34018 5958 34070 6010
rect 34082 5958 34134 6010
rect 34146 5958 34198 6010
rect 34210 5958 34262 6010
rect 34274 5958 34326 6010
rect 7288 5856 7340 5908
rect 30104 5856 30156 5908
rect 19708 5788 19760 5840
rect 23204 5831 23256 5840
rect 23204 5797 23213 5831
rect 23213 5797 23247 5831
rect 23247 5797 23256 5831
rect 23204 5788 23256 5797
rect 22008 5720 22060 5772
rect 6184 5695 6236 5704
rect 6184 5661 6193 5695
rect 6193 5661 6227 5695
rect 6227 5661 6236 5695
rect 6184 5652 6236 5661
rect 20260 5652 20312 5704
rect 22376 5652 22428 5704
rect 26884 5652 26936 5704
rect 27620 5695 27672 5704
rect 27620 5661 27629 5695
rect 27629 5661 27663 5695
rect 27663 5661 27672 5695
rect 27620 5652 27672 5661
rect 6368 5559 6420 5568
rect 6368 5525 6377 5559
rect 6377 5525 6411 5559
rect 6411 5525 6420 5559
rect 6368 5516 6420 5525
rect 28540 5516 28592 5568
rect 10398 5414 10450 5466
rect 10462 5414 10514 5466
rect 10526 5414 10578 5466
rect 10590 5414 10642 5466
rect 10654 5414 10706 5466
rect 19846 5414 19898 5466
rect 19910 5414 19962 5466
rect 19974 5414 20026 5466
rect 20038 5414 20090 5466
rect 20102 5414 20154 5466
rect 29294 5414 29346 5466
rect 29358 5414 29410 5466
rect 29422 5414 29474 5466
rect 29486 5414 29538 5466
rect 29550 5414 29602 5466
rect 22468 5355 22520 5364
rect 22468 5321 22477 5355
rect 22477 5321 22511 5355
rect 22511 5321 22520 5355
rect 22468 5312 22520 5321
rect 26516 5312 26568 5364
rect 19432 5287 19484 5296
rect 19432 5253 19441 5287
rect 19441 5253 19475 5287
rect 19475 5253 19484 5287
rect 19432 5244 19484 5253
rect 20260 5244 20312 5296
rect 6184 5176 6236 5228
rect 6644 5219 6696 5228
rect 6644 5185 6653 5219
rect 6653 5185 6687 5219
rect 6687 5185 6696 5219
rect 6644 5176 6696 5185
rect 20076 5219 20128 5228
rect 20076 5185 20085 5219
rect 20085 5185 20119 5219
rect 20119 5185 20128 5219
rect 20076 5176 20128 5185
rect 20536 5176 20588 5228
rect 22376 5219 22428 5228
rect 22376 5185 22385 5219
rect 22385 5185 22419 5219
rect 22419 5185 22428 5219
rect 22376 5176 22428 5185
rect 22560 5219 22612 5228
rect 22560 5185 22569 5219
rect 22569 5185 22603 5219
rect 22603 5185 22612 5219
rect 22560 5176 22612 5185
rect 27160 5219 27212 5228
rect 27160 5185 27169 5219
rect 27169 5185 27203 5219
rect 27203 5185 27212 5219
rect 27160 5176 27212 5185
rect 19524 5108 19576 5160
rect 20260 5151 20312 5160
rect 20260 5117 20269 5151
rect 20269 5117 20303 5151
rect 20303 5117 20312 5151
rect 20260 5108 20312 5117
rect 24400 5040 24452 5092
rect 7472 4972 7524 5024
rect 20168 5015 20220 5024
rect 20168 4981 20177 5015
rect 20177 4981 20211 5015
rect 20211 4981 20220 5015
rect 20168 4972 20220 4981
rect 5674 4870 5726 4922
rect 5738 4870 5790 4922
rect 5802 4870 5854 4922
rect 5866 4870 5918 4922
rect 5930 4870 5982 4922
rect 15122 4870 15174 4922
rect 15186 4870 15238 4922
rect 15250 4870 15302 4922
rect 15314 4870 15366 4922
rect 15378 4870 15430 4922
rect 24570 4870 24622 4922
rect 24634 4870 24686 4922
rect 24698 4870 24750 4922
rect 24762 4870 24814 4922
rect 24826 4870 24878 4922
rect 34018 4870 34070 4922
rect 34082 4870 34134 4922
rect 34146 4870 34198 4922
rect 34210 4870 34262 4922
rect 34274 4870 34326 4922
rect 2872 4811 2924 4820
rect 2872 4777 2881 4811
rect 2881 4777 2915 4811
rect 2915 4777 2924 4811
rect 2872 4768 2924 4777
rect 4252 4768 4304 4820
rect 19432 4811 19484 4820
rect 19432 4777 19441 4811
rect 19441 4777 19475 4811
rect 19475 4777 19484 4811
rect 19432 4768 19484 4777
rect 20260 4811 20312 4820
rect 20260 4777 20269 4811
rect 20269 4777 20303 4811
rect 20303 4777 20312 4811
rect 20260 4768 20312 4777
rect 22560 4768 22612 4820
rect 3148 4564 3200 4616
rect 6092 4607 6144 4616
rect 6092 4573 6101 4607
rect 6101 4573 6135 4607
rect 6135 4573 6144 4607
rect 6092 4564 6144 4573
rect 7748 4607 7800 4616
rect 7748 4573 7757 4607
rect 7757 4573 7791 4607
rect 7791 4573 7800 4607
rect 7748 4564 7800 4573
rect 14832 4607 14884 4616
rect 14832 4573 14841 4607
rect 14841 4573 14875 4607
rect 14875 4573 14884 4607
rect 14832 4564 14884 4573
rect 31852 4700 31904 4752
rect 23204 4632 23256 4684
rect 20168 4564 20220 4616
rect 20076 4496 20128 4548
rect 20536 4564 20588 4616
rect 27620 4607 27672 4616
rect 20444 4496 20496 4548
rect 22376 4496 22428 4548
rect 27344 4539 27396 4548
rect 27344 4505 27353 4539
rect 27353 4505 27387 4539
rect 27387 4505 27396 4539
rect 27344 4496 27396 4505
rect 27620 4573 27629 4607
rect 27629 4573 27663 4607
rect 27663 4573 27672 4607
rect 27620 4564 27672 4573
rect 28540 4564 28592 4616
rect 1492 4471 1544 4480
rect 1492 4437 1501 4471
rect 1501 4437 1535 4471
rect 1535 4437 1544 4471
rect 1492 4428 1544 4437
rect 5540 4428 5592 4480
rect 7564 4471 7616 4480
rect 7564 4437 7573 4471
rect 7573 4437 7607 4471
rect 7607 4437 7616 4471
rect 7564 4428 7616 4437
rect 14280 4428 14332 4480
rect 15568 4471 15620 4480
rect 15568 4437 15577 4471
rect 15577 4437 15611 4471
rect 15611 4437 15620 4471
rect 15568 4428 15620 4437
rect 23480 4428 23532 4480
rect 27620 4428 27672 4480
rect 10398 4326 10450 4378
rect 10462 4326 10514 4378
rect 10526 4326 10578 4378
rect 10590 4326 10642 4378
rect 10654 4326 10706 4378
rect 19846 4326 19898 4378
rect 19910 4326 19962 4378
rect 19974 4326 20026 4378
rect 20038 4326 20090 4378
rect 20102 4326 20154 4378
rect 29294 4326 29346 4378
rect 29358 4326 29410 4378
rect 29422 4326 29474 4378
rect 29486 4326 29538 4378
rect 29550 4326 29602 4378
rect 3148 4267 3200 4276
rect 3148 4233 3157 4267
rect 3157 4233 3191 4267
rect 3191 4233 3200 4267
rect 3148 4224 3200 4233
rect 4068 4224 4120 4276
rect 7472 4267 7524 4276
rect 7472 4233 7481 4267
rect 7481 4233 7515 4267
rect 7515 4233 7524 4267
rect 7472 4224 7524 4233
rect 27160 4224 27212 4276
rect 27528 4224 27580 4276
rect 2872 4020 2924 4072
rect 2872 3884 2924 3936
rect 4712 4088 4764 4140
rect 5540 4131 5592 4140
rect 5540 4097 5549 4131
rect 5549 4097 5583 4131
rect 5583 4097 5592 4131
rect 5540 4088 5592 4097
rect 6368 4088 6420 4140
rect 7564 4088 7616 4140
rect 11980 4088 12032 4140
rect 14280 4131 14332 4140
rect 14280 4097 14289 4131
rect 14289 4097 14323 4131
rect 14323 4097 14332 4131
rect 14280 4088 14332 4097
rect 14372 4088 14424 4140
rect 14464 4088 14516 4140
rect 18328 4131 18380 4140
rect 18328 4097 18337 4131
rect 18337 4097 18371 4131
rect 18371 4097 18380 4131
rect 18328 4088 18380 4097
rect 10508 4063 10560 4072
rect 10508 4029 10517 4063
rect 10517 4029 10551 4063
rect 10551 4029 10560 4063
rect 10508 4020 10560 4029
rect 9496 3995 9548 4004
rect 9496 3961 9505 3995
rect 9505 3961 9539 3995
rect 9539 3961 9548 3995
rect 9496 3952 9548 3961
rect 4252 3884 4304 3936
rect 7472 3884 7524 3936
rect 10784 3884 10836 3936
rect 15568 4020 15620 4072
rect 14188 3995 14240 4004
rect 14188 3961 14197 3995
rect 14197 3961 14231 3995
rect 14231 3961 14240 3995
rect 14188 3952 14240 3961
rect 17500 4020 17552 4072
rect 23756 4156 23808 4208
rect 27620 4199 27672 4208
rect 27620 4165 27629 4199
rect 27629 4165 27663 4199
rect 27663 4165 27672 4199
rect 27620 4156 27672 4165
rect 20260 4131 20312 4140
rect 20260 4097 20269 4131
rect 20269 4097 20303 4131
rect 20303 4097 20312 4131
rect 20260 4088 20312 4097
rect 20444 4131 20496 4140
rect 20444 4097 20453 4131
rect 20453 4097 20487 4131
rect 20487 4097 20496 4131
rect 20444 4088 20496 4097
rect 23480 4131 23532 4140
rect 23480 4097 23489 4131
rect 23489 4097 23523 4131
rect 23523 4097 23532 4131
rect 23480 4088 23532 4097
rect 27988 4088 28040 4140
rect 30840 4088 30892 4140
rect 14372 3884 14424 3936
rect 14924 3927 14976 3936
rect 14924 3893 14933 3927
rect 14933 3893 14967 3927
rect 14967 3893 14976 3927
rect 14924 3884 14976 3893
rect 19708 3927 19760 3936
rect 19708 3893 19717 3927
rect 19717 3893 19751 3927
rect 19751 3893 19760 3927
rect 19708 3884 19760 3893
rect 20260 3927 20312 3936
rect 20260 3893 20269 3927
rect 20269 3893 20303 3927
rect 20303 3893 20312 3927
rect 20260 3884 20312 3893
rect 24308 3884 24360 3936
rect 28540 3884 28592 3936
rect 5674 3782 5726 3834
rect 5738 3782 5790 3834
rect 5802 3782 5854 3834
rect 5866 3782 5918 3834
rect 5930 3782 5982 3834
rect 15122 3782 15174 3834
rect 15186 3782 15238 3834
rect 15250 3782 15302 3834
rect 15314 3782 15366 3834
rect 15378 3782 15430 3834
rect 24570 3782 24622 3834
rect 24634 3782 24686 3834
rect 24698 3782 24750 3834
rect 24762 3782 24814 3834
rect 24826 3782 24878 3834
rect 34018 3782 34070 3834
rect 34082 3782 34134 3834
rect 34146 3782 34198 3834
rect 34210 3782 34262 3834
rect 34274 3782 34326 3834
rect 12072 3680 12124 3732
rect 14188 3680 14240 3732
rect 16764 3723 16816 3732
rect 16764 3689 16773 3723
rect 16773 3689 16807 3723
rect 16807 3689 16816 3723
rect 16764 3680 16816 3689
rect 20720 3680 20772 3732
rect 31760 3680 31812 3732
rect 36820 3723 36872 3732
rect 36820 3689 36829 3723
rect 36829 3689 36863 3723
rect 36863 3689 36872 3723
rect 36820 3680 36872 3689
rect 11980 3655 12032 3664
rect 11980 3621 11989 3655
rect 11989 3621 12023 3655
rect 12023 3621 12032 3655
rect 11980 3612 12032 3621
rect 10508 3587 10560 3596
rect 10508 3553 10517 3587
rect 10517 3553 10551 3587
rect 10551 3553 10560 3587
rect 10508 3544 10560 3553
rect 2872 3519 2924 3528
rect 1492 3383 1544 3392
rect 1492 3349 1501 3383
rect 1501 3349 1535 3383
rect 1535 3349 1544 3383
rect 1492 3340 1544 3349
rect 2872 3485 2881 3519
rect 2881 3485 2915 3519
rect 2915 3485 2924 3519
rect 2872 3476 2924 3485
rect 10784 3519 10836 3528
rect 10784 3485 10793 3519
rect 10793 3485 10827 3519
rect 10827 3485 10836 3519
rect 10784 3476 10836 3485
rect 14372 3612 14424 3664
rect 12440 3519 12492 3528
rect 12440 3485 12449 3519
rect 12449 3485 12483 3519
rect 12483 3485 12492 3519
rect 12440 3476 12492 3485
rect 14464 3544 14516 3596
rect 14648 3587 14700 3596
rect 14648 3553 14657 3587
rect 14657 3553 14691 3587
rect 14691 3553 14700 3587
rect 31300 3612 31352 3664
rect 14648 3544 14700 3553
rect 14372 3519 14424 3528
rect 14372 3485 14381 3519
rect 14381 3485 14415 3519
rect 14415 3485 14424 3519
rect 14372 3476 14424 3485
rect 20260 3544 20312 3596
rect 22928 3544 22980 3596
rect 24400 3544 24452 3596
rect 26884 3587 26936 3596
rect 26884 3553 26893 3587
rect 26893 3553 26927 3587
rect 26927 3553 26936 3587
rect 26884 3544 26936 3553
rect 31576 3587 31628 3596
rect 31576 3553 31585 3587
rect 31585 3553 31619 3587
rect 31619 3553 31628 3587
rect 31576 3544 31628 3553
rect 33692 3544 33744 3596
rect 14188 3408 14240 3460
rect 14556 3340 14608 3392
rect 19248 3476 19300 3528
rect 21364 3519 21416 3528
rect 21364 3485 21373 3519
rect 21373 3485 21407 3519
rect 21407 3485 21416 3519
rect 21364 3476 21416 3485
rect 27344 3476 27396 3528
rect 27988 3519 28040 3528
rect 27988 3485 27997 3519
rect 27997 3485 28031 3519
rect 28031 3485 28040 3519
rect 27988 3476 28040 3485
rect 28540 3476 28592 3528
rect 31392 3476 31444 3528
rect 31852 3476 31904 3528
rect 32404 3519 32456 3528
rect 32404 3485 32413 3519
rect 32413 3485 32447 3519
rect 32447 3485 32456 3519
rect 32404 3476 32456 3485
rect 16856 3451 16908 3460
rect 16856 3417 16865 3451
rect 16865 3417 16899 3451
rect 16899 3417 16908 3451
rect 16856 3408 16908 3417
rect 22468 3408 22520 3460
rect 29000 3408 29052 3460
rect 30012 3451 30064 3460
rect 30012 3417 30021 3451
rect 30021 3417 30055 3451
rect 30055 3417 30064 3451
rect 30012 3408 30064 3417
rect 33232 3408 33284 3460
rect 16672 3340 16724 3392
rect 23480 3383 23532 3392
rect 23480 3349 23489 3383
rect 23489 3349 23523 3383
rect 23523 3349 23532 3383
rect 23480 3340 23532 3349
rect 31024 3383 31076 3392
rect 31024 3349 31033 3383
rect 31033 3349 31067 3383
rect 31067 3349 31076 3383
rect 31024 3340 31076 3349
rect 37924 3476 37976 3528
rect 37648 3408 37700 3460
rect 37280 3340 37332 3392
rect 38108 3383 38160 3392
rect 38108 3349 38117 3383
rect 38117 3349 38151 3383
rect 38151 3349 38160 3383
rect 38108 3340 38160 3349
rect 10398 3238 10450 3290
rect 10462 3238 10514 3290
rect 10526 3238 10578 3290
rect 10590 3238 10642 3290
rect 10654 3238 10706 3290
rect 19846 3238 19898 3290
rect 19910 3238 19962 3290
rect 19974 3238 20026 3290
rect 20038 3238 20090 3290
rect 20102 3238 20154 3290
rect 29294 3238 29346 3290
rect 29358 3238 29410 3290
rect 29422 3238 29474 3290
rect 29486 3238 29538 3290
rect 29550 3238 29602 3290
rect 2136 3179 2188 3188
rect 2136 3145 2145 3179
rect 2145 3145 2179 3179
rect 2179 3145 2188 3179
rect 2136 3136 2188 3145
rect 5540 3136 5592 3188
rect 12440 3136 12492 3188
rect 37924 3179 37976 3188
rect 37924 3145 37933 3179
rect 37933 3145 37967 3179
rect 37967 3145 37976 3179
rect 37924 3136 37976 3145
rect 14372 3068 14424 3120
rect 14556 3111 14608 3120
rect 14556 3077 14565 3111
rect 14565 3077 14599 3111
rect 14599 3077 14608 3111
rect 14556 3068 14608 3077
rect 14924 3068 14976 3120
rect 31024 3068 31076 3120
rect 31576 3111 31628 3120
rect 31576 3077 31585 3111
rect 31585 3077 31619 3111
rect 31619 3077 31628 3111
rect 31576 3068 31628 3077
rect 23572 3000 23624 3052
rect 24308 3043 24360 3052
rect 24308 3009 24317 3043
rect 24317 3009 24351 3043
rect 24351 3009 24360 3043
rect 24308 3000 24360 3009
rect 24400 3000 24452 3052
rect 31300 3043 31352 3052
rect 31300 3009 31309 3043
rect 31309 3009 31343 3043
rect 31343 3009 31352 3043
rect 31300 3000 31352 3009
rect 31392 3043 31444 3052
rect 31392 3009 31401 3043
rect 31401 3009 31435 3043
rect 31435 3009 31444 3043
rect 38108 3043 38160 3052
rect 31392 3000 31444 3009
rect 38108 3009 38117 3043
rect 38117 3009 38151 3043
rect 38151 3009 38160 3043
rect 38108 3000 38160 3009
rect 39120 3000 39172 3052
rect 14648 2932 14700 2984
rect 17592 2932 17644 2984
rect 38016 2932 38068 2984
rect 27528 2864 27580 2916
rect 2228 2796 2280 2848
rect 12808 2839 12860 2848
rect 12808 2805 12817 2839
rect 12817 2805 12851 2839
rect 12851 2805 12860 2839
rect 12808 2796 12860 2805
rect 14004 2796 14056 2848
rect 14188 2796 14240 2848
rect 17592 2839 17644 2848
rect 17592 2805 17601 2839
rect 17601 2805 17635 2839
rect 17635 2805 17644 2839
rect 17592 2796 17644 2805
rect 20260 2796 20312 2848
rect 28356 2839 28408 2848
rect 28356 2805 28365 2839
rect 28365 2805 28399 2839
rect 28399 2805 28408 2839
rect 28356 2796 28408 2805
rect 31944 2796 31996 2848
rect 34520 2839 34572 2848
rect 34520 2805 34529 2839
rect 34529 2805 34563 2839
rect 34563 2805 34572 2839
rect 34520 2796 34572 2805
rect 36728 2796 36780 2848
rect 37464 2796 37516 2848
rect 5674 2694 5726 2746
rect 5738 2694 5790 2746
rect 5802 2694 5854 2746
rect 5866 2694 5918 2746
rect 5930 2694 5982 2746
rect 15122 2694 15174 2746
rect 15186 2694 15238 2746
rect 15250 2694 15302 2746
rect 15314 2694 15366 2746
rect 15378 2694 15430 2746
rect 24570 2694 24622 2746
rect 24634 2694 24686 2746
rect 24698 2694 24750 2746
rect 24762 2694 24814 2746
rect 24826 2694 24878 2746
rect 34018 2694 34070 2746
rect 34082 2694 34134 2746
rect 34146 2694 34198 2746
rect 34210 2694 34262 2746
rect 34274 2694 34326 2746
rect 14188 2592 14240 2644
rect 14372 2592 14424 2644
rect 16672 2635 16724 2644
rect 16672 2601 16681 2635
rect 16681 2601 16715 2635
rect 16715 2601 16724 2635
rect 16672 2592 16724 2601
rect 16856 2592 16908 2644
rect 19248 2635 19300 2644
rect 19248 2601 19257 2635
rect 19257 2601 19291 2635
rect 19291 2601 19300 2635
rect 19248 2592 19300 2601
rect 20720 2592 20772 2644
rect 21364 2592 21416 2644
rect 22468 2635 22520 2644
rect 22468 2601 22477 2635
rect 22477 2601 22511 2635
rect 22511 2601 22520 2635
rect 22468 2592 22520 2601
rect 22928 2592 22980 2644
rect 29000 2592 29052 2644
rect 30012 2592 30064 2644
rect 31760 2592 31812 2644
rect 32404 2592 32456 2644
rect 33232 2635 33284 2644
rect 33232 2601 33241 2635
rect 33241 2601 33275 2635
rect 33275 2601 33284 2635
rect 33232 2592 33284 2601
rect 33692 2592 33744 2644
rect 36820 2592 36872 2644
rect 37280 2635 37332 2644
rect 37280 2601 37289 2635
rect 37289 2601 37323 2635
rect 37323 2601 37332 2635
rect 37280 2592 37332 2601
rect 37648 2592 37700 2644
rect 14832 2524 14884 2576
rect 16764 2524 16816 2576
rect 2136 2456 2188 2508
rect 2228 2388 2280 2440
rect 4436 2456 4488 2508
rect 5540 2388 5592 2440
rect 6276 2388 6328 2440
rect 7196 2431 7248 2440
rect 7196 2397 7205 2431
rect 7205 2397 7239 2431
rect 7239 2397 7248 2431
rect 7196 2388 7248 2397
rect 8392 2431 8444 2440
rect 8392 2397 8401 2431
rect 8401 2397 8435 2431
rect 8435 2397 8444 2431
rect 8392 2388 8444 2397
rect 12440 2388 12492 2440
rect 12808 2388 12860 2440
rect 14004 2388 14056 2440
rect 15200 2388 15252 2440
rect 16396 2388 16448 2440
rect 17592 2388 17644 2440
rect 18788 2388 18840 2440
rect 20260 2388 20312 2440
rect 19708 2320 19760 2372
rect 22376 2388 22428 2440
rect 23572 2388 23624 2440
rect 27988 2456 28040 2508
rect 27528 2431 27580 2440
rect 27528 2397 27537 2431
rect 27537 2397 27571 2431
rect 27571 2397 27580 2431
rect 27528 2388 27580 2397
rect 28356 2388 28408 2440
rect 29644 2431 29696 2440
rect 29644 2397 29653 2431
rect 29653 2397 29687 2431
rect 29687 2397 29696 2431
rect 29644 2388 29696 2397
rect 30748 2388 30800 2440
rect 31944 2388 31996 2440
rect 33140 2388 33192 2440
rect 34520 2388 34572 2440
rect 35532 2388 35584 2440
rect 37464 2431 37516 2440
rect 37464 2397 37473 2431
rect 37473 2397 37507 2431
rect 37507 2397 37516 2431
rect 37464 2388 37516 2397
rect 38016 2388 38068 2440
rect 1492 2295 1544 2304
rect 1492 2261 1501 2295
rect 1501 2261 1535 2295
rect 1535 2261 1544 2295
rect 1492 2252 1544 2261
rect 2044 2252 2096 2304
rect 3240 2295 3292 2304
rect 3240 2261 3249 2295
rect 3249 2261 3283 2295
rect 3283 2261 3292 2295
rect 3240 2252 3292 2261
rect 4436 2252 4488 2304
rect 5632 2295 5684 2304
rect 5632 2261 5641 2295
rect 5641 2261 5675 2295
rect 5675 2261 5684 2295
rect 5632 2252 5684 2261
rect 6828 2252 6880 2304
rect 8024 2252 8076 2304
rect 9220 2252 9272 2304
rect 11612 2252 11664 2304
rect 18788 2252 18840 2304
rect 21180 2295 21232 2304
rect 21180 2261 21189 2295
rect 21189 2261 21223 2295
rect 21223 2261 21232 2295
rect 21180 2252 21232 2261
rect 24768 2252 24820 2304
rect 27160 2252 27212 2304
rect 10398 2150 10450 2202
rect 10462 2150 10514 2202
rect 10526 2150 10578 2202
rect 10590 2150 10642 2202
rect 10654 2150 10706 2202
rect 19846 2150 19898 2202
rect 19910 2150 19962 2202
rect 19974 2150 20026 2202
rect 20038 2150 20090 2202
rect 20102 2150 20154 2202
rect 29294 2150 29346 2202
rect 29358 2150 29410 2202
rect 29422 2150 29474 2202
rect 29486 2150 29538 2202
rect 29550 2150 29602 2202
<< metal2 >>
rect 2870 35200 2926 36000
rect 8574 35200 8630 36000
rect 14278 35200 14334 36000
rect 19982 35306 20038 36000
rect 25686 35306 25742 36000
rect 19982 35278 20300 35306
rect 19982 35200 20038 35278
rect 1398 34368 1454 34377
rect 1398 34303 1454 34312
rect 1412 33114 1440 34303
rect 1492 33312 1544 33318
rect 1492 33254 1544 33260
rect 1400 33108 1452 33114
rect 1400 33050 1452 33056
rect 1504 33017 1532 33254
rect 1490 33008 1546 33017
rect 1490 32943 1546 32952
rect 2228 32768 2280 32774
rect 2228 32710 2280 32716
rect 2240 32570 2268 32710
rect 2228 32564 2280 32570
rect 2228 32506 2280 32512
rect 1768 32224 1820 32230
rect 1768 32166 1820 32172
rect 1492 31680 1544 31686
rect 1490 31648 1492 31657
rect 1544 31648 1546 31657
rect 1490 31583 1546 31592
rect 1676 30728 1728 30734
rect 1676 30670 1728 30676
rect 1492 30592 1544 30598
rect 1492 30534 1544 30540
rect 1504 30297 1532 30534
rect 1490 30288 1546 30297
rect 1490 30223 1546 30232
rect 1688 29850 1716 30670
rect 1676 29844 1728 29850
rect 1676 29786 1728 29792
rect 1492 29028 1544 29034
rect 1492 28970 1544 28976
rect 1504 28937 1532 28970
rect 1490 28928 1546 28937
rect 1490 28863 1546 28872
rect 1492 27872 1544 27878
rect 1492 27814 1544 27820
rect 1504 27577 1532 27814
rect 1490 27568 1546 27577
rect 1490 27503 1546 27512
rect 1492 26240 1544 26246
rect 1490 26208 1492 26217
rect 1780 26234 1808 32166
rect 2688 31816 2740 31822
rect 2688 31758 2740 31764
rect 2700 31482 2728 31758
rect 2688 31476 2740 31482
rect 2688 31418 2740 31424
rect 2884 30818 2912 35200
rect 8588 33590 8616 35200
rect 10398 33756 10706 33765
rect 10398 33754 10404 33756
rect 10460 33754 10484 33756
rect 10540 33754 10564 33756
rect 10620 33754 10644 33756
rect 10700 33754 10706 33756
rect 10460 33702 10462 33754
rect 10642 33702 10644 33754
rect 10398 33700 10404 33702
rect 10460 33700 10484 33702
rect 10540 33700 10564 33702
rect 10620 33700 10644 33702
rect 10700 33700 10706 33702
rect 10398 33691 10706 33700
rect 19846 33756 20154 33765
rect 19846 33754 19852 33756
rect 19908 33754 19932 33756
rect 19988 33754 20012 33756
rect 20068 33754 20092 33756
rect 20148 33754 20154 33756
rect 19908 33702 19910 33754
rect 20090 33702 20092 33754
rect 19846 33700 19852 33702
rect 19908 33700 19932 33702
rect 19988 33700 20012 33702
rect 20068 33700 20092 33702
rect 20148 33700 20154 33702
rect 19846 33691 20154 33700
rect 8576 33584 8628 33590
rect 8576 33526 8628 33532
rect 9128 33584 9180 33590
rect 9128 33526 9180 33532
rect 5674 33212 5982 33221
rect 5674 33210 5680 33212
rect 5736 33210 5760 33212
rect 5816 33210 5840 33212
rect 5896 33210 5920 33212
rect 5976 33210 5982 33212
rect 5736 33158 5738 33210
rect 5918 33158 5920 33210
rect 5674 33156 5680 33158
rect 5736 33156 5760 33158
rect 5816 33156 5840 33158
rect 5896 33156 5920 33158
rect 5976 33156 5982 33158
rect 5674 33147 5982 33156
rect 9140 33114 9168 33526
rect 20272 33522 20300 35278
rect 25686 35278 25820 35306
rect 25686 35200 25742 35278
rect 25792 33522 25820 35278
rect 31390 35200 31446 36000
rect 31496 35278 31708 35306
rect 31404 35170 31432 35200
rect 31496 35170 31524 35278
rect 31404 35142 31524 35170
rect 29294 33756 29602 33765
rect 29294 33754 29300 33756
rect 29356 33754 29380 33756
rect 29436 33754 29460 33756
rect 29516 33754 29540 33756
rect 29596 33754 29602 33756
rect 29356 33702 29358 33754
rect 29538 33702 29540 33754
rect 29294 33700 29300 33702
rect 29356 33700 29380 33702
rect 29436 33700 29460 33702
rect 29516 33700 29540 33702
rect 29596 33700 29602 33702
rect 29294 33691 29602 33700
rect 14096 33516 14148 33522
rect 14096 33458 14148 33464
rect 20260 33516 20312 33522
rect 20260 33458 20312 33464
rect 25780 33516 25832 33522
rect 31680 33504 31708 35278
rect 37094 35200 37150 36000
rect 37108 33522 37136 35200
rect 31760 33516 31812 33522
rect 31680 33476 31760 33504
rect 25780 33458 25832 33464
rect 31760 33458 31812 33464
rect 37096 33516 37148 33522
rect 37096 33458 37148 33464
rect 9404 33312 9456 33318
rect 9404 33254 9456 33260
rect 9128 33108 9180 33114
rect 9128 33050 9180 33056
rect 9036 32972 9088 32978
rect 9036 32914 9088 32920
rect 9048 32502 9076 32914
rect 9036 32496 9088 32502
rect 9036 32438 9088 32444
rect 3332 32428 3384 32434
rect 3332 32370 3384 32376
rect 6644 32428 6696 32434
rect 6644 32370 6696 32376
rect 3344 32026 3372 32370
rect 3976 32360 4028 32366
rect 3976 32302 4028 32308
rect 3332 32020 3384 32026
rect 3332 31962 3384 31968
rect 3424 31340 3476 31346
rect 3424 31282 3476 31288
rect 3148 31272 3200 31278
rect 3148 31214 3200 31220
rect 2792 30790 2912 30818
rect 2044 29028 2096 29034
rect 2044 28970 2096 28976
rect 1544 26208 1546 26217
rect 1490 26143 1546 26152
rect 1688 26206 1808 26234
rect 1492 25152 1544 25158
rect 1492 25094 1544 25100
rect 1504 24857 1532 25094
rect 1490 24848 1546 24857
rect 1490 24783 1546 24792
rect 1492 23520 1544 23526
rect 1490 23488 1492 23497
rect 1544 23488 1546 23497
rect 1490 23423 1546 23432
rect 1400 22432 1452 22438
rect 1400 22374 1452 22380
rect 1412 22137 1440 22374
rect 1398 22128 1454 22137
rect 1398 22063 1454 22072
rect 1492 20800 1544 20806
rect 1490 20768 1492 20777
rect 1544 20768 1546 20777
rect 1490 20703 1546 20712
rect 1492 19712 1544 19718
rect 1492 19654 1544 19660
rect 1504 19417 1532 19654
rect 1490 19408 1546 19417
rect 1490 19343 1546 19352
rect 1492 18080 1544 18086
rect 1490 18048 1492 18057
rect 1544 18048 1546 18057
rect 1490 17983 1546 17992
rect 1492 16992 1544 16998
rect 1492 16934 1544 16940
rect 1504 16697 1532 16934
rect 1584 16720 1636 16726
rect 1490 16688 1546 16697
rect 1584 16662 1636 16668
rect 1490 16623 1546 16632
rect 1492 15360 1544 15366
rect 1490 15328 1492 15337
rect 1544 15328 1546 15337
rect 1490 15263 1546 15272
rect 1492 14272 1544 14278
rect 1492 14214 1544 14220
rect 1504 13977 1532 14214
rect 1490 13968 1546 13977
rect 1490 13903 1546 13912
rect 1492 12640 1544 12646
rect 1490 12608 1492 12617
rect 1544 12608 1546 12617
rect 1490 12543 1546 12552
rect 1492 11552 1544 11558
rect 1492 11494 1544 11500
rect 1504 11257 1532 11494
rect 1490 11248 1546 11257
rect 1490 11183 1546 11192
rect 1492 9920 1544 9926
rect 1490 9888 1492 9897
rect 1544 9888 1546 9897
rect 1490 9823 1546 9832
rect 1492 8832 1544 8838
rect 1492 8774 1544 8780
rect 1504 8537 1532 8774
rect 1490 8528 1546 8537
rect 1490 8463 1546 8472
rect 1492 7200 1544 7206
rect 1490 7168 1492 7177
rect 1544 7168 1546 7177
rect 1490 7103 1546 7112
rect 1596 6322 1624 16662
rect 1688 14414 1716 26206
rect 1860 23724 1912 23730
rect 1860 23666 1912 23672
rect 1768 20936 1820 20942
rect 1768 20878 1820 20884
rect 1780 20602 1808 20878
rect 1768 20596 1820 20602
rect 1768 20538 1820 20544
rect 1676 14408 1728 14414
rect 1676 14350 1728 14356
rect 1872 13462 1900 23666
rect 1952 18284 2004 18290
rect 1952 18226 2004 18232
rect 1964 18086 1992 18226
rect 1952 18080 2004 18086
rect 1952 18022 2004 18028
rect 1860 13456 1912 13462
rect 1860 13398 1912 13404
rect 1964 9450 1992 18022
rect 2056 13190 2084 28970
rect 2320 27872 2372 27878
rect 2320 27814 2372 27820
rect 2228 25152 2280 25158
rect 2228 25094 2280 25100
rect 2240 24954 2268 25094
rect 2228 24948 2280 24954
rect 2228 24890 2280 24896
rect 2332 24818 2360 27814
rect 2412 26376 2464 26382
rect 2412 26318 2464 26324
rect 2424 25702 2452 26318
rect 2412 25696 2464 25702
rect 2412 25638 2464 25644
rect 2320 24812 2372 24818
rect 2320 24754 2372 24760
rect 2228 20800 2280 20806
rect 2228 20742 2280 20748
rect 2240 18086 2268 20742
rect 2792 20602 2820 30790
rect 2964 29640 3016 29646
rect 2964 29582 3016 29588
rect 2976 29034 3004 29582
rect 2964 29028 3016 29034
rect 2964 28970 3016 28976
rect 2872 27464 2924 27470
rect 2872 27406 2924 27412
rect 2884 26586 2912 27406
rect 2872 26580 2924 26586
rect 2872 26522 2924 26528
rect 2976 26382 3004 28970
rect 3056 27600 3108 27606
rect 3056 27542 3108 27548
rect 3068 27130 3096 27542
rect 3056 27124 3108 27130
rect 3056 27066 3108 27072
rect 2964 26376 3016 26382
rect 2964 26318 3016 26324
rect 3068 26234 3096 27066
rect 3160 26382 3188 31214
rect 3436 30258 3464 31282
rect 3988 30802 4016 32302
rect 4988 32224 5040 32230
rect 4988 32166 5040 32172
rect 5000 30938 5028 32166
rect 5674 32124 5982 32133
rect 5674 32122 5680 32124
rect 5736 32122 5760 32124
rect 5816 32122 5840 32124
rect 5896 32122 5920 32124
rect 5976 32122 5982 32124
rect 5736 32070 5738 32122
rect 5918 32070 5920 32122
rect 5674 32068 5680 32070
rect 5736 32068 5760 32070
rect 5816 32068 5840 32070
rect 5896 32068 5920 32070
rect 5976 32068 5982 32070
rect 5674 32059 5982 32068
rect 6656 32026 6684 32370
rect 8024 32224 8076 32230
rect 8024 32166 8076 32172
rect 6644 32020 6696 32026
rect 6644 31962 6696 31968
rect 8036 31958 8064 32166
rect 8024 31952 8076 31958
rect 8024 31894 8076 31900
rect 6460 31816 6512 31822
rect 6460 31758 6512 31764
rect 6472 31482 6500 31758
rect 8036 31482 8064 31894
rect 8760 31680 8812 31686
rect 8760 31622 8812 31628
rect 6460 31476 6512 31482
rect 6460 31418 6512 31424
rect 8024 31476 8076 31482
rect 8024 31418 8076 31424
rect 8772 31346 8800 31622
rect 9048 31346 9076 32438
rect 9128 31816 9180 31822
rect 9128 31758 9180 31764
rect 6552 31340 6604 31346
rect 6552 31282 6604 31288
rect 8760 31340 8812 31346
rect 8760 31282 8812 31288
rect 9036 31340 9088 31346
rect 9036 31282 9088 31288
rect 5674 31036 5982 31045
rect 5674 31034 5680 31036
rect 5736 31034 5760 31036
rect 5816 31034 5840 31036
rect 5896 31034 5920 31036
rect 5976 31034 5982 31036
rect 5736 30982 5738 31034
rect 5918 30982 5920 31034
rect 5674 30980 5680 30982
rect 5736 30980 5760 30982
rect 5816 30980 5840 30982
rect 5896 30980 5920 30982
rect 5976 30980 5982 30982
rect 5674 30971 5982 30980
rect 4988 30932 5040 30938
rect 4988 30874 5040 30880
rect 3976 30796 4028 30802
rect 3976 30738 4028 30744
rect 6564 30734 6592 31282
rect 6920 31272 6972 31278
rect 6920 31214 6972 31220
rect 6932 30802 6960 31214
rect 9140 30938 9168 31758
rect 9128 30932 9180 30938
rect 9128 30874 9180 30880
rect 6920 30796 6972 30802
rect 6920 30738 6972 30744
rect 4252 30728 4304 30734
rect 4252 30670 4304 30676
rect 6552 30728 6604 30734
rect 6552 30670 6604 30676
rect 4264 30394 4292 30670
rect 4252 30388 4304 30394
rect 4252 30330 4304 30336
rect 3424 30252 3476 30258
rect 3424 30194 3476 30200
rect 4160 30184 4212 30190
rect 4160 30126 4212 30132
rect 4172 29510 4200 30126
rect 5674 29948 5982 29957
rect 5674 29946 5680 29948
rect 5736 29946 5760 29948
rect 5816 29946 5840 29948
rect 5896 29946 5920 29948
rect 5976 29946 5982 29948
rect 5736 29894 5738 29946
rect 5918 29894 5920 29946
rect 5674 29892 5680 29894
rect 5736 29892 5760 29894
rect 5816 29892 5840 29894
rect 5896 29892 5920 29894
rect 5976 29892 5982 29894
rect 5674 29883 5982 29892
rect 4160 29504 4212 29510
rect 4160 29446 4212 29452
rect 4620 29504 4672 29510
rect 4620 29446 4672 29452
rect 3240 27328 3292 27334
rect 3240 27270 3292 27276
rect 3252 26994 3280 27270
rect 3976 27056 4028 27062
rect 3976 26998 4028 27004
rect 3240 26988 3292 26994
rect 3240 26930 3292 26936
rect 3148 26376 3200 26382
rect 3148 26318 3200 26324
rect 3884 26376 3936 26382
rect 3884 26318 3936 26324
rect 2884 26206 3096 26234
rect 2884 23526 2912 26206
rect 3608 24064 3660 24070
rect 3608 24006 3660 24012
rect 3620 23730 3648 24006
rect 3608 23724 3660 23730
rect 3608 23666 3660 23672
rect 2872 23520 2924 23526
rect 2872 23462 2924 23468
rect 2780 20596 2832 20602
rect 2780 20538 2832 20544
rect 2228 18080 2280 18086
rect 2228 18022 2280 18028
rect 2240 16726 2268 18022
rect 2228 16720 2280 16726
rect 2228 16662 2280 16668
rect 2780 16448 2832 16454
rect 2780 16390 2832 16396
rect 2792 16114 2820 16390
rect 2780 16108 2832 16114
rect 2780 16050 2832 16056
rect 2044 13184 2096 13190
rect 2044 13126 2096 13132
rect 2136 12096 2188 12102
rect 2136 12038 2188 12044
rect 1952 9444 2004 9450
rect 1952 9386 2004 9392
rect 1584 6316 1636 6322
rect 1584 6258 1636 6264
rect 1492 6112 1544 6118
rect 1492 6054 1544 6060
rect 1504 5817 1532 6054
rect 1490 5808 1546 5817
rect 1490 5743 1546 5752
rect 1492 4480 1544 4486
rect 1490 4448 1492 4457
rect 1544 4448 1546 4457
rect 1490 4383 1546 4392
rect 1492 3392 1544 3398
rect 1492 3334 1544 3340
rect 1504 3097 1532 3334
rect 2148 3194 2176 12038
rect 2228 11552 2280 11558
rect 2228 11494 2280 11500
rect 2240 11286 2268 11494
rect 2228 11280 2280 11286
rect 2228 11222 2280 11228
rect 2884 9042 2912 23462
rect 3896 22778 3924 26318
rect 3988 26314 4016 26998
rect 3976 26308 4028 26314
rect 3976 26250 4028 26256
rect 3988 24206 4016 26250
rect 4344 25696 4396 25702
rect 4344 25638 4396 25644
rect 3976 24200 4028 24206
rect 3976 24142 4028 24148
rect 4160 24200 4212 24206
rect 4160 24142 4212 24148
rect 3884 22772 3936 22778
rect 3884 22714 3936 22720
rect 3896 22506 3924 22714
rect 3884 22500 3936 22506
rect 3884 22442 3936 22448
rect 3056 22432 3108 22438
rect 3056 22374 3108 22380
rect 3068 21554 3096 22374
rect 3056 21548 3108 21554
rect 3056 21490 3108 21496
rect 2964 21344 3016 21350
rect 2964 21286 3016 21292
rect 2976 20942 3004 21286
rect 2964 20936 3016 20942
rect 2964 20878 3016 20884
rect 3884 20936 3936 20942
rect 3884 20878 3936 20884
rect 3608 18624 3660 18630
rect 3608 18566 3660 18572
rect 3620 18290 3648 18566
rect 3896 18290 3924 20878
rect 4172 19310 4200 24142
rect 4160 19304 4212 19310
rect 4160 19246 4212 19252
rect 3976 19168 4028 19174
rect 3976 19110 4028 19116
rect 3988 18766 4016 19110
rect 3976 18760 4028 18766
rect 3976 18702 4028 18708
rect 3608 18284 3660 18290
rect 3608 18226 3660 18232
rect 3884 18284 3936 18290
rect 3884 18226 3936 18232
rect 3976 17604 4028 17610
rect 3976 17546 4028 17552
rect 3988 16590 4016 17546
rect 4160 16788 4212 16794
rect 4160 16730 4212 16736
rect 4172 16590 4200 16730
rect 2964 16584 3016 16590
rect 2964 16526 3016 16532
rect 3976 16584 4028 16590
rect 3976 16526 4028 16532
rect 4160 16584 4212 16590
rect 4212 16546 4292 16574
rect 4160 16526 4212 16532
rect 2976 16250 3004 16526
rect 2964 16244 3016 16250
rect 2964 16186 3016 16192
rect 3792 14408 3844 14414
rect 3792 14350 3844 14356
rect 3332 12980 3384 12986
rect 3332 12922 3384 12928
rect 3148 12844 3200 12850
rect 3148 12786 3200 12792
rect 3160 12646 3188 12786
rect 3148 12640 3200 12646
rect 3148 12582 3200 12588
rect 3160 12102 3188 12582
rect 3148 12096 3200 12102
rect 3148 12038 3200 12044
rect 3344 11694 3372 12922
rect 3608 12640 3660 12646
rect 3608 12582 3660 12588
rect 3424 12096 3476 12102
rect 3424 12038 3476 12044
rect 3436 11762 3464 12038
rect 3620 11762 3648 12582
rect 3804 12306 3832 14350
rect 3792 12300 3844 12306
rect 3792 12242 3844 12248
rect 4160 12232 4212 12238
rect 4160 12174 4212 12180
rect 4172 11898 4200 12174
rect 4160 11892 4212 11898
rect 4160 11834 4212 11840
rect 3424 11756 3476 11762
rect 3424 11698 3476 11704
rect 3608 11756 3660 11762
rect 3608 11698 3660 11704
rect 3332 11688 3384 11694
rect 3332 11630 3384 11636
rect 3344 10810 3372 11630
rect 3332 10804 3384 10810
rect 3332 10746 3384 10752
rect 3700 9444 3752 9450
rect 3700 9386 3752 9392
rect 3712 9110 3740 9386
rect 3700 9104 3752 9110
rect 3700 9046 3752 9052
rect 2872 9036 2924 9042
rect 2872 8978 2924 8984
rect 2688 8900 2740 8906
rect 2688 8842 2740 8848
rect 2700 8634 2728 8842
rect 2872 8832 2924 8838
rect 3700 8832 3752 8838
rect 2924 8780 3004 8786
rect 2872 8774 3004 8780
rect 3700 8774 3752 8780
rect 2884 8758 3004 8774
rect 2688 8628 2740 8634
rect 2688 8570 2740 8576
rect 2976 8566 3004 8758
rect 2964 8560 3016 8566
rect 2964 8502 3016 8508
rect 3712 8498 3740 8774
rect 3700 8492 3752 8498
rect 3700 8434 3752 8440
rect 3240 8288 3292 8294
rect 3240 8230 3292 8236
rect 4068 8288 4120 8294
rect 4068 8230 4120 8236
rect 3252 7886 3280 8230
rect 4080 7886 4108 8230
rect 3240 7880 3292 7886
rect 3240 7822 3292 7828
rect 3792 7880 3844 7886
rect 3792 7822 3844 7828
rect 4068 7880 4120 7886
rect 4068 7822 4120 7828
rect 3148 7812 3200 7818
rect 3148 7754 3200 7760
rect 3160 6118 3188 7754
rect 3608 7744 3660 7750
rect 3608 7686 3660 7692
rect 3620 6322 3648 7686
rect 3804 6390 3832 7822
rect 3792 6384 3844 6390
rect 3792 6326 3844 6332
rect 3608 6316 3660 6322
rect 3608 6258 3660 6264
rect 3148 6112 3200 6118
rect 3148 6054 3200 6060
rect 2872 4820 2924 4826
rect 2872 4762 2924 4768
rect 2884 4078 2912 4762
rect 3160 4622 3188 6054
rect 4264 4826 4292 16546
rect 4356 12434 4384 25638
rect 4632 24206 4660 29446
rect 5674 28860 5982 28869
rect 5674 28858 5680 28860
rect 5736 28858 5760 28860
rect 5816 28858 5840 28860
rect 5896 28858 5920 28860
rect 5976 28858 5982 28860
rect 5736 28806 5738 28858
rect 5918 28806 5920 28858
rect 5674 28804 5680 28806
rect 5736 28804 5760 28806
rect 5816 28804 5840 28806
rect 5896 28804 5920 28806
rect 5976 28804 5982 28806
rect 5674 28795 5982 28804
rect 5674 27772 5982 27781
rect 5674 27770 5680 27772
rect 5736 27770 5760 27772
rect 5816 27770 5840 27772
rect 5896 27770 5920 27772
rect 5976 27770 5982 27772
rect 5736 27718 5738 27770
rect 5918 27718 5920 27770
rect 5674 27716 5680 27718
rect 5736 27716 5760 27718
rect 5816 27716 5840 27718
rect 5896 27716 5920 27718
rect 5976 27716 5982 27718
rect 5674 27707 5982 27716
rect 6932 27470 6960 30738
rect 9128 28552 9180 28558
rect 9128 28494 9180 28500
rect 8392 28416 8444 28422
rect 8392 28358 8444 28364
rect 8404 28082 8432 28358
rect 8392 28076 8444 28082
rect 8392 28018 8444 28024
rect 8116 28008 8168 28014
rect 8116 27950 8168 27956
rect 5080 27464 5132 27470
rect 5080 27406 5132 27412
rect 5540 27464 5592 27470
rect 5540 27406 5592 27412
rect 6736 27464 6788 27470
rect 6736 27406 6788 27412
rect 6920 27464 6972 27470
rect 6920 27406 6972 27412
rect 5092 26994 5120 27406
rect 5552 27130 5580 27406
rect 5724 27396 5776 27402
rect 5724 27338 5776 27344
rect 5736 27282 5764 27338
rect 5644 27254 5764 27282
rect 6552 27328 6604 27334
rect 6552 27270 6604 27276
rect 5540 27124 5592 27130
rect 5540 27066 5592 27072
rect 5644 26994 5672 27254
rect 6564 26994 6592 27270
rect 6748 27062 6776 27406
rect 6736 27056 6788 27062
rect 6736 26998 6788 27004
rect 5080 26988 5132 26994
rect 5080 26930 5132 26936
rect 5632 26988 5684 26994
rect 5632 26930 5684 26936
rect 6552 26988 6604 26994
rect 6552 26930 6604 26936
rect 5674 26684 5982 26693
rect 5674 26682 5680 26684
rect 5736 26682 5760 26684
rect 5816 26682 5840 26684
rect 5896 26682 5920 26684
rect 5976 26682 5982 26684
rect 5736 26630 5738 26682
rect 5918 26630 5920 26682
rect 5674 26628 5680 26630
rect 5736 26628 5760 26630
rect 5816 26628 5840 26630
rect 5896 26628 5920 26630
rect 5976 26628 5982 26630
rect 5674 26619 5982 26628
rect 5674 25596 5982 25605
rect 5674 25594 5680 25596
rect 5736 25594 5760 25596
rect 5816 25594 5840 25596
rect 5896 25594 5920 25596
rect 5976 25594 5982 25596
rect 5736 25542 5738 25594
rect 5918 25542 5920 25594
rect 5674 25540 5680 25542
rect 5736 25540 5760 25542
rect 5816 25540 5840 25542
rect 5896 25540 5920 25542
rect 5976 25540 5982 25542
rect 5674 25531 5982 25540
rect 5674 24508 5982 24517
rect 5674 24506 5680 24508
rect 5736 24506 5760 24508
rect 5816 24506 5840 24508
rect 5896 24506 5920 24508
rect 5976 24506 5982 24508
rect 5736 24454 5738 24506
rect 5918 24454 5920 24506
rect 5674 24452 5680 24454
rect 5736 24452 5760 24454
rect 5816 24452 5840 24454
rect 5896 24452 5920 24454
rect 5976 24452 5982 24454
rect 5674 24443 5982 24452
rect 4620 24200 4672 24206
rect 4620 24142 4672 24148
rect 5674 23420 5982 23429
rect 5674 23418 5680 23420
rect 5736 23418 5760 23420
rect 5816 23418 5840 23420
rect 5896 23418 5920 23420
rect 5976 23418 5982 23420
rect 5736 23366 5738 23418
rect 5918 23366 5920 23418
rect 5674 23364 5680 23366
rect 5736 23364 5760 23366
rect 5816 23364 5840 23366
rect 5896 23364 5920 23366
rect 5976 23364 5982 23366
rect 5674 23355 5982 23364
rect 6932 23186 6960 27406
rect 8128 27402 8156 27950
rect 8392 27872 8444 27878
rect 8392 27814 8444 27820
rect 8404 27606 8432 27814
rect 9140 27674 9168 28494
rect 9128 27668 9180 27674
rect 9128 27610 9180 27616
rect 8392 27600 8444 27606
rect 8392 27542 8444 27548
rect 7380 27396 7432 27402
rect 7380 27338 7432 27344
rect 8116 27396 8168 27402
rect 8116 27338 8168 27344
rect 7392 26450 7420 27338
rect 7840 26988 7892 26994
rect 7840 26930 7892 26936
rect 7656 26784 7708 26790
rect 7656 26726 7708 26732
rect 7380 26444 7432 26450
rect 7380 26386 7432 26392
rect 7668 26382 7696 26726
rect 7656 26376 7708 26382
rect 7656 26318 7708 26324
rect 7852 26042 7880 26930
rect 8128 26234 8156 27338
rect 8404 26586 8432 27542
rect 9220 27464 9272 27470
rect 9220 27406 9272 27412
rect 8392 26580 8444 26586
rect 8392 26522 8444 26528
rect 8036 26206 8156 26234
rect 7840 26036 7892 26042
rect 7840 25978 7892 25984
rect 7380 25832 7432 25838
rect 7380 25774 7432 25780
rect 6920 23180 6972 23186
rect 6920 23122 6972 23128
rect 5448 23112 5500 23118
rect 5448 23054 5500 23060
rect 5460 22642 5488 23054
rect 6000 22976 6052 22982
rect 6000 22918 6052 22924
rect 4620 22636 4672 22642
rect 4620 22578 4672 22584
rect 5448 22636 5500 22642
rect 5448 22578 5500 22584
rect 4632 19378 4660 22578
rect 5674 22332 5982 22341
rect 5674 22330 5680 22332
rect 5736 22330 5760 22332
rect 5816 22330 5840 22332
rect 5896 22330 5920 22332
rect 5976 22330 5982 22332
rect 5736 22278 5738 22330
rect 5918 22278 5920 22330
rect 5674 22276 5680 22278
rect 5736 22276 5760 22278
rect 5816 22276 5840 22278
rect 5896 22276 5920 22278
rect 5976 22276 5982 22278
rect 5674 22267 5982 22276
rect 6012 22030 6040 22918
rect 7392 22574 7420 25774
rect 8036 23866 8064 26206
rect 8404 23866 8432 26522
rect 9232 25906 9260 27406
rect 9220 25900 9272 25906
rect 9220 25842 9272 25848
rect 9232 24206 9260 25842
rect 8944 24200 8996 24206
rect 8944 24142 8996 24148
rect 9220 24200 9272 24206
rect 9220 24142 9272 24148
rect 8024 23860 8076 23866
rect 8024 23802 8076 23808
rect 8392 23860 8444 23866
rect 8392 23802 8444 23808
rect 8956 23186 8984 24142
rect 8944 23180 8996 23186
rect 8944 23122 8996 23128
rect 9036 23112 9088 23118
rect 9036 23054 9088 23060
rect 7380 22568 7432 22574
rect 7380 22510 7432 22516
rect 6920 22432 6972 22438
rect 6920 22374 6972 22380
rect 6932 22030 6960 22374
rect 6000 22024 6052 22030
rect 6000 21966 6052 21972
rect 6920 22024 6972 22030
rect 6920 21966 6972 21972
rect 6000 21888 6052 21894
rect 6000 21830 6052 21836
rect 7012 21888 7064 21894
rect 7012 21830 7064 21836
rect 5674 21244 5982 21253
rect 5674 21242 5680 21244
rect 5736 21242 5760 21244
rect 5816 21242 5840 21244
rect 5896 21242 5920 21244
rect 5976 21242 5982 21244
rect 5736 21190 5738 21242
rect 5918 21190 5920 21242
rect 5674 21188 5680 21190
rect 5736 21188 5760 21190
rect 5816 21188 5840 21190
rect 5896 21188 5920 21190
rect 5976 21188 5982 21190
rect 5674 21179 5982 21188
rect 6012 20942 6040 21830
rect 7024 20942 7052 21830
rect 6000 20936 6052 20942
rect 6000 20878 6052 20884
rect 6644 20936 6696 20942
rect 6644 20878 6696 20884
rect 7012 20936 7064 20942
rect 7012 20878 7064 20884
rect 5674 20156 5982 20165
rect 5674 20154 5680 20156
rect 5736 20154 5760 20156
rect 5816 20154 5840 20156
rect 5896 20154 5920 20156
rect 5976 20154 5982 20156
rect 5736 20102 5738 20154
rect 5918 20102 5920 20154
rect 5674 20100 5680 20102
rect 5736 20100 5760 20102
rect 5816 20100 5840 20102
rect 5896 20100 5920 20102
rect 5976 20100 5982 20102
rect 5674 20091 5982 20100
rect 6656 20058 6684 20878
rect 6736 20800 6788 20806
rect 6736 20742 6788 20748
rect 6644 20052 6696 20058
rect 6644 19994 6696 20000
rect 6276 19848 6328 19854
rect 6276 19790 6328 19796
rect 4620 19372 4672 19378
rect 4620 19314 4672 19320
rect 4632 18222 4660 19314
rect 5674 19068 5982 19077
rect 5674 19066 5680 19068
rect 5736 19066 5760 19068
rect 5816 19066 5840 19068
rect 5896 19066 5920 19068
rect 5976 19066 5982 19068
rect 5736 19014 5738 19066
rect 5918 19014 5920 19066
rect 5674 19012 5680 19014
rect 5736 19012 5760 19014
rect 5816 19012 5840 19014
rect 5896 19012 5920 19014
rect 5976 19012 5982 19014
rect 5674 19003 5982 19012
rect 6288 18766 6316 19790
rect 6748 18970 6776 20742
rect 7104 19372 7156 19378
rect 7104 19314 7156 19320
rect 7012 19168 7064 19174
rect 7012 19110 7064 19116
rect 6736 18964 6788 18970
rect 6736 18906 6788 18912
rect 7024 18766 7052 19110
rect 6276 18760 6328 18766
rect 6276 18702 6328 18708
rect 7012 18760 7064 18766
rect 7012 18702 7064 18708
rect 4620 18216 4672 18222
rect 4620 18158 4672 18164
rect 4632 17746 4660 18158
rect 5674 17980 5982 17989
rect 5674 17978 5680 17980
rect 5736 17978 5760 17980
rect 5816 17978 5840 17980
rect 5896 17978 5920 17980
rect 5976 17978 5982 17980
rect 5736 17926 5738 17978
rect 5918 17926 5920 17978
rect 5674 17924 5680 17926
rect 5736 17924 5760 17926
rect 5816 17924 5840 17926
rect 5896 17924 5920 17926
rect 5976 17924 5982 17926
rect 5674 17915 5982 17924
rect 4620 17740 4672 17746
rect 4620 17682 4672 17688
rect 5674 16892 5982 16901
rect 5674 16890 5680 16892
rect 5736 16890 5760 16892
rect 5816 16890 5840 16892
rect 5896 16890 5920 16892
rect 5976 16890 5982 16892
rect 5736 16838 5738 16890
rect 5918 16838 5920 16890
rect 5674 16836 5680 16838
rect 5736 16836 5760 16838
rect 5816 16836 5840 16838
rect 5896 16836 5920 16838
rect 5976 16836 5982 16838
rect 5674 16827 5982 16836
rect 6288 16590 6316 18702
rect 7116 18426 7144 19314
rect 7104 18420 7156 18426
rect 7104 18362 7156 18368
rect 8300 18352 8352 18358
rect 8300 18294 8352 18300
rect 7288 18216 7340 18222
rect 7288 18158 7340 18164
rect 7300 17542 7328 18158
rect 8208 17672 8260 17678
rect 8208 17614 8260 17620
rect 7288 17536 7340 17542
rect 7288 17478 7340 17484
rect 8220 16658 8248 17614
rect 6920 16652 6972 16658
rect 6920 16594 6972 16600
rect 8208 16652 8260 16658
rect 8208 16594 8260 16600
rect 6276 16584 6328 16590
rect 6276 16526 6328 16532
rect 6932 16522 6960 16594
rect 6920 16516 6972 16522
rect 6920 16458 6972 16464
rect 5674 15804 5982 15813
rect 5674 15802 5680 15804
rect 5736 15802 5760 15804
rect 5816 15802 5840 15804
rect 5896 15802 5920 15804
rect 5976 15802 5982 15804
rect 5736 15750 5738 15802
rect 5918 15750 5920 15802
rect 5674 15748 5680 15750
rect 5736 15748 5760 15750
rect 5816 15748 5840 15750
rect 5896 15748 5920 15750
rect 5976 15748 5982 15750
rect 5674 15739 5982 15748
rect 5674 14716 5982 14725
rect 5674 14714 5680 14716
rect 5736 14714 5760 14716
rect 5816 14714 5840 14716
rect 5896 14714 5920 14716
rect 5976 14714 5982 14716
rect 5736 14662 5738 14714
rect 5918 14662 5920 14714
rect 5674 14660 5680 14662
rect 5736 14660 5760 14662
rect 5816 14660 5840 14662
rect 5896 14660 5920 14662
rect 5976 14660 5982 14662
rect 5674 14651 5982 14660
rect 6000 14340 6052 14346
rect 6000 14282 6052 14288
rect 5674 13628 5982 13637
rect 5674 13626 5680 13628
rect 5736 13626 5760 13628
rect 5816 13626 5840 13628
rect 5896 13626 5920 13628
rect 5976 13626 5982 13628
rect 5736 13574 5738 13626
rect 5918 13574 5920 13626
rect 5674 13572 5680 13574
rect 5736 13572 5760 13574
rect 5816 13572 5840 13574
rect 5896 13572 5920 13574
rect 5976 13572 5982 13574
rect 5674 13563 5982 13572
rect 6012 13530 6040 14282
rect 6000 13524 6052 13530
rect 6000 13466 6052 13472
rect 5674 12540 5982 12549
rect 5674 12538 5680 12540
rect 5736 12538 5760 12540
rect 5816 12538 5840 12540
rect 5896 12538 5920 12540
rect 5976 12538 5982 12540
rect 5736 12486 5738 12538
rect 5918 12486 5920 12538
rect 5674 12484 5680 12486
rect 5736 12484 5760 12486
rect 5816 12484 5840 12486
rect 5896 12484 5920 12486
rect 5976 12484 5982 12486
rect 5674 12475 5982 12484
rect 5540 12436 5592 12442
rect 4356 12406 4476 12434
rect 4448 8362 4476 12406
rect 5540 12378 5592 12384
rect 5172 12164 5224 12170
rect 5172 12106 5224 12112
rect 5184 11898 5212 12106
rect 5172 11892 5224 11898
rect 5172 11834 5224 11840
rect 4896 10464 4948 10470
rect 4896 10406 4948 10412
rect 4908 10062 4936 10406
rect 4896 10056 4948 10062
rect 4896 9998 4948 10004
rect 4712 9920 4764 9926
rect 4712 9862 4764 9868
rect 4436 8356 4488 8362
rect 4436 8298 4488 8304
rect 4252 4820 4304 4826
rect 4252 4762 4304 4768
rect 3148 4616 3200 4622
rect 3148 4558 3200 4564
rect 3160 4282 3188 4558
rect 3148 4276 3200 4282
rect 3148 4218 3200 4224
rect 4068 4276 4120 4282
rect 4068 4218 4120 4224
rect 2872 4072 2924 4078
rect 2872 4014 2924 4020
rect 4080 4026 4108 4218
rect 4080 3998 4292 4026
rect 4264 3942 4292 3998
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 4252 3936 4304 3942
rect 4252 3878 4304 3884
rect 2884 3534 2912 3878
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 2136 3188 2188 3194
rect 2136 3130 2188 3136
rect 1490 3088 1546 3097
rect 1490 3023 1546 3032
rect 2148 2514 2176 3130
rect 2228 2848 2280 2854
rect 2228 2790 2280 2796
rect 2136 2508 2188 2514
rect 2136 2450 2188 2456
rect 2240 2446 2268 2790
rect 4448 2514 4476 8298
rect 4724 4146 4752 9862
rect 4988 9376 5040 9382
rect 4988 9318 5040 9324
rect 5000 9042 5028 9318
rect 4988 9036 5040 9042
rect 4988 8978 5040 8984
rect 5000 8634 5028 8978
rect 4988 8628 5040 8634
rect 4988 8570 5040 8576
rect 5552 4706 5580 12378
rect 6276 11552 6328 11558
rect 6276 11494 6328 11500
rect 5674 11452 5982 11461
rect 5674 11450 5680 11452
rect 5736 11450 5760 11452
rect 5816 11450 5840 11452
rect 5896 11450 5920 11452
rect 5976 11450 5982 11452
rect 5736 11398 5738 11450
rect 5918 11398 5920 11450
rect 5674 11396 5680 11398
rect 5736 11396 5760 11398
rect 5816 11396 5840 11398
rect 5896 11396 5920 11398
rect 5976 11396 5982 11398
rect 5674 11387 5982 11396
rect 5674 10364 5982 10373
rect 5674 10362 5680 10364
rect 5736 10362 5760 10364
rect 5816 10362 5840 10364
rect 5896 10362 5920 10364
rect 5976 10362 5982 10364
rect 5736 10310 5738 10362
rect 5918 10310 5920 10362
rect 5674 10308 5680 10310
rect 5736 10308 5760 10310
rect 5816 10308 5840 10310
rect 5896 10308 5920 10310
rect 5976 10308 5982 10310
rect 5674 10299 5982 10308
rect 5674 9276 5982 9285
rect 5674 9274 5680 9276
rect 5736 9274 5760 9276
rect 5816 9274 5840 9276
rect 5896 9274 5920 9276
rect 5976 9274 5982 9276
rect 5736 9222 5738 9274
rect 5918 9222 5920 9274
rect 5674 9220 5680 9222
rect 5736 9220 5760 9222
rect 5816 9220 5840 9222
rect 5896 9220 5920 9222
rect 5976 9220 5982 9222
rect 5674 9211 5982 9220
rect 6184 8832 6236 8838
rect 6184 8774 6236 8780
rect 5674 8188 5982 8197
rect 5674 8186 5680 8188
rect 5736 8186 5760 8188
rect 5816 8186 5840 8188
rect 5896 8186 5920 8188
rect 5976 8186 5982 8188
rect 5736 8134 5738 8186
rect 5918 8134 5920 8186
rect 5674 8132 5680 8134
rect 5736 8132 5760 8134
rect 5816 8132 5840 8134
rect 5896 8132 5920 8134
rect 5976 8132 5982 8134
rect 5674 8123 5982 8132
rect 6092 7744 6144 7750
rect 6092 7686 6144 7692
rect 5674 7100 5982 7109
rect 5674 7098 5680 7100
rect 5736 7098 5760 7100
rect 5816 7098 5840 7100
rect 5896 7098 5920 7100
rect 5976 7098 5982 7100
rect 5736 7046 5738 7098
rect 5918 7046 5920 7098
rect 5674 7044 5680 7046
rect 5736 7044 5760 7046
rect 5816 7044 5840 7046
rect 5896 7044 5920 7046
rect 5976 7044 5982 7046
rect 5674 7035 5982 7044
rect 5674 6012 5982 6021
rect 5674 6010 5680 6012
rect 5736 6010 5760 6012
rect 5816 6010 5840 6012
rect 5896 6010 5920 6012
rect 5976 6010 5982 6012
rect 5736 5958 5738 6010
rect 5918 5958 5920 6010
rect 5674 5956 5680 5958
rect 5736 5956 5760 5958
rect 5816 5956 5840 5958
rect 5896 5956 5920 5958
rect 5976 5956 5982 5958
rect 5674 5947 5982 5956
rect 5674 4924 5982 4933
rect 5674 4922 5680 4924
rect 5736 4922 5760 4924
rect 5816 4922 5840 4924
rect 5896 4922 5920 4924
rect 5976 4922 5982 4924
rect 5736 4870 5738 4922
rect 5918 4870 5920 4922
rect 5674 4868 5680 4870
rect 5736 4868 5760 4870
rect 5816 4868 5840 4870
rect 5896 4868 5920 4870
rect 5976 4868 5982 4870
rect 5674 4859 5982 4868
rect 5552 4678 5672 4706
rect 5540 4480 5592 4486
rect 5540 4422 5592 4428
rect 5552 4146 5580 4422
rect 4712 4140 4764 4146
rect 4712 4082 4764 4088
rect 5540 4140 5592 4146
rect 5540 4082 5592 4088
rect 5644 4026 5672 4678
rect 6104 4622 6132 7686
rect 6196 6322 6224 8774
rect 6184 6316 6236 6322
rect 6184 6258 6236 6264
rect 6196 5710 6224 6258
rect 6184 5704 6236 5710
rect 6184 5646 6236 5652
rect 6196 5234 6224 5646
rect 6184 5228 6236 5234
rect 6184 5170 6236 5176
rect 6092 4616 6144 4622
rect 6092 4558 6144 4564
rect 5552 3998 5672 4026
rect 5552 3194 5580 3998
rect 5674 3836 5982 3845
rect 5674 3834 5680 3836
rect 5736 3834 5760 3836
rect 5816 3834 5840 3836
rect 5896 3834 5920 3836
rect 5976 3834 5982 3836
rect 5736 3782 5738 3834
rect 5918 3782 5920 3834
rect 5674 3780 5680 3782
rect 5736 3780 5760 3782
rect 5816 3780 5840 3782
rect 5896 3780 5920 3782
rect 5976 3780 5982 3782
rect 5674 3771 5982 3780
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 4436 2508 4488 2514
rect 4436 2450 4488 2456
rect 5552 2446 5580 3130
rect 5674 2748 5982 2757
rect 5674 2746 5680 2748
rect 5736 2746 5760 2748
rect 5816 2746 5840 2748
rect 5896 2746 5920 2748
rect 5976 2746 5982 2748
rect 5736 2694 5738 2746
rect 5918 2694 5920 2746
rect 5674 2692 5680 2694
rect 5736 2692 5760 2694
rect 5816 2692 5840 2694
rect 5896 2692 5920 2694
rect 5976 2692 5982 2694
rect 5674 2683 5982 2692
rect 6288 2446 6316 11494
rect 6932 9450 6960 16458
rect 7104 16448 7156 16454
rect 7104 16390 7156 16396
rect 7116 10742 7144 16390
rect 8312 16182 8340 18294
rect 8852 17536 8904 17542
rect 8852 17478 8904 17484
rect 8864 16574 8892 17478
rect 9048 16794 9076 23054
rect 9416 19378 9444 33254
rect 12532 32904 12584 32910
rect 12532 32846 12584 32852
rect 10398 32668 10706 32677
rect 10398 32666 10404 32668
rect 10460 32666 10484 32668
rect 10540 32666 10564 32668
rect 10620 32666 10644 32668
rect 10700 32666 10706 32668
rect 10460 32614 10462 32666
rect 10642 32614 10644 32666
rect 10398 32612 10404 32614
rect 10460 32612 10484 32614
rect 10540 32612 10564 32614
rect 10620 32612 10644 32614
rect 10700 32612 10706 32614
rect 10398 32603 10706 32612
rect 11796 32428 11848 32434
rect 11796 32370 11848 32376
rect 10876 32224 10928 32230
rect 10876 32166 10928 32172
rect 10398 31580 10706 31589
rect 10398 31578 10404 31580
rect 10460 31578 10484 31580
rect 10540 31578 10564 31580
rect 10620 31578 10644 31580
rect 10700 31578 10706 31580
rect 10460 31526 10462 31578
rect 10642 31526 10644 31578
rect 10398 31524 10404 31526
rect 10460 31524 10484 31526
rect 10540 31524 10564 31526
rect 10620 31524 10644 31526
rect 10700 31524 10706 31526
rect 10398 31515 10706 31524
rect 9864 30728 9916 30734
rect 9864 30670 9916 30676
rect 9876 30598 9904 30670
rect 9864 30592 9916 30598
rect 9864 30534 9916 30540
rect 9876 27334 9904 30534
rect 10398 30492 10706 30501
rect 10398 30490 10404 30492
rect 10460 30490 10484 30492
rect 10540 30490 10564 30492
rect 10620 30490 10644 30492
rect 10700 30490 10706 30492
rect 10460 30438 10462 30490
rect 10642 30438 10644 30490
rect 10398 30436 10404 30438
rect 10460 30436 10484 30438
rect 10540 30436 10564 30438
rect 10620 30436 10644 30438
rect 10700 30436 10706 30438
rect 10398 30427 10706 30436
rect 10398 29404 10706 29413
rect 10398 29402 10404 29404
rect 10460 29402 10484 29404
rect 10540 29402 10564 29404
rect 10620 29402 10644 29404
rect 10700 29402 10706 29404
rect 10460 29350 10462 29402
rect 10642 29350 10644 29402
rect 10398 29348 10404 29350
rect 10460 29348 10484 29350
rect 10540 29348 10564 29350
rect 10620 29348 10644 29350
rect 10700 29348 10706 29350
rect 10398 29339 10706 29348
rect 10398 28316 10706 28325
rect 10398 28314 10404 28316
rect 10460 28314 10484 28316
rect 10540 28314 10564 28316
rect 10620 28314 10644 28316
rect 10700 28314 10706 28316
rect 10460 28262 10462 28314
rect 10642 28262 10644 28314
rect 10398 28260 10404 28262
rect 10460 28260 10484 28262
rect 10540 28260 10564 28262
rect 10620 28260 10644 28262
rect 10700 28260 10706 28262
rect 10398 28251 10706 28260
rect 9864 27328 9916 27334
rect 9864 27270 9916 27276
rect 9876 26790 9904 27270
rect 10398 27228 10706 27237
rect 10398 27226 10404 27228
rect 10460 27226 10484 27228
rect 10540 27226 10564 27228
rect 10620 27226 10644 27228
rect 10700 27226 10706 27228
rect 10460 27174 10462 27226
rect 10642 27174 10644 27226
rect 10398 27172 10404 27174
rect 10460 27172 10484 27174
rect 10540 27172 10564 27174
rect 10620 27172 10644 27174
rect 10700 27172 10706 27174
rect 10398 27163 10706 27172
rect 9864 26784 9916 26790
rect 9864 26726 9916 26732
rect 10398 26140 10706 26149
rect 10398 26138 10404 26140
rect 10460 26138 10484 26140
rect 10540 26138 10564 26140
rect 10620 26138 10644 26140
rect 10700 26138 10706 26140
rect 10460 26086 10462 26138
rect 10642 26086 10644 26138
rect 10398 26084 10404 26086
rect 10460 26084 10484 26086
rect 10540 26084 10564 26086
rect 10620 26084 10644 26086
rect 10700 26084 10706 26086
rect 10398 26075 10706 26084
rect 10398 25052 10706 25061
rect 10398 25050 10404 25052
rect 10460 25050 10484 25052
rect 10540 25050 10564 25052
rect 10620 25050 10644 25052
rect 10700 25050 10706 25052
rect 10460 24998 10462 25050
rect 10642 24998 10644 25050
rect 10398 24996 10404 24998
rect 10460 24996 10484 24998
rect 10540 24996 10564 24998
rect 10620 24996 10644 24998
rect 10700 24996 10706 24998
rect 10398 24987 10706 24996
rect 10398 23964 10706 23973
rect 10398 23962 10404 23964
rect 10460 23962 10484 23964
rect 10540 23962 10564 23964
rect 10620 23962 10644 23964
rect 10700 23962 10706 23964
rect 10460 23910 10462 23962
rect 10642 23910 10644 23962
rect 10398 23908 10404 23910
rect 10460 23908 10484 23910
rect 10540 23908 10564 23910
rect 10620 23908 10644 23910
rect 10700 23908 10706 23910
rect 10398 23899 10706 23908
rect 9496 23792 9548 23798
rect 9496 23734 9548 23740
rect 9508 23662 9536 23734
rect 9864 23724 9916 23730
rect 9864 23666 9916 23672
rect 9496 23656 9548 23662
rect 9496 23598 9548 23604
rect 9508 22778 9536 23598
rect 9876 23322 9904 23666
rect 9956 23520 10008 23526
rect 9956 23462 10008 23468
rect 9864 23316 9916 23322
rect 9864 23258 9916 23264
rect 9588 23180 9640 23186
rect 9588 23122 9640 23128
rect 9496 22772 9548 22778
rect 9496 22714 9548 22720
rect 9600 20346 9628 23122
rect 9968 23050 9996 23462
rect 9956 23044 10008 23050
rect 9956 22986 10008 22992
rect 10398 22876 10706 22885
rect 10398 22874 10404 22876
rect 10460 22874 10484 22876
rect 10540 22874 10564 22876
rect 10620 22874 10644 22876
rect 10700 22874 10706 22876
rect 10460 22822 10462 22874
rect 10642 22822 10644 22874
rect 10398 22820 10404 22822
rect 10460 22820 10484 22822
rect 10540 22820 10564 22822
rect 10620 22820 10644 22822
rect 10700 22820 10706 22822
rect 10398 22811 10706 22820
rect 10140 22636 10192 22642
rect 10140 22578 10192 22584
rect 10152 22234 10180 22578
rect 10140 22228 10192 22234
rect 10140 22170 10192 22176
rect 10048 22024 10100 22030
rect 10048 21966 10100 21972
rect 9600 20318 9720 20346
rect 9588 20256 9640 20262
rect 9588 20198 9640 20204
rect 9404 19372 9456 19378
rect 9404 19314 9456 19320
rect 9128 18216 9180 18222
rect 9128 18158 9180 18164
rect 9036 16788 9088 16794
rect 9036 16730 9088 16736
rect 8864 16546 8984 16574
rect 8300 16176 8352 16182
rect 8300 16118 8352 16124
rect 8852 15972 8904 15978
rect 8852 15914 8904 15920
rect 8392 15632 8444 15638
rect 8392 15574 8444 15580
rect 7748 14340 7800 14346
rect 7748 14282 7800 14288
rect 7196 14272 7248 14278
rect 7196 14214 7248 14220
rect 7104 10736 7156 10742
rect 7104 10678 7156 10684
rect 6920 9444 6972 9450
rect 6920 9386 6972 9392
rect 6644 9376 6696 9382
rect 6644 9318 6696 9324
rect 6656 8974 6684 9318
rect 6644 8968 6696 8974
rect 6644 8910 6696 8916
rect 6932 8616 6960 9386
rect 7012 8628 7064 8634
rect 6932 8588 7012 8616
rect 7012 8570 7064 8576
rect 7116 8566 7144 10678
rect 7104 8560 7156 8566
rect 7104 8502 7156 8508
rect 6920 8356 6972 8362
rect 6920 8298 6972 8304
rect 6932 6798 6960 8298
rect 7116 7750 7144 8502
rect 7104 7744 7156 7750
rect 7104 7686 7156 7692
rect 6920 6792 6972 6798
rect 6920 6734 6972 6740
rect 6644 6656 6696 6662
rect 6644 6598 6696 6604
rect 6368 5568 6420 5574
rect 6368 5510 6420 5516
rect 6380 4146 6408 5510
rect 6656 5234 6684 6598
rect 6644 5228 6696 5234
rect 6644 5170 6696 5176
rect 6368 4140 6420 4146
rect 6368 4082 6420 4088
rect 7208 2446 7236 14214
rect 7760 14074 7788 14282
rect 7748 14068 7800 14074
rect 7748 14010 7800 14016
rect 7288 13320 7340 13326
rect 7288 13262 7340 13268
rect 7380 13320 7432 13326
rect 7380 13262 7432 13268
rect 7300 12306 7328 13262
rect 7288 12300 7340 12306
rect 7288 12242 7340 12248
rect 7392 10470 7420 13262
rect 7380 10464 7432 10470
rect 7380 10406 7432 10412
rect 7380 8832 7432 8838
rect 7380 8774 7432 8780
rect 7392 8566 7420 8774
rect 7380 8560 7432 8566
rect 7380 8502 7432 8508
rect 7288 8084 7340 8090
rect 7288 8026 7340 8032
rect 7300 7206 7328 8026
rect 7392 7818 7420 8502
rect 7748 8356 7800 8362
rect 7748 8298 7800 8304
rect 7564 8288 7616 8294
rect 7564 8230 7616 8236
rect 7380 7812 7432 7818
rect 7380 7754 7432 7760
rect 7392 7546 7420 7754
rect 7576 7750 7604 8230
rect 7564 7744 7616 7750
rect 7564 7686 7616 7692
rect 7380 7540 7432 7546
rect 7380 7482 7432 7488
rect 7288 7200 7340 7206
rect 7288 7142 7340 7148
rect 7300 5914 7328 7142
rect 7576 6934 7604 7686
rect 7564 6928 7616 6934
rect 7564 6870 7616 6876
rect 7288 5908 7340 5914
rect 7288 5850 7340 5856
rect 7472 5024 7524 5030
rect 7472 4966 7524 4972
rect 7484 4282 7512 4966
rect 7760 4622 7788 8298
rect 7748 4616 7800 4622
rect 7748 4558 7800 4564
rect 7564 4480 7616 4486
rect 7564 4422 7616 4428
rect 7472 4276 7524 4282
rect 7472 4218 7524 4224
rect 7484 3942 7512 4218
rect 7576 4146 7604 4422
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7472 3936 7524 3942
rect 7472 3878 7524 3884
rect 8404 2446 8432 15574
rect 8864 15434 8892 15914
rect 8852 15428 8904 15434
rect 8852 15370 8904 15376
rect 8864 14822 8892 15370
rect 8852 14816 8904 14822
rect 8852 14758 8904 14764
rect 8864 13530 8892 14758
rect 8852 13524 8904 13530
rect 8852 13466 8904 13472
rect 8864 12442 8892 13466
rect 8956 13190 8984 16546
rect 9036 15904 9088 15910
rect 9036 15846 9088 15852
rect 9048 14482 9076 15846
rect 9036 14476 9088 14482
rect 9036 14418 9088 14424
rect 8944 13184 8996 13190
rect 8944 13126 8996 13132
rect 8852 12436 8904 12442
rect 8852 12378 8904 12384
rect 8852 8832 8904 8838
rect 8852 8774 8904 8780
rect 8864 8634 8892 8774
rect 8852 8628 8904 8634
rect 8852 8570 8904 8576
rect 9048 7954 9076 14418
rect 9140 11898 9168 18158
rect 9416 16726 9444 19314
rect 9496 18828 9548 18834
rect 9496 18770 9548 18776
rect 9404 16720 9456 16726
rect 9404 16662 9456 16668
rect 9404 16108 9456 16114
rect 9404 16050 9456 16056
rect 9416 15638 9444 16050
rect 9508 15910 9536 18770
rect 9600 18358 9628 20198
rect 9692 19854 9720 20318
rect 9680 19848 9732 19854
rect 9680 19790 9732 19796
rect 9588 18352 9640 18358
rect 9588 18294 9640 18300
rect 9692 16794 9720 19790
rect 10060 18970 10088 21966
rect 10398 21788 10706 21797
rect 10398 21786 10404 21788
rect 10460 21786 10484 21788
rect 10540 21786 10564 21788
rect 10620 21786 10644 21788
rect 10700 21786 10706 21788
rect 10460 21734 10462 21786
rect 10642 21734 10644 21786
rect 10398 21732 10404 21734
rect 10460 21732 10484 21734
rect 10540 21732 10564 21734
rect 10620 21732 10644 21734
rect 10700 21732 10706 21734
rect 10398 21723 10706 21732
rect 10398 20700 10706 20709
rect 10398 20698 10404 20700
rect 10460 20698 10484 20700
rect 10540 20698 10564 20700
rect 10620 20698 10644 20700
rect 10700 20698 10706 20700
rect 10460 20646 10462 20698
rect 10642 20646 10644 20698
rect 10398 20644 10404 20646
rect 10460 20644 10484 20646
rect 10540 20644 10564 20646
rect 10620 20644 10644 20646
rect 10700 20644 10706 20646
rect 10398 20635 10706 20644
rect 10398 19612 10706 19621
rect 10398 19610 10404 19612
rect 10460 19610 10484 19612
rect 10540 19610 10564 19612
rect 10620 19610 10644 19612
rect 10700 19610 10706 19612
rect 10460 19558 10462 19610
rect 10642 19558 10644 19610
rect 10398 19556 10404 19558
rect 10460 19556 10484 19558
rect 10540 19556 10564 19558
rect 10620 19556 10644 19558
rect 10700 19556 10706 19558
rect 10398 19547 10706 19556
rect 10048 18964 10100 18970
rect 10048 18906 10100 18912
rect 9864 18760 9916 18766
rect 9864 18702 9916 18708
rect 9876 17882 9904 18702
rect 10398 18524 10706 18533
rect 10398 18522 10404 18524
rect 10460 18522 10484 18524
rect 10540 18522 10564 18524
rect 10620 18522 10644 18524
rect 10700 18522 10706 18524
rect 10460 18470 10462 18522
rect 10642 18470 10644 18522
rect 10398 18468 10404 18470
rect 10460 18468 10484 18470
rect 10540 18468 10564 18470
rect 10620 18468 10644 18470
rect 10700 18468 10706 18470
rect 10398 18459 10706 18468
rect 10888 18222 10916 32166
rect 11520 31952 11572 31958
rect 11520 31894 11572 31900
rect 11532 29850 11560 31894
rect 11704 31340 11756 31346
rect 11704 31282 11756 31288
rect 11716 30394 11744 31282
rect 11808 30666 11836 32370
rect 12544 31890 12572 32846
rect 12900 32564 12952 32570
rect 12900 32506 12952 32512
rect 12912 32230 12940 32506
rect 12900 32224 12952 32230
rect 12900 32166 12952 32172
rect 12532 31884 12584 31890
rect 12532 31826 12584 31832
rect 12256 31816 12308 31822
rect 12256 31758 12308 31764
rect 12268 31482 12296 31758
rect 12544 31754 12572 31826
rect 12544 31726 12664 31754
rect 12256 31476 12308 31482
rect 12256 31418 12308 31424
rect 11796 30660 11848 30666
rect 11796 30602 11848 30608
rect 11704 30388 11756 30394
rect 11704 30330 11756 30336
rect 11520 29844 11572 29850
rect 11520 29786 11572 29792
rect 11808 29170 11836 30602
rect 12440 30252 12492 30258
rect 12440 30194 12492 30200
rect 12452 30054 12480 30194
rect 12440 30048 12492 30054
rect 12440 29990 12492 29996
rect 11796 29164 11848 29170
rect 11796 29106 11848 29112
rect 12452 29102 12480 29990
rect 12636 29646 12664 31726
rect 12716 30796 12768 30802
rect 12716 30738 12768 30744
rect 12532 29640 12584 29646
rect 12532 29582 12584 29588
rect 12624 29640 12676 29646
rect 12624 29582 12676 29588
rect 12544 29306 12572 29582
rect 12532 29300 12584 29306
rect 12532 29242 12584 29248
rect 12440 29096 12492 29102
rect 12440 29038 12492 29044
rect 12452 28626 12480 29038
rect 12440 28620 12492 28626
rect 12440 28562 12492 28568
rect 12256 28552 12308 28558
rect 12256 28494 12308 28500
rect 12268 27946 12296 28494
rect 12636 28422 12664 29582
rect 12624 28416 12676 28422
rect 12624 28358 12676 28364
rect 12256 27940 12308 27946
rect 12256 27882 12308 27888
rect 12164 26240 12216 26246
rect 12164 26182 12216 26188
rect 12176 25906 12204 26182
rect 12164 25900 12216 25906
rect 12164 25842 12216 25848
rect 11704 25832 11756 25838
rect 11704 25774 11756 25780
rect 11716 23118 11744 25774
rect 12268 23526 12296 27882
rect 12348 26376 12400 26382
rect 12348 26318 12400 26324
rect 12360 25498 12388 26318
rect 12440 25696 12492 25702
rect 12440 25638 12492 25644
rect 12348 25492 12400 25498
rect 12348 25434 12400 25440
rect 12452 25242 12480 25638
rect 12728 25362 12756 30738
rect 12716 25356 12768 25362
rect 12716 25298 12768 25304
rect 12360 25214 12480 25242
rect 12256 23520 12308 23526
rect 12256 23462 12308 23468
rect 11704 23112 11756 23118
rect 11704 23054 11756 23060
rect 11716 22234 11744 23054
rect 11704 22228 11756 22234
rect 11704 22170 11756 22176
rect 12072 21956 12124 21962
rect 12072 21898 12124 21904
rect 11704 19780 11756 19786
rect 11704 19722 11756 19728
rect 11716 19514 11744 19722
rect 11704 19508 11756 19514
rect 11704 19450 11756 19456
rect 11336 19372 11388 19378
rect 11336 19314 11388 19320
rect 11348 18698 11376 19314
rect 11152 18692 11204 18698
rect 11152 18634 11204 18640
rect 11336 18692 11388 18698
rect 11336 18634 11388 18640
rect 11164 18358 11192 18634
rect 11152 18352 11204 18358
rect 11152 18294 11204 18300
rect 10876 18216 10928 18222
rect 10876 18158 10928 18164
rect 9864 17876 9916 17882
rect 9864 17818 9916 17824
rect 10968 17604 11020 17610
rect 10968 17546 11020 17552
rect 10398 17436 10706 17445
rect 10398 17434 10404 17436
rect 10460 17434 10484 17436
rect 10540 17434 10564 17436
rect 10620 17434 10644 17436
rect 10700 17434 10706 17436
rect 10460 17382 10462 17434
rect 10642 17382 10644 17434
rect 10398 17380 10404 17382
rect 10460 17380 10484 17382
rect 10540 17380 10564 17382
rect 10620 17380 10644 17382
rect 10700 17380 10706 17382
rect 10398 17371 10706 17380
rect 9680 16788 9732 16794
rect 9680 16730 9732 16736
rect 9588 16584 9640 16590
rect 9588 16526 9640 16532
rect 9496 15904 9548 15910
rect 9496 15846 9548 15852
rect 9404 15632 9456 15638
rect 9404 15574 9456 15580
rect 9600 14074 9628 16526
rect 9692 15706 9720 16730
rect 9956 16720 10008 16726
rect 9956 16662 10008 16668
rect 9968 16590 9996 16662
rect 9956 16584 10008 16590
rect 9956 16526 10008 16532
rect 10784 16584 10836 16590
rect 10784 16526 10836 16532
rect 10398 16348 10706 16357
rect 10398 16346 10404 16348
rect 10460 16346 10484 16348
rect 10540 16346 10564 16348
rect 10620 16346 10644 16348
rect 10700 16346 10706 16348
rect 10460 16294 10462 16346
rect 10642 16294 10644 16346
rect 10398 16292 10404 16294
rect 10460 16292 10484 16294
rect 10540 16292 10564 16294
rect 10620 16292 10644 16294
rect 10700 16292 10706 16294
rect 10398 16283 10706 16292
rect 10796 16250 10824 16526
rect 10980 16522 11008 17546
rect 12084 16658 12112 21898
rect 12360 21894 12388 25214
rect 12728 24614 12756 25298
rect 12716 24608 12768 24614
rect 12716 24550 12768 24556
rect 12164 21888 12216 21894
rect 12164 21830 12216 21836
rect 12348 21888 12400 21894
rect 12348 21830 12400 21836
rect 11704 16652 11756 16658
rect 11704 16594 11756 16600
rect 12072 16652 12124 16658
rect 12072 16594 12124 16600
rect 10968 16516 11020 16522
rect 10968 16458 11020 16464
rect 11336 16448 11388 16454
rect 11336 16390 11388 16396
rect 10784 16244 10836 16250
rect 10784 16186 10836 16192
rect 11060 16176 11112 16182
rect 11060 16118 11112 16124
rect 10140 16040 10192 16046
rect 10140 15982 10192 15988
rect 10324 16040 10376 16046
rect 10324 15982 10376 15988
rect 9680 15700 9732 15706
rect 9680 15642 9732 15648
rect 9680 15360 9732 15366
rect 9680 15302 9732 15308
rect 9692 14414 9720 15302
rect 10152 14958 10180 15982
rect 10140 14952 10192 14958
rect 10140 14894 10192 14900
rect 9680 14408 9732 14414
rect 9680 14350 9732 14356
rect 9588 14068 9640 14074
rect 9588 14010 9640 14016
rect 9312 13320 9364 13326
rect 9312 13262 9364 13268
rect 9324 12986 9352 13262
rect 9312 12980 9364 12986
rect 9312 12922 9364 12928
rect 9600 12238 9628 14010
rect 10152 12434 10180 14894
rect 10336 14482 10364 15982
rect 11072 15434 11100 16118
rect 11348 15978 11376 16390
rect 11716 16250 11744 16594
rect 11704 16244 11756 16250
rect 11704 16186 11756 16192
rect 11704 16040 11756 16046
rect 11704 15982 11756 15988
rect 11336 15972 11388 15978
rect 11336 15914 11388 15920
rect 11716 15638 11744 15982
rect 11704 15632 11756 15638
rect 11704 15574 11756 15580
rect 11060 15428 11112 15434
rect 11060 15370 11112 15376
rect 10398 15260 10706 15269
rect 10398 15258 10404 15260
rect 10460 15258 10484 15260
rect 10540 15258 10564 15260
rect 10620 15258 10644 15260
rect 10700 15258 10706 15260
rect 10460 15206 10462 15258
rect 10642 15206 10644 15258
rect 10398 15204 10404 15206
rect 10460 15204 10484 15206
rect 10540 15204 10564 15206
rect 10620 15204 10644 15206
rect 10700 15204 10706 15206
rect 10398 15195 10706 15204
rect 11072 15026 11100 15370
rect 11060 15020 11112 15026
rect 11060 14962 11112 14968
rect 10324 14476 10376 14482
rect 10324 14418 10376 14424
rect 10398 14172 10706 14181
rect 10398 14170 10404 14172
rect 10460 14170 10484 14172
rect 10540 14170 10564 14172
rect 10620 14170 10644 14172
rect 10700 14170 10706 14172
rect 10460 14118 10462 14170
rect 10642 14118 10644 14170
rect 10398 14116 10404 14118
rect 10460 14116 10484 14118
rect 10540 14116 10564 14118
rect 10620 14116 10644 14118
rect 10700 14116 10706 14118
rect 10398 14107 10706 14116
rect 10398 13084 10706 13093
rect 10398 13082 10404 13084
rect 10460 13082 10484 13084
rect 10540 13082 10564 13084
rect 10620 13082 10644 13084
rect 10700 13082 10706 13084
rect 10460 13030 10462 13082
rect 10642 13030 10644 13082
rect 10398 13028 10404 13030
rect 10460 13028 10484 13030
rect 10540 13028 10564 13030
rect 10620 13028 10644 13030
rect 10700 13028 10706 13030
rect 10398 13019 10706 13028
rect 9968 12406 10180 12434
rect 9588 12232 9640 12238
rect 9588 12174 9640 12180
rect 9220 12096 9272 12102
rect 9220 12038 9272 12044
rect 9128 11892 9180 11898
rect 9128 11834 9180 11840
rect 9232 11762 9260 12038
rect 9220 11756 9272 11762
rect 9220 11698 9272 11704
rect 9968 11558 9996 12406
rect 10398 11996 10706 12005
rect 10398 11994 10404 11996
rect 10460 11994 10484 11996
rect 10540 11994 10564 11996
rect 10620 11994 10644 11996
rect 10700 11994 10706 11996
rect 10460 11942 10462 11994
rect 10642 11942 10644 11994
rect 10398 11940 10404 11942
rect 10460 11940 10484 11942
rect 10540 11940 10564 11942
rect 10620 11940 10644 11942
rect 10700 11940 10706 11942
rect 10398 11931 10706 11940
rect 10048 11824 10100 11830
rect 10048 11766 10100 11772
rect 9956 11552 10008 11558
rect 9956 11494 10008 11500
rect 10060 11354 10088 11766
rect 11796 11756 11848 11762
rect 11796 11698 11848 11704
rect 10140 11688 10192 11694
rect 10140 11630 10192 11636
rect 10048 11348 10100 11354
rect 10048 11290 10100 11296
rect 10152 11150 10180 11630
rect 10140 11144 10192 11150
rect 10140 11086 10192 11092
rect 10152 8498 10180 11086
rect 10398 10908 10706 10917
rect 10398 10906 10404 10908
rect 10460 10906 10484 10908
rect 10540 10906 10564 10908
rect 10620 10906 10644 10908
rect 10700 10906 10706 10908
rect 10460 10854 10462 10906
rect 10642 10854 10644 10906
rect 10398 10852 10404 10854
rect 10460 10852 10484 10854
rect 10540 10852 10564 10854
rect 10620 10852 10644 10854
rect 10700 10852 10706 10854
rect 10398 10843 10706 10852
rect 10398 9820 10706 9829
rect 10398 9818 10404 9820
rect 10460 9818 10484 9820
rect 10540 9818 10564 9820
rect 10620 9818 10644 9820
rect 10700 9818 10706 9820
rect 10460 9766 10462 9818
rect 10642 9766 10644 9818
rect 10398 9764 10404 9766
rect 10460 9764 10484 9766
rect 10540 9764 10564 9766
rect 10620 9764 10644 9766
rect 10700 9764 10706 9766
rect 10398 9755 10706 9764
rect 10398 8732 10706 8741
rect 10398 8730 10404 8732
rect 10460 8730 10484 8732
rect 10540 8730 10564 8732
rect 10620 8730 10644 8732
rect 10700 8730 10706 8732
rect 10460 8678 10462 8730
rect 10642 8678 10644 8730
rect 10398 8676 10404 8678
rect 10460 8676 10484 8678
rect 10540 8676 10564 8678
rect 10620 8676 10644 8678
rect 10700 8676 10706 8678
rect 10398 8667 10706 8676
rect 10140 8492 10192 8498
rect 10140 8434 10192 8440
rect 9036 7948 9088 7954
rect 9036 7890 9088 7896
rect 9496 7812 9548 7818
rect 9496 7754 9548 7760
rect 9956 7812 10008 7818
rect 9956 7754 10008 7760
rect 9508 4010 9536 7754
rect 9968 7546 9996 7754
rect 9956 7540 10008 7546
rect 9956 7482 10008 7488
rect 10152 7410 10180 8434
rect 11808 7954 11836 11698
rect 11796 7948 11848 7954
rect 11796 7890 11848 7896
rect 10398 7644 10706 7653
rect 10398 7642 10404 7644
rect 10460 7642 10484 7644
rect 10540 7642 10564 7644
rect 10620 7642 10644 7644
rect 10700 7642 10706 7644
rect 10460 7590 10462 7642
rect 10642 7590 10644 7642
rect 10398 7588 10404 7590
rect 10460 7588 10484 7590
rect 10540 7588 10564 7590
rect 10620 7588 10644 7590
rect 10700 7588 10706 7590
rect 10398 7579 10706 7588
rect 11808 7546 11836 7890
rect 12072 7812 12124 7818
rect 12072 7754 12124 7760
rect 11796 7540 11848 7546
rect 11796 7482 11848 7488
rect 10140 7404 10192 7410
rect 10140 7346 10192 7352
rect 10398 6556 10706 6565
rect 10398 6554 10404 6556
rect 10460 6554 10484 6556
rect 10540 6554 10564 6556
rect 10620 6554 10644 6556
rect 10700 6554 10706 6556
rect 10460 6502 10462 6554
rect 10642 6502 10644 6554
rect 10398 6500 10404 6502
rect 10460 6500 10484 6502
rect 10540 6500 10564 6502
rect 10620 6500 10644 6502
rect 10700 6500 10706 6502
rect 10398 6491 10706 6500
rect 10398 5468 10706 5477
rect 10398 5466 10404 5468
rect 10460 5466 10484 5468
rect 10540 5466 10564 5468
rect 10620 5466 10644 5468
rect 10700 5466 10706 5468
rect 10460 5414 10462 5466
rect 10642 5414 10644 5466
rect 10398 5412 10404 5414
rect 10460 5412 10484 5414
rect 10540 5412 10564 5414
rect 10620 5412 10644 5414
rect 10700 5412 10706 5414
rect 10398 5403 10706 5412
rect 10398 4380 10706 4389
rect 10398 4378 10404 4380
rect 10460 4378 10484 4380
rect 10540 4378 10564 4380
rect 10620 4378 10644 4380
rect 10700 4378 10706 4380
rect 10460 4326 10462 4378
rect 10642 4326 10644 4378
rect 10398 4324 10404 4326
rect 10460 4324 10484 4326
rect 10540 4324 10564 4326
rect 10620 4324 10644 4326
rect 10700 4324 10706 4326
rect 10398 4315 10706 4324
rect 11980 4140 12032 4146
rect 11980 4082 12032 4088
rect 10508 4072 10560 4078
rect 10508 4014 10560 4020
rect 9496 4004 9548 4010
rect 9496 3946 9548 3952
rect 10520 3602 10548 4014
rect 10784 3936 10836 3942
rect 10784 3878 10836 3884
rect 10508 3596 10560 3602
rect 10508 3538 10560 3544
rect 10796 3534 10824 3878
rect 11992 3670 12020 4082
rect 12084 3738 12112 7754
rect 12176 7342 12204 21830
rect 12256 18624 12308 18630
rect 12256 18566 12308 18572
rect 12268 15978 12296 18566
rect 12912 18426 12940 32166
rect 13176 31272 13228 31278
rect 13176 31214 13228 31220
rect 13188 30802 13216 31214
rect 13176 30796 13228 30802
rect 13176 30738 13228 30744
rect 13820 30184 13872 30190
rect 13820 30126 13872 30132
rect 12992 29164 13044 29170
rect 12992 29106 13044 29112
rect 13004 28762 13032 29106
rect 13832 29102 13860 30126
rect 13820 29096 13872 29102
rect 13820 29038 13872 29044
rect 13452 28960 13504 28966
rect 13452 28902 13504 28908
rect 12992 28756 13044 28762
rect 12992 28698 13044 28704
rect 13464 28626 13492 28902
rect 13832 28626 13860 29038
rect 13452 28620 13504 28626
rect 13452 28562 13504 28568
rect 13820 28620 13872 28626
rect 13820 28562 13872 28568
rect 13464 27878 13492 28562
rect 13452 27872 13504 27878
rect 13452 27814 13504 27820
rect 13268 24948 13320 24954
rect 13268 24890 13320 24896
rect 13280 23730 13308 24890
rect 13268 23724 13320 23730
rect 13268 23666 13320 23672
rect 12992 22432 13044 22438
rect 12992 22374 13044 22380
rect 13004 22030 13032 22374
rect 12992 22024 13044 22030
rect 12992 21966 13044 21972
rect 12900 18420 12952 18426
rect 12900 18362 12952 18368
rect 12912 18222 12940 18362
rect 12900 18216 12952 18222
rect 12900 18158 12952 18164
rect 13268 18216 13320 18222
rect 13268 18158 13320 18164
rect 12348 16448 12400 16454
rect 12348 16390 12400 16396
rect 12360 16114 12388 16390
rect 12348 16108 12400 16114
rect 12348 16050 12400 16056
rect 12256 15972 12308 15978
rect 12256 15914 12308 15920
rect 12268 15502 12296 15914
rect 12256 15496 12308 15502
rect 12256 15438 12308 15444
rect 13280 12646 13308 18158
rect 13464 17338 13492 27814
rect 13544 24608 13596 24614
rect 13544 24550 13596 24556
rect 13556 23798 13584 24550
rect 13544 23792 13596 23798
rect 13544 23734 13596 23740
rect 13556 22506 13584 23734
rect 13832 22574 13860 28562
rect 14108 28558 14136 33458
rect 15122 33212 15430 33221
rect 15122 33210 15128 33212
rect 15184 33210 15208 33212
rect 15264 33210 15288 33212
rect 15344 33210 15368 33212
rect 15424 33210 15430 33212
rect 15184 33158 15186 33210
rect 15366 33158 15368 33210
rect 15122 33156 15128 33158
rect 15184 33156 15208 33158
rect 15264 33156 15288 33158
rect 15344 33156 15368 33158
rect 15424 33156 15430 33158
rect 15122 33147 15430 33156
rect 24570 33212 24878 33221
rect 24570 33210 24576 33212
rect 24632 33210 24656 33212
rect 24712 33210 24736 33212
rect 24792 33210 24816 33212
rect 24872 33210 24878 33212
rect 24632 33158 24634 33210
rect 24814 33158 24816 33210
rect 24570 33156 24576 33158
rect 24632 33156 24656 33158
rect 24712 33156 24736 33158
rect 24792 33156 24816 33158
rect 24872 33156 24878 33158
rect 24570 33147 24878 33156
rect 34018 33212 34326 33221
rect 34018 33210 34024 33212
rect 34080 33210 34104 33212
rect 34160 33210 34184 33212
rect 34240 33210 34264 33212
rect 34320 33210 34326 33212
rect 34080 33158 34082 33210
rect 34262 33158 34264 33210
rect 34018 33156 34024 33158
rect 34080 33156 34104 33158
rect 34160 33156 34184 33158
rect 34240 33156 34264 33158
rect 34320 33156 34326 33158
rect 34018 33147 34326 33156
rect 19846 32668 20154 32677
rect 19846 32666 19852 32668
rect 19908 32666 19932 32668
rect 19988 32666 20012 32668
rect 20068 32666 20092 32668
rect 20148 32666 20154 32668
rect 19908 32614 19910 32666
rect 20090 32614 20092 32666
rect 19846 32612 19852 32614
rect 19908 32612 19932 32614
rect 19988 32612 20012 32614
rect 20068 32612 20092 32614
rect 20148 32612 20154 32614
rect 19846 32603 20154 32612
rect 29294 32668 29602 32677
rect 29294 32666 29300 32668
rect 29356 32666 29380 32668
rect 29436 32666 29460 32668
rect 29516 32666 29540 32668
rect 29596 32666 29602 32668
rect 29356 32614 29358 32666
rect 29538 32614 29540 32666
rect 29294 32612 29300 32614
rect 29356 32612 29380 32614
rect 29436 32612 29460 32614
rect 29516 32612 29540 32614
rect 29596 32612 29602 32614
rect 29294 32603 29602 32612
rect 17224 32496 17276 32502
rect 17224 32438 17276 32444
rect 16396 32428 16448 32434
rect 16396 32370 16448 32376
rect 15122 32124 15430 32133
rect 15122 32122 15128 32124
rect 15184 32122 15208 32124
rect 15264 32122 15288 32124
rect 15344 32122 15368 32124
rect 15424 32122 15430 32124
rect 15184 32070 15186 32122
rect 15366 32070 15368 32122
rect 15122 32068 15128 32070
rect 15184 32068 15208 32070
rect 15264 32068 15288 32070
rect 15344 32068 15368 32070
rect 15424 32068 15430 32070
rect 15122 32059 15430 32068
rect 16408 31958 16436 32370
rect 16396 31952 16448 31958
rect 16396 31894 16448 31900
rect 17236 31822 17264 32438
rect 18328 32224 18380 32230
rect 18328 32166 18380 32172
rect 22376 32224 22428 32230
rect 22376 32166 22428 32172
rect 18340 31958 18368 32166
rect 18788 32020 18840 32026
rect 18788 31962 18840 31968
rect 18328 31952 18380 31958
rect 18328 31894 18380 31900
rect 16212 31816 16264 31822
rect 16212 31758 16264 31764
rect 17224 31816 17276 31822
rect 17224 31758 17276 31764
rect 17592 31816 17644 31822
rect 17592 31758 17644 31764
rect 16224 31482 16252 31758
rect 16212 31476 16264 31482
rect 16212 31418 16264 31424
rect 15844 31340 15896 31346
rect 15844 31282 15896 31288
rect 15660 31272 15712 31278
rect 15660 31214 15712 31220
rect 15122 31036 15430 31045
rect 15122 31034 15128 31036
rect 15184 31034 15208 31036
rect 15264 31034 15288 31036
rect 15344 31034 15368 31036
rect 15424 31034 15430 31036
rect 15184 30982 15186 31034
rect 15366 30982 15368 31034
rect 15122 30980 15128 30982
rect 15184 30980 15208 30982
rect 15264 30980 15288 30982
rect 15344 30980 15368 30982
rect 15424 30980 15430 30982
rect 15122 30971 15430 30980
rect 15672 30938 15700 31214
rect 15660 30932 15712 30938
rect 15660 30874 15712 30880
rect 15122 29948 15430 29957
rect 15122 29946 15128 29948
rect 15184 29946 15208 29948
rect 15264 29946 15288 29948
rect 15344 29946 15368 29948
rect 15424 29946 15430 29948
rect 15184 29894 15186 29946
rect 15366 29894 15368 29946
rect 15122 29892 15128 29894
rect 15184 29892 15208 29894
rect 15264 29892 15288 29894
rect 15344 29892 15368 29894
rect 15424 29892 15430 29894
rect 15122 29883 15430 29892
rect 15122 28860 15430 28869
rect 15122 28858 15128 28860
rect 15184 28858 15208 28860
rect 15264 28858 15288 28860
rect 15344 28858 15368 28860
rect 15424 28858 15430 28860
rect 15184 28806 15186 28858
rect 15366 28806 15368 28858
rect 15122 28804 15128 28806
rect 15184 28804 15208 28806
rect 15264 28804 15288 28806
rect 15344 28804 15368 28806
rect 15424 28804 15430 28806
rect 15122 28795 15430 28804
rect 14004 28552 14056 28558
rect 14004 28494 14056 28500
rect 14096 28552 14148 28558
rect 14096 28494 14148 28500
rect 14016 26586 14044 28494
rect 15122 27772 15430 27781
rect 15122 27770 15128 27772
rect 15184 27770 15208 27772
rect 15264 27770 15288 27772
rect 15344 27770 15368 27772
rect 15424 27770 15430 27772
rect 15184 27718 15186 27770
rect 15366 27718 15368 27770
rect 15122 27716 15128 27718
rect 15184 27716 15208 27718
rect 15264 27716 15288 27718
rect 15344 27716 15368 27718
rect 15424 27716 15430 27718
rect 15122 27707 15430 27716
rect 14924 26784 14976 26790
rect 14924 26726 14976 26732
rect 14004 26580 14056 26586
rect 14004 26522 14056 26528
rect 14936 26450 14964 26726
rect 15122 26684 15430 26693
rect 15122 26682 15128 26684
rect 15184 26682 15208 26684
rect 15264 26682 15288 26684
rect 15344 26682 15368 26684
rect 15424 26682 15430 26684
rect 15184 26630 15186 26682
rect 15366 26630 15368 26682
rect 15122 26628 15128 26630
rect 15184 26628 15208 26630
rect 15264 26628 15288 26630
rect 15344 26628 15368 26630
rect 15424 26628 15430 26630
rect 15122 26619 15430 26628
rect 14924 26444 14976 26450
rect 14924 26386 14976 26392
rect 15016 26376 15068 26382
rect 15016 26318 15068 26324
rect 15568 26376 15620 26382
rect 15568 26318 15620 26324
rect 15028 25294 15056 26318
rect 15122 25596 15430 25605
rect 15122 25594 15128 25596
rect 15184 25594 15208 25596
rect 15264 25594 15288 25596
rect 15344 25594 15368 25596
rect 15424 25594 15430 25596
rect 15184 25542 15186 25594
rect 15366 25542 15368 25594
rect 15122 25540 15128 25542
rect 15184 25540 15208 25542
rect 15264 25540 15288 25542
rect 15344 25540 15368 25542
rect 15424 25540 15430 25542
rect 15122 25531 15430 25540
rect 15580 25362 15608 26318
rect 15568 25356 15620 25362
rect 15568 25298 15620 25304
rect 15016 25288 15068 25294
rect 15016 25230 15068 25236
rect 15028 24818 15056 25230
rect 15016 24812 15068 24818
rect 15016 24754 15068 24760
rect 13912 23724 13964 23730
rect 13912 23666 13964 23672
rect 13924 23526 13952 23666
rect 13912 23520 13964 23526
rect 13912 23462 13964 23468
rect 13820 22568 13872 22574
rect 13820 22510 13872 22516
rect 13544 22500 13596 22506
rect 13544 22442 13596 22448
rect 13452 17332 13504 17338
rect 13452 17274 13504 17280
rect 13820 15088 13872 15094
rect 13820 15030 13872 15036
rect 13832 13462 13860 15030
rect 13820 13456 13872 13462
rect 13820 13398 13872 13404
rect 13832 12730 13860 13398
rect 13740 12702 13860 12730
rect 13268 12640 13320 12646
rect 13268 12582 13320 12588
rect 13636 12640 13688 12646
rect 13636 12582 13688 12588
rect 12716 12300 12768 12306
rect 12716 12242 12768 12248
rect 12728 11898 12756 12242
rect 13648 12238 13676 12582
rect 13740 12306 13768 12702
rect 13820 12640 13872 12646
rect 13820 12582 13872 12588
rect 13728 12300 13780 12306
rect 13728 12242 13780 12248
rect 13268 12232 13320 12238
rect 13268 12174 13320 12180
rect 13636 12232 13688 12238
rect 13636 12174 13688 12180
rect 13176 12096 13228 12102
rect 13176 12038 13228 12044
rect 12716 11892 12768 11898
rect 12716 11834 12768 11840
rect 13188 11830 13216 12038
rect 13176 11824 13228 11830
rect 13176 11766 13228 11772
rect 13280 11150 13308 12174
rect 13648 11762 13676 12174
rect 13636 11756 13688 11762
rect 13636 11698 13688 11704
rect 13648 11354 13676 11698
rect 13832 11626 13860 12582
rect 13820 11620 13872 11626
rect 13820 11562 13872 11568
rect 13924 11370 13952 23462
rect 15028 22642 15056 24754
rect 15122 24508 15430 24517
rect 15122 24506 15128 24508
rect 15184 24506 15208 24508
rect 15264 24506 15288 24508
rect 15344 24506 15368 24508
rect 15424 24506 15430 24508
rect 15184 24454 15186 24506
rect 15366 24454 15368 24506
rect 15122 24452 15128 24454
rect 15184 24452 15208 24454
rect 15264 24452 15288 24454
rect 15344 24452 15368 24454
rect 15424 24452 15430 24454
rect 15122 24443 15430 24452
rect 15122 23420 15430 23429
rect 15122 23418 15128 23420
rect 15184 23418 15208 23420
rect 15264 23418 15288 23420
rect 15344 23418 15368 23420
rect 15424 23418 15430 23420
rect 15184 23366 15186 23418
rect 15366 23366 15368 23418
rect 15122 23364 15128 23366
rect 15184 23364 15208 23366
rect 15264 23364 15288 23366
rect 15344 23364 15368 23366
rect 15424 23364 15430 23366
rect 15122 23355 15430 23364
rect 15580 23322 15608 25298
rect 15672 24614 15700 30874
rect 15856 29170 15884 31282
rect 15844 29164 15896 29170
rect 15844 29106 15896 29112
rect 17236 29102 17264 31758
rect 17604 31482 17632 31758
rect 17592 31476 17644 31482
rect 17592 31418 17644 31424
rect 17500 29164 17552 29170
rect 17500 29106 17552 29112
rect 17224 29096 17276 29102
rect 17224 29038 17276 29044
rect 16672 29028 16724 29034
rect 16672 28970 16724 28976
rect 16684 28558 16712 28970
rect 17236 28694 17264 29038
rect 17512 28762 17540 29106
rect 18340 29034 18368 31894
rect 18328 29028 18380 29034
rect 18328 28970 18380 28976
rect 17500 28756 17552 28762
rect 17500 28698 17552 28704
rect 17224 28688 17276 28694
rect 17224 28630 17276 28636
rect 16672 28552 16724 28558
rect 16672 28494 16724 28500
rect 16028 26376 16080 26382
rect 16028 26318 16080 26324
rect 15752 26240 15804 26246
rect 15752 26182 15804 26188
rect 15764 25906 15792 26182
rect 16040 26042 16068 26318
rect 17040 26240 17092 26246
rect 17040 26182 17092 26188
rect 16028 26036 16080 26042
rect 16028 25978 16080 25984
rect 15752 25900 15804 25906
rect 15752 25842 15804 25848
rect 17052 25702 17080 26182
rect 17040 25696 17092 25702
rect 17040 25638 17092 25644
rect 15844 25288 15896 25294
rect 15844 25230 15896 25236
rect 15856 24954 15884 25230
rect 17052 25158 17080 25638
rect 17040 25152 17092 25158
rect 17040 25094 17092 25100
rect 15844 24948 15896 24954
rect 15844 24890 15896 24896
rect 15660 24608 15712 24614
rect 15660 24550 15712 24556
rect 16856 23724 16908 23730
rect 16856 23666 16908 23672
rect 16672 23520 16724 23526
rect 16672 23462 16724 23468
rect 15568 23316 15620 23322
rect 15568 23258 15620 23264
rect 14740 22636 14792 22642
rect 14740 22578 14792 22584
rect 15016 22636 15068 22642
rect 15016 22578 15068 22584
rect 14752 22098 14780 22578
rect 15122 22332 15430 22341
rect 15122 22330 15128 22332
rect 15184 22330 15208 22332
rect 15264 22330 15288 22332
rect 15344 22330 15368 22332
rect 15424 22330 15430 22332
rect 15184 22278 15186 22330
rect 15366 22278 15368 22330
rect 15122 22276 15128 22278
rect 15184 22276 15208 22278
rect 15264 22276 15288 22278
rect 15344 22276 15368 22278
rect 15424 22276 15430 22278
rect 15122 22267 15430 22276
rect 14740 22092 14792 22098
rect 14740 22034 14792 22040
rect 14832 21956 14884 21962
rect 14832 21898 14884 21904
rect 14844 20058 14872 21898
rect 15122 21244 15430 21253
rect 15122 21242 15128 21244
rect 15184 21242 15208 21244
rect 15264 21242 15288 21244
rect 15344 21242 15368 21244
rect 15424 21242 15430 21244
rect 15184 21190 15186 21242
rect 15366 21190 15368 21242
rect 15122 21188 15128 21190
rect 15184 21188 15208 21190
rect 15264 21188 15288 21190
rect 15344 21188 15368 21190
rect 15424 21188 15430 21190
rect 15122 21179 15430 21188
rect 15122 20156 15430 20165
rect 15122 20154 15128 20156
rect 15184 20154 15208 20156
rect 15264 20154 15288 20156
rect 15344 20154 15368 20156
rect 15424 20154 15430 20156
rect 15184 20102 15186 20154
rect 15366 20102 15368 20154
rect 15122 20100 15128 20102
rect 15184 20100 15208 20102
rect 15264 20100 15288 20102
rect 15344 20100 15368 20102
rect 15424 20100 15430 20102
rect 15122 20091 15430 20100
rect 14832 20052 14884 20058
rect 14832 19994 14884 20000
rect 14556 19780 14608 19786
rect 14556 19722 14608 19728
rect 14568 18290 14596 19722
rect 14844 19378 14872 19994
rect 15580 19922 15608 23258
rect 16684 23118 16712 23462
rect 16672 23112 16724 23118
rect 16672 23054 16724 23060
rect 16868 22778 16896 23666
rect 17052 22982 17080 25094
rect 17040 22976 17092 22982
rect 17040 22918 17092 22924
rect 16856 22772 16908 22778
rect 16856 22714 16908 22720
rect 17052 20058 17080 22918
rect 18800 21554 18828 31962
rect 22388 31958 22416 32166
rect 24570 32124 24878 32133
rect 24570 32122 24576 32124
rect 24632 32122 24656 32124
rect 24712 32122 24736 32124
rect 24792 32122 24816 32124
rect 24872 32122 24878 32124
rect 24632 32070 24634 32122
rect 24814 32070 24816 32122
rect 24570 32068 24576 32070
rect 24632 32068 24656 32070
rect 24712 32068 24736 32070
rect 24792 32068 24816 32070
rect 24872 32068 24878 32070
rect 24570 32059 24878 32068
rect 34018 32124 34326 32133
rect 34018 32122 34024 32124
rect 34080 32122 34104 32124
rect 34160 32122 34184 32124
rect 34240 32122 34264 32124
rect 34320 32122 34326 32124
rect 34080 32070 34082 32122
rect 34262 32070 34264 32122
rect 34018 32068 34024 32070
rect 34080 32068 34104 32070
rect 34160 32068 34184 32070
rect 34240 32068 34264 32070
rect 34320 32068 34326 32070
rect 34018 32059 34326 32068
rect 23480 32020 23532 32026
rect 23480 31962 23532 31968
rect 25412 32020 25464 32026
rect 25412 31962 25464 31968
rect 29000 32020 29052 32026
rect 29000 31962 29052 31968
rect 22376 31952 22428 31958
rect 22376 31894 22428 31900
rect 20720 31816 20772 31822
rect 20720 31758 20772 31764
rect 22100 31816 22152 31822
rect 22100 31758 22152 31764
rect 19846 31580 20154 31589
rect 19846 31578 19852 31580
rect 19908 31578 19932 31580
rect 19988 31578 20012 31580
rect 20068 31578 20092 31580
rect 20148 31578 20154 31580
rect 19908 31526 19910 31578
rect 20090 31526 20092 31578
rect 19846 31524 19852 31526
rect 19908 31524 19932 31526
rect 19988 31524 20012 31526
rect 20068 31524 20092 31526
rect 20148 31524 20154 31526
rect 19846 31515 20154 31524
rect 20732 31482 20760 31758
rect 22112 31482 22140 31758
rect 20720 31476 20772 31482
rect 20720 31418 20772 31424
rect 22100 31476 22152 31482
rect 22100 31418 22152 31424
rect 21180 31340 21232 31346
rect 21180 31282 21232 31288
rect 21364 31340 21416 31346
rect 21364 31282 21416 31288
rect 19524 31272 19576 31278
rect 19524 31214 19576 31220
rect 19432 29028 19484 29034
rect 19432 28970 19484 28976
rect 19444 27946 19472 28970
rect 19340 27940 19392 27946
rect 19340 27882 19392 27888
rect 19432 27940 19484 27946
rect 19432 27882 19484 27888
rect 19352 27334 19380 27882
rect 19340 27328 19392 27334
rect 19340 27270 19392 27276
rect 19352 21690 19380 27270
rect 19340 21684 19392 21690
rect 19340 21626 19392 21632
rect 18788 21548 18840 21554
rect 18788 21490 18840 21496
rect 19248 21548 19300 21554
rect 19248 21490 19300 21496
rect 19260 20806 19288 21490
rect 19248 20800 19300 20806
rect 19248 20742 19300 20748
rect 19260 20534 19288 20742
rect 19248 20528 19300 20534
rect 19248 20470 19300 20476
rect 17224 20392 17276 20398
rect 17224 20334 17276 20340
rect 17040 20052 17092 20058
rect 17040 19994 17092 20000
rect 15568 19916 15620 19922
rect 15568 19858 15620 19864
rect 17040 19848 17092 19854
rect 17040 19790 17092 19796
rect 17052 19514 17080 19790
rect 17040 19508 17092 19514
rect 17040 19450 17092 19456
rect 14832 19372 14884 19378
rect 14832 19314 14884 19320
rect 17236 19310 17264 20334
rect 17224 19304 17276 19310
rect 17224 19246 17276 19252
rect 15122 19068 15430 19077
rect 15122 19066 15128 19068
rect 15184 19066 15208 19068
rect 15264 19066 15288 19068
rect 15344 19066 15368 19068
rect 15424 19066 15430 19068
rect 15184 19014 15186 19066
rect 15366 19014 15368 19066
rect 15122 19012 15128 19014
rect 15184 19012 15208 19014
rect 15264 19012 15288 19014
rect 15344 19012 15368 19014
rect 15424 19012 15430 19014
rect 15122 19003 15430 19012
rect 14372 18284 14424 18290
rect 14372 18226 14424 18232
rect 14556 18284 14608 18290
rect 14556 18226 14608 18232
rect 14280 18080 14332 18086
rect 14280 18022 14332 18028
rect 14292 17882 14320 18022
rect 14280 17876 14332 17882
rect 14280 17818 14332 17824
rect 14384 17678 14412 18226
rect 14372 17672 14424 17678
rect 14372 17614 14424 17620
rect 14568 16590 14596 18226
rect 15122 17980 15430 17989
rect 15122 17978 15128 17980
rect 15184 17978 15208 17980
rect 15264 17978 15288 17980
rect 15344 17978 15368 17980
rect 15424 17978 15430 17980
rect 15184 17926 15186 17978
rect 15366 17926 15368 17978
rect 15122 17924 15128 17926
rect 15184 17924 15208 17926
rect 15264 17924 15288 17926
rect 15344 17924 15368 17926
rect 15424 17924 15430 17926
rect 15122 17915 15430 17924
rect 14740 17672 14792 17678
rect 14740 17614 14792 17620
rect 15476 17672 15528 17678
rect 15476 17614 15528 17620
rect 14556 16584 14608 16590
rect 14556 16526 14608 16532
rect 14372 16516 14424 16522
rect 14372 16458 14424 16464
rect 14384 15502 14412 16458
rect 14372 15496 14424 15502
rect 14372 15438 14424 15444
rect 14556 15496 14608 15502
rect 14556 15438 14608 15444
rect 14568 15094 14596 15438
rect 14556 15088 14608 15094
rect 14556 15030 14608 15036
rect 14556 13320 14608 13326
rect 14556 13262 14608 13268
rect 14464 12844 14516 12850
rect 14464 12786 14516 12792
rect 14004 12776 14056 12782
rect 14004 12718 14056 12724
rect 14372 12776 14424 12782
rect 14372 12718 14424 12724
rect 14016 12374 14044 12718
rect 14004 12368 14056 12374
rect 14004 12310 14056 12316
rect 14384 12306 14412 12718
rect 14372 12300 14424 12306
rect 14372 12242 14424 12248
rect 14372 12164 14424 12170
rect 14372 12106 14424 12112
rect 14384 11762 14412 12106
rect 14476 12102 14504 12786
rect 14464 12096 14516 12102
rect 14464 12038 14516 12044
rect 14476 11898 14504 12038
rect 14568 11898 14596 13262
rect 14648 12708 14700 12714
rect 14648 12650 14700 12656
rect 14660 12102 14688 12650
rect 14648 12096 14700 12102
rect 14648 12038 14700 12044
rect 14464 11892 14516 11898
rect 14464 11834 14516 11840
rect 14556 11892 14608 11898
rect 14556 11834 14608 11840
rect 14372 11756 14424 11762
rect 14372 11698 14424 11704
rect 14280 11552 14332 11558
rect 14280 11494 14332 11500
rect 13636 11348 13688 11354
rect 13636 11290 13688 11296
rect 13832 11342 13952 11370
rect 14292 11354 14320 11494
rect 14280 11348 14332 11354
rect 13268 11144 13320 11150
rect 13268 11086 13320 11092
rect 13280 9654 13308 11086
rect 13268 9648 13320 9654
rect 13268 9590 13320 9596
rect 13832 8906 13860 11342
rect 14280 11290 14332 11296
rect 14568 11286 14596 11834
rect 14556 11280 14608 11286
rect 14556 11222 14608 11228
rect 14568 10742 14596 11222
rect 14660 11150 14688 12038
rect 14752 11762 14780 17614
rect 15122 16892 15430 16901
rect 15122 16890 15128 16892
rect 15184 16890 15208 16892
rect 15264 16890 15288 16892
rect 15344 16890 15368 16892
rect 15424 16890 15430 16892
rect 15184 16838 15186 16890
rect 15366 16838 15368 16890
rect 15122 16836 15128 16838
rect 15184 16836 15208 16838
rect 15264 16836 15288 16838
rect 15344 16836 15368 16838
rect 15424 16836 15430 16838
rect 15122 16827 15430 16836
rect 14832 16176 14884 16182
rect 14832 16118 14884 16124
rect 14844 15502 14872 16118
rect 15122 15804 15430 15813
rect 15122 15802 15128 15804
rect 15184 15802 15208 15804
rect 15264 15802 15288 15804
rect 15344 15802 15368 15804
rect 15424 15802 15430 15804
rect 15184 15750 15186 15802
rect 15366 15750 15368 15802
rect 15122 15748 15128 15750
rect 15184 15748 15208 15750
rect 15264 15748 15288 15750
rect 15344 15748 15368 15750
rect 15424 15748 15430 15750
rect 15122 15739 15430 15748
rect 14832 15496 14884 15502
rect 14832 15438 14884 15444
rect 14844 15026 14872 15438
rect 14832 15020 14884 15026
rect 14832 14962 14884 14968
rect 15122 14716 15430 14725
rect 15122 14714 15128 14716
rect 15184 14714 15208 14716
rect 15264 14714 15288 14716
rect 15344 14714 15368 14716
rect 15424 14714 15430 14716
rect 15184 14662 15186 14714
rect 15366 14662 15368 14714
rect 15122 14660 15128 14662
rect 15184 14660 15208 14662
rect 15264 14660 15288 14662
rect 15344 14660 15368 14662
rect 15424 14660 15430 14662
rect 15122 14651 15430 14660
rect 15488 14414 15516 17614
rect 19444 17610 19472 27882
rect 19536 26790 19564 31214
rect 21192 30734 21220 31282
rect 21376 30938 21404 31282
rect 21364 30932 21416 30938
rect 21364 30874 21416 30880
rect 20812 30728 20864 30734
rect 20812 30670 20864 30676
rect 21180 30728 21232 30734
rect 21180 30670 21232 30676
rect 19846 30492 20154 30501
rect 19846 30490 19852 30492
rect 19908 30490 19932 30492
rect 19988 30490 20012 30492
rect 20068 30490 20092 30492
rect 20148 30490 20154 30492
rect 19908 30438 19910 30490
rect 20090 30438 20092 30490
rect 19846 30436 19852 30438
rect 19908 30436 19932 30438
rect 19988 30436 20012 30438
rect 20068 30436 20092 30438
rect 20148 30436 20154 30438
rect 19846 30427 20154 30436
rect 19846 29404 20154 29413
rect 19846 29402 19852 29404
rect 19908 29402 19932 29404
rect 19988 29402 20012 29404
rect 20068 29402 20092 29404
rect 20148 29402 20154 29404
rect 19908 29350 19910 29402
rect 20090 29350 20092 29402
rect 19846 29348 19852 29350
rect 19908 29348 19932 29350
rect 19988 29348 20012 29350
rect 20068 29348 20092 29350
rect 20148 29348 20154 29350
rect 19846 29339 20154 29348
rect 20720 28552 20772 28558
rect 20720 28494 20772 28500
rect 19846 28316 20154 28325
rect 19846 28314 19852 28316
rect 19908 28314 19932 28316
rect 19988 28314 20012 28316
rect 20068 28314 20092 28316
rect 20148 28314 20154 28316
rect 19908 28262 19910 28314
rect 20090 28262 20092 28314
rect 19846 28260 19852 28262
rect 19908 28260 19932 28262
rect 19988 28260 20012 28262
rect 20068 28260 20092 28262
rect 20148 28260 20154 28262
rect 19846 28251 20154 28260
rect 19708 27872 19760 27878
rect 19708 27814 19760 27820
rect 19524 26784 19576 26790
rect 19524 26726 19576 26732
rect 19536 24206 19564 26726
rect 19616 26308 19668 26314
rect 19616 26250 19668 26256
rect 19628 24818 19656 26250
rect 19720 25158 19748 27814
rect 20732 27402 20760 28494
rect 20720 27396 20772 27402
rect 20720 27338 20772 27344
rect 19846 27228 20154 27237
rect 19846 27226 19852 27228
rect 19908 27226 19932 27228
rect 19988 27226 20012 27228
rect 20068 27226 20092 27228
rect 20148 27226 20154 27228
rect 19908 27174 19910 27226
rect 20090 27174 20092 27226
rect 19846 27172 19852 27174
rect 19908 27172 19932 27174
rect 19988 27172 20012 27174
rect 20068 27172 20092 27174
rect 20148 27172 20154 27174
rect 19846 27163 20154 27172
rect 20732 26790 20760 27338
rect 20720 26784 20772 26790
rect 20720 26726 20772 26732
rect 19846 26140 20154 26149
rect 19846 26138 19852 26140
rect 19908 26138 19932 26140
rect 19988 26138 20012 26140
rect 20068 26138 20092 26140
rect 20148 26138 20154 26140
rect 19908 26086 19910 26138
rect 20090 26086 20092 26138
rect 19846 26084 19852 26086
rect 19908 26084 19932 26086
rect 19988 26084 20012 26086
rect 20068 26084 20092 26086
rect 20148 26084 20154 26086
rect 19846 26075 20154 26084
rect 20536 25288 20588 25294
rect 20536 25230 20588 25236
rect 19708 25152 19760 25158
rect 19708 25094 19760 25100
rect 19616 24812 19668 24818
rect 19616 24754 19668 24760
rect 19524 24200 19576 24206
rect 19524 24142 19576 24148
rect 17960 17604 18012 17610
rect 17960 17546 18012 17552
rect 19432 17604 19484 17610
rect 19432 17546 19484 17552
rect 17776 17536 17828 17542
rect 17776 17478 17828 17484
rect 17788 17338 17816 17478
rect 17776 17332 17828 17338
rect 17776 17274 17828 17280
rect 17788 17082 17816 17274
rect 17972 17202 18000 17546
rect 17960 17196 18012 17202
rect 17960 17138 18012 17144
rect 19064 17196 19116 17202
rect 19064 17138 19116 17144
rect 17696 17054 17816 17082
rect 16120 16720 16172 16726
rect 16120 16662 16172 16668
rect 15844 16516 15896 16522
rect 15844 16458 15896 16464
rect 15856 15638 15884 16458
rect 16132 15978 16160 16662
rect 16120 15972 16172 15978
rect 16120 15914 16172 15920
rect 15844 15632 15896 15638
rect 15844 15574 15896 15580
rect 15752 15496 15804 15502
rect 15752 15438 15804 15444
rect 15764 14958 15792 15438
rect 15752 14952 15804 14958
rect 15752 14894 15804 14900
rect 15764 14550 15792 14894
rect 15752 14544 15804 14550
rect 15752 14486 15804 14492
rect 15856 14482 15884 15574
rect 16132 15026 16160 15914
rect 17696 15026 17724 17054
rect 17776 16992 17828 16998
rect 17776 16934 17828 16940
rect 18788 16992 18840 16998
rect 18788 16934 18840 16940
rect 17788 16454 17816 16934
rect 17776 16448 17828 16454
rect 17776 16390 17828 16396
rect 18800 15162 18828 16934
rect 18788 15156 18840 15162
rect 18788 15098 18840 15104
rect 16120 15020 16172 15026
rect 16120 14962 16172 14968
rect 17684 15020 17736 15026
rect 17684 14962 17736 14968
rect 17500 14952 17552 14958
rect 17500 14894 17552 14900
rect 17512 14482 17540 14894
rect 15844 14476 15896 14482
rect 15844 14418 15896 14424
rect 17500 14476 17552 14482
rect 17500 14418 17552 14424
rect 15476 14408 15528 14414
rect 15476 14350 15528 14356
rect 17592 14408 17644 14414
rect 17592 14350 17644 14356
rect 15488 14006 15516 14350
rect 15476 14000 15528 14006
rect 15476 13942 15528 13948
rect 17604 13938 17632 14350
rect 17592 13932 17644 13938
rect 17592 13874 17644 13880
rect 15122 13628 15430 13637
rect 15122 13626 15128 13628
rect 15184 13626 15208 13628
rect 15264 13626 15288 13628
rect 15344 13626 15368 13628
rect 15424 13626 15430 13628
rect 15184 13574 15186 13626
rect 15366 13574 15368 13626
rect 15122 13572 15128 13574
rect 15184 13572 15208 13574
rect 15264 13572 15288 13574
rect 15344 13572 15368 13574
rect 15424 13572 15430 13574
rect 15122 13563 15430 13572
rect 16488 13388 16540 13394
rect 16488 13330 16540 13336
rect 14832 12640 14884 12646
rect 14832 12582 14884 12588
rect 14844 12374 14872 12582
rect 15122 12540 15430 12549
rect 15122 12538 15128 12540
rect 15184 12538 15208 12540
rect 15264 12538 15288 12540
rect 15344 12538 15368 12540
rect 15424 12538 15430 12540
rect 15184 12486 15186 12538
rect 15366 12486 15368 12538
rect 15122 12484 15128 12486
rect 15184 12484 15208 12486
rect 15264 12484 15288 12486
rect 15344 12484 15368 12486
rect 15424 12484 15430 12486
rect 15122 12475 15430 12484
rect 14832 12368 14884 12374
rect 14832 12310 14884 12316
rect 14740 11756 14792 11762
rect 14740 11698 14792 11704
rect 14844 11286 14872 12310
rect 16500 12170 16528 13330
rect 17696 13326 17724 14962
rect 18236 14000 18288 14006
rect 18236 13942 18288 13948
rect 18052 13796 18104 13802
rect 18052 13738 18104 13744
rect 17684 13320 17736 13326
rect 17684 13262 17736 13268
rect 18064 12782 18092 13738
rect 18052 12776 18104 12782
rect 18052 12718 18104 12724
rect 16488 12164 16540 12170
rect 16488 12106 16540 12112
rect 15122 11452 15430 11461
rect 15122 11450 15128 11452
rect 15184 11450 15208 11452
rect 15264 11450 15288 11452
rect 15344 11450 15368 11452
rect 15424 11450 15430 11452
rect 15184 11398 15186 11450
rect 15366 11398 15368 11450
rect 15122 11396 15128 11398
rect 15184 11396 15208 11398
rect 15264 11396 15288 11398
rect 15344 11396 15368 11398
rect 15424 11396 15430 11398
rect 15122 11387 15430 11396
rect 14832 11280 14884 11286
rect 14832 11222 14884 11228
rect 16500 11150 16528 12106
rect 18064 11762 18092 12718
rect 18248 11762 18276 13942
rect 18788 13184 18840 13190
rect 18788 13126 18840 13132
rect 18800 12918 18828 13126
rect 19076 12918 19104 17138
rect 19536 16574 19564 24142
rect 19628 20466 19656 24754
rect 19720 24274 19748 25094
rect 19846 25052 20154 25061
rect 19846 25050 19852 25052
rect 19908 25050 19932 25052
rect 19988 25050 20012 25052
rect 20068 25050 20092 25052
rect 20148 25050 20154 25052
rect 19908 24998 19910 25050
rect 20090 24998 20092 25050
rect 19846 24996 19852 24998
rect 19908 24996 19932 24998
rect 19988 24996 20012 24998
rect 20068 24996 20092 24998
rect 20148 24996 20154 24998
rect 19846 24987 20154 24996
rect 19708 24268 19760 24274
rect 19708 24210 19760 24216
rect 19846 23964 20154 23973
rect 19846 23962 19852 23964
rect 19908 23962 19932 23964
rect 19988 23962 20012 23964
rect 20068 23962 20092 23964
rect 20148 23962 20154 23964
rect 19908 23910 19910 23962
rect 20090 23910 20092 23962
rect 19846 23908 19852 23910
rect 19908 23908 19932 23910
rect 19988 23908 20012 23910
rect 20068 23908 20092 23910
rect 20148 23908 20154 23910
rect 19846 23899 20154 23908
rect 19846 22876 20154 22885
rect 19846 22874 19852 22876
rect 19908 22874 19932 22876
rect 19988 22874 20012 22876
rect 20068 22874 20092 22876
rect 20148 22874 20154 22876
rect 19908 22822 19910 22874
rect 20090 22822 20092 22874
rect 19846 22820 19852 22822
rect 19908 22820 19932 22822
rect 19988 22820 20012 22822
rect 20068 22820 20092 22822
rect 20148 22820 20154 22822
rect 19846 22811 20154 22820
rect 19846 21788 20154 21797
rect 19846 21786 19852 21788
rect 19908 21786 19932 21788
rect 19988 21786 20012 21788
rect 20068 21786 20092 21788
rect 20148 21786 20154 21788
rect 19908 21734 19910 21786
rect 20090 21734 20092 21786
rect 19846 21732 19852 21734
rect 19908 21732 19932 21734
rect 19988 21732 20012 21734
rect 20068 21732 20092 21734
rect 20148 21732 20154 21734
rect 19846 21723 20154 21732
rect 19708 21548 19760 21554
rect 19708 21490 19760 21496
rect 20352 21548 20404 21554
rect 20352 21490 20404 21496
rect 19720 20602 19748 21490
rect 20260 21344 20312 21350
rect 20260 21286 20312 21292
rect 20272 20942 20300 21286
rect 20260 20936 20312 20942
rect 20260 20878 20312 20884
rect 19846 20700 20154 20709
rect 19846 20698 19852 20700
rect 19908 20698 19932 20700
rect 19988 20698 20012 20700
rect 20068 20698 20092 20700
rect 20148 20698 20154 20700
rect 19908 20646 19910 20698
rect 20090 20646 20092 20698
rect 19846 20644 19852 20646
rect 19908 20644 19932 20646
rect 19988 20644 20012 20646
rect 20068 20644 20092 20646
rect 20148 20644 20154 20646
rect 19846 20635 20154 20644
rect 19708 20596 19760 20602
rect 19708 20538 19760 20544
rect 19616 20460 19668 20466
rect 19616 20402 19668 20408
rect 19628 17338 19656 20402
rect 20364 19786 20392 21490
rect 20548 19922 20576 25230
rect 20628 24064 20680 24070
rect 20628 24006 20680 24012
rect 20640 23730 20668 24006
rect 20628 23724 20680 23730
rect 20628 23666 20680 23672
rect 20824 22642 20852 30670
rect 21192 28626 21220 30670
rect 21180 28620 21232 28626
rect 21180 28562 21232 28568
rect 21272 28484 21324 28490
rect 21272 28426 21324 28432
rect 21284 28082 21312 28426
rect 20996 28076 21048 28082
rect 20996 28018 21048 28024
rect 21272 28076 21324 28082
rect 21272 28018 21324 28024
rect 21008 27674 21036 28018
rect 23492 28014 23520 31962
rect 25044 31816 25096 31822
rect 25044 31758 25096 31764
rect 25320 31816 25372 31822
rect 25320 31758 25372 31764
rect 24570 31036 24878 31045
rect 24570 31034 24576 31036
rect 24632 31034 24656 31036
rect 24712 31034 24736 31036
rect 24792 31034 24816 31036
rect 24872 31034 24878 31036
rect 24632 30982 24634 31034
rect 24814 30982 24816 31034
rect 24570 30980 24576 30982
rect 24632 30980 24656 30982
rect 24712 30980 24736 30982
rect 24792 30980 24816 30982
rect 24872 30980 24878 30982
rect 24570 30971 24878 30980
rect 25056 30938 25084 31758
rect 25332 30938 25360 31758
rect 25044 30932 25096 30938
rect 25044 30874 25096 30880
rect 25320 30932 25372 30938
rect 25320 30874 25372 30880
rect 23940 30796 23992 30802
rect 23940 30738 23992 30744
rect 23952 29714 23980 30738
rect 24492 30728 24544 30734
rect 24492 30670 24544 30676
rect 25228 30728 25280 30734
rect 25228 30670 25280 30676
rect 24400 30252 24452 30258
rect 24400 30194 24452 30200
rect 23940 29708 23992 29714
rect 23940 29650 23992 29656
rect 24124 29640 24176 29646
rect 24124 29582 24176 29588
rect 24136 28082 24164 29582
rect 24412 29306 24440 30194
rect 24504 30190 24532 30670
rect 24492 30184 24544 30190
rect 24492 30126 24544 30132
rect 24400 29300 24452 29306
rect 24400 29242 24452 29248
rect 24124 28076 24176 28082
rect 24124 28018 24176 28024
rect 23480 28008 23532 28014
rect 23480 27950 23532 27956
rect 20996 27668 21048 27674
rect 20996 27610 21048 27616
rect 23492 27606 23520 27950
rect 23480 27600 23532 27606
rect 23480 27542 23532 27548
rect 24136 27538 24164 28018
rect 24308 27872 24360 27878
rect 24308 27814 24360 27820
rect 24124 27532 24176 27538
rect 24124 27474 24176 27480
rect 24136 27130 24164 27474
rect 24124 27124 24176 27130
rect 24124 27066 24176 27072
rect 23572 26988 23624 26994
rect 23572 26930 23624 26936
rect 21272 26784 21324 26790
rect 21272 26726 21324 26732
rect 20996 25288 21048 25294
rect 20996 25230 21048 25236
rect 21008 24682 21036 25230
rect 20996 24676 21048 24682
rect 20996 24618 21048 24624
rect 21008 24274 21036 24618
rect 20996 24268 21048 24274
rect 20996 24210 21048 24216
rect 20904 23724 20956 23730
rect 20904 23666 20956 23672
rect 20812 22636 20864 22642
rect 20812 22578 20864 22584
rect 20916 21146 20944 23666
rect 20996 23520 21048 23526
rect 20996 23462 21048 23468
rect 20904 21140 20956 21146
rect 20904 21082 20956 21088
rect 21008 20806 21036 23462
rect 20996 20800 21048 20806
rect 20996 20742 21048 20748
rect 20536 19916 20588 19922
rect 20536 19858 20588 19864
rect 20352 19780 20404 19786
rect 20352 19722 20404 19728
rect 19846 19612 20154 19621
rect 19846 19610 19852 19612
rect 19908 19610 19932 19612
rect 19988 19610 20012 19612
rect 20068 19610 20092 19612
rect 20148 19610 20154 19612
rect 19908 19558 19910 19610
rect 20090 19558 20092 19610
rect 19846 19556 19852 19558
rect 19908 19556 19932 19558
rect 19988 19556 20012 19558
rect 20068 19556 20092 19558
rect 20148 19556 20154 19558
rect 19846 19547 20154 19556
rect 20904 18964 20956 18970
rect 20904 18906 20956 18912
rect 20628 18692 20680 18698
rect 20628 18634 20680 18640
rect 19846 18524 20154 18533
rect 19846 18522 19852 18524
rect 19908 18522 19932 18524
rect 19988 18522 20012 18524
rect 20068 18522 20092 18524
rect 20148 18522 20154 18524
rect 19908 18470 19910 18522
rect 20090 18470 20092 18522
rect 19846 18468 19852 18470
rect 19908 18468 19932 18470
rect 19988 18468 20012 18470
rect 20068 18468 20092 18470
rect 20148 18468 20154 18470
rect 19846 18459 20154 18468
rect 19846 17436 20154 17445
rect 19846 17434 19852 17436
rect 19908 17434 19932 17436
rect 19988 17434 20012 17436
rect 20068 17434 20092 17436
rect 20148 17434 20154 17436
rect 19908 17382 19910 17434
rect 20090 17382 20092 17434
rect 19846 17380 19852 17382
rect 19908 17380 19932 17382
rect 19988 17380 20012 17382
rect 20068 17380 20092 17382
rect 20148 17380 20154 17382
rect 19846 17371 20154 17380
rect 19616 17332 19668 17338
rect 19616 17274 19668 17280
rect 19800 17264 19852 17270
rect 19800 17206 19852 17212
rect 19812 16658 19840 17206
rect 19800 16652 19852 16658
rect 19800 16594 19852 16600
rect 19444 16546 19564 16574
rect 19340 14408 19392 14414
rect 19340 14350 19392 14356
rect 18788 12912 18840 12918
rect 18788 12854 18840 12860
rect 19064 12912 19116 12918
rect 19064 12854 19116 12860
rect 18052 11756 18104 11762
rect 18052 11698 18104 11704
rect 18236 11756 18288 11762
rect 18236 11698 18288 11704
rect 16672 11620 16724 11626
rect 16672 11562 16724 11568
rect 16684 11218 16712 11562
rect 18052 11552 18104 11558
rect 18052 11494 18104 11500
rect 16672 11212 16724 11218
rect 16672 11154 16724 11160
rect 14648 11144 14700 11150
rect 14648 11086 14700 11092
rect 16028 11144 16080 11150
rect 16028 11086 16080 11092
rect 16488 11144 16540 11150
rect 16488 11086 16540 11092
rect 14556 10736 14608 10742
rect 14556 10678 14608 10684
rect 15122 10364 15430 10373
rect 15122 10362 15128 10364
rect 15184 10362 15208 10364
rect 15264 10362 15288 10364
rect 15344 10362 15368 10364
rect 15424 10362 15430 10364
rect 15184 10310 15186 10362
rect 15366 10310 15368 10362
rect 15122 10308 15128 10310
rect 15184 10308 15208 10310
rect 15264 10308 15288 10310
rect 15344 10308 15368 10310
rect 15424 10308 15430 10310
rect 15122 10299 15430 10308
rect 16040 10130 16068 11086
rect 16672 11008 16724 11014
rect 16672 10950 16724 10956
rect 16684 10742 16712 10950
rect 18064 10810 18092 11494
rect 18052 10804 18104 10810
rect 18052 10746 18104 10752
rect 19076 10742 19104 12854
rect 19352 12850 19380 14350
rect 19340 12844 19392 12850
rect 19340 12786 19392 12792
rect 19444 12782 19472 16546
rect 19846 16348 20154 16357
rect 19846 16346 19852 16348
rect 19908 16346 19932 16348
rect 19988 16346 20012 16348
rect 20068 16346 20092 16348
rect 20148 16346 20154 16348
rect 19908 16294 19910 16346
rect 20090 16294 20092 16346
rect 19846 16292 19852 16294
rect 19908 16292 19932 16294
rect 19988 16292 20012 16294
rect 20068 16292 20092 16294
rect 20148 16292 20154 16294
rect 19846 16283 20154 16292
rect 20640 16250 20668 18634
rect 20916 16574 20944 18906
rect 20824 16546 20944 16574
rect 20628 16244 20680 16250
rect 20628 16186 20680 16192
rect 19846 15260 20154 15269
rect 19846 15258 19852 15260
rect 19908 15258 19932 15260
rect 19988 15258 20012 15260
rect 20068 15258 20092 15260
rect 20148 15258 20154 15260
rect 19908 15206 19910 15258
rect 20090 15206 20092 15258
rect 19846 15204 19852 15206
rect 19908 15204 19932 15206
rect 19988 15204 20012 15206
rect 20068 15204 20092 15206
rect 20148 15204 20154 15206
rect 19846 15195 20154 15204
rect 20720 14272 20772 14278
rect 20720 14214 20772 14220
rect 19846 14172 20154 14181
rect 19846 14170 19852 14172
rect 19908 14170 19932 14172
rect 19988 14170 20012 14172
rect 20068 14170 20092 14172
rect 20148 14170 20154 14172
rect 19908 14118 19910 14170
rect 20090 14118 20092 14170
rect 19846 14116 19852 14118
rect 19908 14116 19932 14118
rect 19988 14116 20012 14118
rect 20068 14116 20092 14118
rect 20148 14116 20154 14118
rect 19846 14107 20154 14116
rect 20732 13938 20760 14214
rect 20720 13932 20772 13938
rect 20720 13874 20772 13880
rect 19616 13388 19668 13394
rect 19616 13330 19668 13336
rect 19524 13320 19576 13326
rect 19524 13262 19576 13268
rect 19536 12986 19564 13262
rect 19524 12980 19576 12986
rect 19524 12922 19576 12928
rect 19432 12776 19484 12782
rect 19432 12718 19484 12724
rect 19628 12646 19656 13330
rect 19846 13084 20154 13093
rect 19846 13082 19852 13084
rect 19908 13082 19932 13084
rect 19988 13082 20012 13084
rect 20068 13082 20092 13084
rect 20148 13082 20154 13084
rect 19908 13030 19910 13082
rect 20090 13030 20092 13082
rect 19846 13028 19852 13030
rect 19908 13028 19932 13030
rect 19988 13028 20012 13030
rect 20068 13028 20092 13030
rect 20148 13028 20154 13030
rect 19846 13019 20154 13028
rect 19616 12640 19668 12646
rect 19616 12582 19668 12588
rect 16672 10736 16724 10742
rect 16672 10678 16724 10684
rect 17868 10736 17920 10742
rect 17868 10678 17920 10684
rect 19064 10736 19116 10742
rect 19064 10678 19116 10684
rect 16684 10130 16712 10678
rect 17592 10464 17644 10470
rect 17592 10406 17644 10412
rect 16028 10124 16080 10130
rect 16028 10066 16080 10072
rect 16672 10124 16724 10130
rect 16672 10066 16724 10072
rect 15122 9276 15430 9285
rect 15122 9274 15128 9276
rect 15184 9274 15208 9276
rect 15264 9274 15288 9276
rect 15344 9274 15368 9276
rect 15424 9274 15430 9276
rect 15184 9222 15186 9274
rect 15366 9222 15368 9274
rect 15122 9220 15128 9222
rect 15184 9220 15208 9222
rect 15264 9220 15288 9222
rect 15344 9220 15368 9222
rect 15424 9220 15430 9222
rect 15122 9211 15430 9220
rect 13820 8900 13872 8906
rect 13820 8842 13872 8848
rect 13832 8566 13860 8842
rect 13820 8560 13872 8566
rect 13820 8502 13872 8508
rect 13728 8492 13780 8498
rect 13728 8434 13780 8440
rect 13084 8288 13136 8294
rect 13084 8230 13136 8236
rect 13096 7818 13124 8230
rect 13740 7886 13768 8434
rect 17500 8424 17552 8430
rect 17500 8366 17552 8372
rect 15122 8188 15430 8197
rect 15122 8186 15128 8188
rect 15184 8186 15208 8188
rect 15264 8186 15288 8188
rect 15344 8186 15368 8188
rect 15424 8186 15430 8188
rect 15184 8134 15186 8186
rect 15366 8134 15368 8186
rect 15122 8132 15128 8134
rect 15184 8132 15208 8134
rect 15264 8132 15288 8134
rect 15344 8132 15368 8134
rect 15424 8132 15430 8134
rect 15122 8123 15430 8132
rect 13728 7880 13780 7886
rect 13728 7822 13780 7828
rect 13084 7812 13136 7818
rect 13084 7754 13136 7760
rect 14096 7744 14148 7750
rect 14096 7686 14148 7692
rect 14108 7410 14136 7686
rect 17408 7472 17460 7478
rect 17408 7414 17460 7420
rect 14096 7404 14148 7410
rect 14096 7346 14148 7352
rect 12164 7336 12216 7342
rect 12164 7278 12216 7284
rect 12992 7336 13044 7342
rect 12992 7278 13044 7284
rect 13004 7002 13032 7278
rect 15122 7100 15430 7109
rect 15122 7098 15128 7100
rect 15184 7098 15208 7100
rect 15264 7098 15288 7100
rect 15344 7098 15368 7100
rect 15424 7098 15430 7100
rect 15184 7046 15186 7098
rect 15366 7046 15368 7098
rect 15122 7044 15128 7046
rect 15184 7044 15208 7046
rect 15264 7044 15288 7046
rect 15344 7044 15368 7046
rect 15424 7044 15430 7046
rect 15122 7035 15430 7044
rect 12992 6996 13044 7002
rect 12992 6938 13044 6944
rect 17420 6934 17448 7414
rect 17512 6934 17540 8366
rect 17408 6928 17460 6934
rect 17408 6870 17460 6876
rect 17500 6928 17552 6934
rect 17500 6870 17552 6876
rect 15122 6012 15430 6021
rect 15122 6010 15128 6012
rect 15184 6010 15208 6012
rect 15264 6010 15288 6012
rect 15344 6010 15368 6012
rect 15424 6010 15430 6012
rect 15184 5958 15186 6010
rect 15366 5958 15368 6010
rect 15122 5956 15128 5958
rect 15184 5956 15208 5958
rect 15264 5956 15288 5958
rect 15344 5956 15368 5958
rect 15424 5956 15430 5958
rect 15122 5947 15430 5956
rect 15122 4924 15430 4933
rect 15122 4922 15128 4924
rect 15184 4922 15208 4924
rect 15264 4922 15288 4924
rect 15344 4922 15368 4924
rect 15424 4922 15430 4924
rect 15184 4870 15186 4922
rect 15366 4870 15368 4922
rect 15122 4868 15128 4870
rect 15184 4868 15208 4870
rect 15264 4868 15288 4870
rect 15344 4868 15368 4870
rect 15424 4868 15430 4870
rect 15122 4859 15430 4868
rect 14832 4616 14884 4622
rect 14832 4558 14884 4564
rect 14280 4480 14332 4486
rect 14280 4422 14332 4428
rect 14292 4146 14320 4422
rect 14280 4140 14332 4146
rect 14280 4082 14332 4088
rect 14372 4140 14424 4146
rect 14372 4082 14424 4088
rect 14464 4140 14516 4146
rect 14464 4082 14516 4088
rect 14188 4004 14240 4010
rect 14188 3946 14240 3952
rect 14200 3738 14228 3946
rect 14384 3942 14412 4082
rect 14372 3936 14424 3942
rect 14372 3878 14424 3884
rect 12072 3732 12124 3738
rect 12072 3674 12124 3680
rect 14188 3732 14240 3738
rect 14188 3674 14240 3680
rect 14384 3670 14412 3878
rect 11980 3664 12032 3670
rect 11980 3606 12032 3612
rect 14372 3664 14424 3670
rect 14372 3606 14424 3612
rect 14476 3602 14504 4082
rect 14464 3596 14516 3602
rect 14464 3538 14516 3544
rect 14648 3596 14700 3602
rect 14648 3538 14700 3544
rect 10784 3528 10836 3534
rect 10784 3470 10836 3476
rect 12440 3528 12492 3534
rect 12440 3470 12492 3476
rect 14372 3528 14424 3534
rect 14372 3470 14424 3476
rect 10398 3292 10706 3301
rect 10398 3290 10404 3292
rect 10460 3290 10484 3292
rect 10540 3290 10564 3292
rect 10620 3290 10644 3292
rect 10700 3290 10706 3292
rect 10460 3238 10462 3290
rect 10642 3238 10644 3290
rect 10398 3236 10404 3238
rect 10460 3236 10484 3238
rect 10540 3236 10564 3238
rect 10620 3236 10644 3238
rect 10700 3236 10706 3238
rect 10398 3227 10706 3236
rect 12452 3194 12480 3470
rect 14188 3460 14240 3466
rect 14188 3402 14240 3408
rect 12440 3188 12492 3194
rect 12440 3130 12492 3136
rect 12452 2446 12480 3130
rect 14200 2854 14228 3402
rect 14384 3126 14412 3470
rect 14556 3392 14608 3398
rect 14556 3334 14608 3340
rect 14568 3126 14596 3334
rect 14372 3120 14424 3126
rect 14372 3062 14424 3068
rect 14556 3120 14608 3126
rect 14556 3062 14608 3068
rect 12808 2848 12860 2854
rect 12808 2790 12860 2796
rect 14004 2848 14056 2854
rect 14004 2790 14056 2796
rect 14188 2848 14240 2854
rect 14188 2790 14240 2796
rect 12820 2446 12848 2790
rect 14016 2446 14044 2790
rect 14200 2650 14228 2790
rect 14384 2650 14412 3062
rect 14660 2990 14688 3538
rect 14648 2984 14700 2990
rect 14648 2926 14700 2932
rect 14188 2644 14240 2650
rect 14188 2586 14240 2592
rect 14372 2644 14424 2650
rect 14372 2586 14424 2592
rect 14844 2582 14872 4558
rect 15568 4480 15620 4486
rect 15568 4422 15620 4428
rect 15580 4078 15608 4422
rect 17512 4078 17540 6870
rect 15568 4072 15620 4078
rect 15568 4014 15620 4020
rect 17500 4072 17552 4078
rect 17500 4014 17552 4020
rect 14924 3936 14976 3942
rect 14924 3878 14976 3884
rect 14936 3126 14964 3878
rect 15122 3836 15430 3845
rect 15122 3834 15128 3836
rect 15184 3834 15208 3836
rect 15264 3834 15288 3836
rect 15344 3834 15368 3836
rect 15424 3834 15430 3836
rect 15184 3782 15186 3834
rect 15366 3782 15368 3834
rect 15122 3780 15128 3782
rect 15184 3780 15208 3782
rect 15264 3780 15288 3782
rect 15344 3780 15368 3782
rect 15424 3780 15430 3782
rect 15122 3771 15430 3780
rect 16764 3732 16816 3738
rect 16764 3674 16816 3680
rect 16672 3392 16724 3398
rect 16672 3334 16724 3340
rect 14924 3120 14976 3126
rect 14924 3062 14976 3068
rect 15122 2748 15430 2757
rect 15122 2746 15128 2748
rect 15184 2746 15208 2748
rect 15264 2746 15288 2748
rect 15344 2746 15368 2748
rect 15424 2746 15430 2748
rect 15184 2694 15186 2746
rect 15366 2694 15368 2746
rect 15122 2692 15128 2694
rect 15184 2692 15208 2694
rect 15264 2692 15288 2694
rect 15344 2692 15368 2694
rect 15424 2692 15430 2694
rect 15122 2683 15430 2692
rect 16684 2650 16712 3334
rect 16672 2644 16724 2650
rect 16672 2586 16724 2592
rect 16776 2582 16804 3674
rect 16856 3460 16908 3466
rect 16856 3402 16908 3408
rect 16868 2650 16896 3402
rect 17604 2990 17632 10406
rect 17880 8974 17908 10678
rect 18972 10668 19024 10674
rect 18972 10610 19024 10616
rect 18984 10470 19012 10610
rect 18972 10464 19024 10470
rect 18972 10406 19024 10412
rect 18984 9654 19012 10406
rect 18972 9648 19024 9654
rect 18972 9590 19024 9596
rect 17868 8968 17920 8974
rect 17868 8910 17920 8916
rect 18984 8634 19012 9590
rect 18972 8628 19024 8634
rect 18972 8570 19024 8576
rect 17776 8492 17828 8498
rect 17776 8434 17828 8440
rect 17788 6662 17816 8434
rect 18236 7948 18288 7954
rect 18236 7890 18288 7896
rect 18052 7812 18104 7818
rect 18052 7754 18104 7760
rect 18064 7206 18092 7754
rect 18248 7410 18276 7890
rect 18236 7404 18288 7410
rect 18236 7346 18288 7352
rect 17960 7200 18012 7206
rect 17960 7142 18012 7148
rect 18052 7200 18104 7206
rect 18052 7142 18104 7148
rect 17972 6798 18000 7142
rect 18064 6866 18092 7142
rect 18052 6860 18104 6866
rect 18052 6802 18104 6808
rect 17960 6792 18012 6798
rect 17960 6734 18012 6740
rect 17776 6656 17828 6662
rect 17776 6598 17828 6604
rect 18248 6390 18276 7346
rect 19524 6792 19576 6798
rect 19524 6734 19576 6740
rect 18328 6656 18380 6662
rect 18328 6598 18380 6604
rect 18236 6384 18288 6390
rect 18236 6326 18288 6332
rect 18340 4146 18368 6598
rect 19432 5296 19484 5302
rect 19432 5238 19484 5244
rect 19444 4826 19472 5238
rect 19536 5166 19564 6734
rect 19524 5160 19576 5166
rect 19524 5102 19576 5108
rect 19432 4820 19484 4826
rect 19432 4762 19484 4768
rect 19628 4434 19656 12582
rect 19846 11996 20154 12005
rect 19846 11994 19852 11996
rect 19908 11994 19932 11996
rect 19988 11994 20012 11996
rect 20068 11994 20092 11996
rect 20148 11994 20154 11996
rect 19908 11942 19910 11994
rect 20090 11942 20092 11994
rect 19846 11940 19852 11942
rect 19908 11940 19932 11942
rect 19988 11940 20012 11942
rect 20068 11940 20092 11942
rect 20148 11940 20154 11942
rect 19846 11931 20154 11940
rect 19846 10908 20154 10917
rect 19846 10906 19852 10908
rect 19908 10906 19932 10908
rect 19988 10906 20012 10908
rect 20068 10906 20092 10908
rect 20148 10906 20154 10908
rect 19908 10854 19910 10906
rect 20090 10854 20092 10906
rect 19846 10852 19852 10854
rect 19908 10852 19932 10854
rect 19988 10852 20012 10854
rect 20068 10852 20092 10854
rect 20148 10852 20154 10854
rect 19846 10843 20154 10852
rect 20824 9994 20852 16546
rect 20904 14000 20956 14006
rect 20904 13942 20956 13948
rect 20916 13258 20944 13942
rect 20904 13252 20956 13258
rect 20904 13194 20956 13200
rect 21008 13190 21036 20742
rect 21088 16652 21140 16658
rect 21088 16594 21140 16600
rect 21100 14006 21128 16594
rect 21180 16516 21232 16522
rect 21180 16458 21232 16464
rect 21088 14000 21140 14006
rect 21088 13942 21140 13948
rect 21192 13802 21220 16458
rect 21180 13796 21232 13802
rect 21180 13738 21232 13744
rect 21192 13530 21220 13738
rect 21284 13530 21312 26726
rect 21824 26376 21876 26382
rect 21824 26318 21876 26324
rect 21836 25498 21864 26318
rect 22836 25696 22888 25702
rect 22836 25638 22888 25644
rect 21824 25492 21876 25498
rect 21824 25434 21876 25440
rect 21836 25362 21864 25434
rect 21824 25356 21876 25362
rect 21824 25298 21876 25304
rect 21836 25242 21864 25298
rect 21744 25214 21864 25242
rect 22100 25288 22152 25294
rect 22100 25230 22152 25236
rect 21744 23730 21772 25214
rect 21824 25152 21876 25158
rect 21824 25094 21876 25100
rect 21836 24818 21864 25094
rect 21824 24812 21876 24818
rect 21824 24754 21876 24760
rect 22112 24614 22140 25230
rect 22848 25158 22876 25638
rect 22836 25152 22888 25158
rect 22836 25094 22888 25100
rect 22100 24608 22152 24614
rect 22100 24550 22152 24556
rect 21732 23724 21784 23730
rect 21732 23666 21784 23672
rect 22848 23526 22876 25094
rect 22836 23520 22888 23526
rect 22836 23462 22888 23468
rect 23480 22092 23532 22098
rect 23480 22034 23532 22040
rect 23492 21690 23520 22034
rect 23480 21684 23532 21690
rect 23480 21626 23532 21632
rect 23584 21570 23612 26930
rect 23664 22024 23716 22030
rect 23664 21966 23716 21972
rect 23676 21690 23704 21966
rect 23664 21684 23716 21690
rect 23664 21626 23716 21632
rect 23492 21554 23612 21570
rect 23480 21548 23612 21554
rect 23532 21542 23612 21548
rect 23480 21490 23532 21496
rect 23388 21480 23440 21486
rect 23388 21422 23440 21428
rect 22928 20528 22980 20534
rect 22928 20470 22980 20476
rect 22008 19712 22060 19718
rect 22008 19654 22060 19660
rect 22020 19378 22048 19654
rect 22008 19372 22060 19378
rect 22008 19314 22060 19320
rect 21640 19168 21692 19174
rect 21640 19110 21692 19116
rect 21652 18766 21680 19110
rect 21640 18760 21692 18766
rect 21640 18702 21692 18708
rect 22100 17536 22152 17542
rect 22100 17478 22152 17484
rect 22112 17270 22140 17478
rect 22100 17264 22152 17270
rect 22100 17206 22152 17212
rect 22284 17264 22336 17270
rect 22284 17206 22336 17212
rect 21456 16992 21508 16998
rect 21456 16934 21508 16940
rect 21468 16454 21496 16934
rect 22112 16522 22140 17206
rect 22296 16726 22324 17206
rect 22284 16720 22336 16726
rect 22284 16662 22336 16668
rect 22836 16652 22888 16658
rect 22836 16594 22888 16600
rect 22100 16516 22152 16522
rect 22100 16458 22152 16464
rect 22284 16516 22336 16522
rect 22284 16458 22336 16464
rect 21456 16448 21508 16454
rect 21456 16390 21508 16396
rect 21824 16448 21876 16454
rect 21824 16390 21876 16396
rect 21836 14482 21864 16390
rect 22008 15020 22060 15026
rect 22008 14962 22060 14968
rect 21824 14476 21876 14482
rect 21824 14418 21876 14424
rect 21916 14272 21968 14278
rect 21916 14214 21968 14220
rect 21824 14000 21876 14006
rect 21824 13942 21876 13948
rect 21836 13870 21864 13942
rect 21824 13864 21876 13870
rect 21824 13806 21876 13812
rect 21928 13734 21956 14214
rect 22020 14074 22048 14962
rect 22192 14408 22244 14414
rect 22192 14350 22244 14356
rect 22204 14074 22232 14350
rect 22008 14068 22060 14074
rect 22008 14010 22060 14016
rect 22192 14068 22244 14074
rect 22192 14010 22244 14016
rect 21916 13728 21968 13734
rect 21916 13670 21968 13676
rect 21180 13524 21232 13530
rect 21180 13466 21232 13472
rect 21272 13524 21324 13530
rect 21272 13466 21324 13472
rect 21928 13326 21956 13670
rect 21916 13320 21968 13326
rect 21916 13262 21968 13268
rect 20996 13184 21048 13190
rect 20996 13126 21048 13132
rect 21916 13184 21968 13190
rect 21916 13126 21968 13132
rect 21928 12986 21956 13126
rect 21916 12980 21968 12986
rect 21916 12922 21968 12928
rect 22020 12850 22048 14010
rect 22204 13326 22232 14010
rect 22296 13870 22324 16458
rect 22468 14476 22520 14482
rect 22468 14418 22520 14424
rect 22480 13988 22508 14418
rect 22848 14278 22876 16594
rect 22836 14272 22888 14278
rect 22836 14214 22888 14220
rect 22560 14000 22612 14006
rect 22480 13960 22560 13988
rect 22284 13864 22336 13870
rect 22284 13806 22336 13812
rect 22480 13326 22508 13960
rect 22560 13942 22612 13948
rect 22192 13320 22244 13326
rect 22192 13262 22244 13268
rect 22468 13320 22520 13326
rect 22468 13262 22520 13268
rect 22204 12918 22232 13262
rect 22192 12912 22244 12918
rect 22192 12854 22244 12860
rect 22008 12844 22060 12850
rect 22008 12786 22060 12792
rect 22468 12640 22520 12646
rect 22468 12582 22520 12588
rect 22480 10742 22508 12582
rect 22940 10810 22968 20470
rect 23400 20398 23428 21422
rect 23388 20392 23440 20398
rect 23388 20334 23440 20340
rect 23400 18834 23428 20334
rect 23388 18828 23440 18834
rect 23388 18770 23440 18776
rect 23492 16794 23520 21490
rect 23572 17672 23624 17678
rect 23572 17614 23624 17620
rect 23480 16788 23532 16794
rect 23480 16730 23532 16736
rect 23480 16652 23532 16658
rect 23480 16594 23532 16600
rect 23492 15026 23520 16594
rect 23584 16590 23612 17614
rect 23572 16584 23624 16590
rect 23572 16526 23624 16532
rect 23480 15020 23532 15026
rect 23480 14962 23532 14968
rect 23584 14006 23612 16526
rect 23664 16516 23716 16522
rect 23664 16458 23716 16464
rect 23676 14482 23704 16458
rect 24320 15978 24348 27814
rect 24504 26234 24532 30126
rect 24570 29948 24878 29957
rect 24570 29946 24576 29948
rect 24632 29946 24656 29948
rect 24712 29946 24736 29948
rect 24792 29946 24816 29948
rect 24872 29946 24878 29948
rect 24632 29894 24634 29946
rect 24814 29894 24816 29946
rect 24570 29892 24576 29894
rect 24632 29892 24656 29894
rect 24712 29892 24736 29894
rect 24792 29892 24816 29894
rect 24872 29892 24878 29894
rect 24570 29883 24878 29892
rect 25240 29850 25268 30670
rect 25424 30054 25452 31962
rect 28264 31816 28316 31822
rect 28264 31758 28316 31764
rect 28172 31748 28224 31754
rect 28172 31690 28224 31696
rect 28184 31278 28212 31690
rect 28172 31272 28224 31278
rect 28172 31214 28224 31220
rect 25412 30048 25464 30054
rect 25412 29990 25464 29996
rect 25228 29844 25280 29850
rect 25228 29786 25280 29792
rect 24768 29708 24820 29714
rect 24768 29650 24820 29656
rect 24780 29578 24808 29650
rect 24768 29572 24820 29578
rect 24768 29514 24820 29520
rect 24952 29164 25004 29170
rect 24952 29106 25004 29112
rect 24570 28860 24878 28869
rect 24570 28858 24576 28860
rect 24632 28858 24656 28860
rect 24712 28858 24736 28860
rect 24792 28858 24816 28860
rect 24872 28858 24878 28860
rect 24632 28806 24634 28858
rect 24814 28806 24816 28858
rect 24570 28804 24576 28806
rect 24632 28804 24656 28806
rect 24712 28804 24736 28806
rect 24792 28804 24816 28806
rect 24872 28804 24878 28806
rect 24570 28795 24878 28804
rect 24964 28218 24992 29106
rect 24952 28212 25004 28218
rect 24952 28154 25004 28160
rect 24570 27772 24878 27781
rect 24570 27770 24576 27772
rect 24632 27770 24656 27772
rect 24712 27770 24736 27772
rect 24792 27770 24816 27772
rect 24872 27770 24878 27772
rect 24632 27718 24634 27770
rect 24814 27718 24816 27770
rect 24570 27716 24576 27718
rect 24632 27716 24656 27718
rect 24712 27716 24736 27718
rect 24792 27716 24816 27718
rect 24872 27716 24878 27718
rect 24570 27707 24878 27716
rect 24952 27396 25004 27402
rect 24952 27338 25004 27344
rect 24570 26684 24878 26693
rect 24570 26682 24576 26684
rect 24632 26682 24656 26684
rect 24712 26682 24736 26684
rect 24792 26682 24816 26684
rect 24872 26682 24878 26684
rect 24632 26630 24634 26682
rect 24814 26630 24816 26682
rect 24570 26628 24576 26630
rect 24632 26628 24656 26630
rect 24712 26628 24736 26630
rect 24792 26628 24816 26630
rect 24872 26628 24878 26630
rect 24570 26619 24878 26628
rect 24860 26376 24912 26382
rect 24860 26318 24912 26324
rect 24412 26206 24532 26234
rect 24412 22098 24440 26206
rect 24872 26042 24900 26318
rect 24860 26036 24912 26042
rect 24860 25978 24912 25984
rect 24570 25596 24878 25605
rect 24570 25594 24576 25596
rect 24632 25594 24656 25596
rect 24712 25594 24736 25596
rect 24792 25594 24816 25596
rect 24872 25594 24878 25596
rect 24632 25542 24634 25594
rect 24814 25542 24816 25594
rect 24570 25540 24576 25542
rect 24632 25540 24656 25542
rect 24712 25540 24736 25542
rect 24792 25540 24816 25542
rect 24872 25540 24878 25542
rect 24570 25531 24878 25540
rect 24570 24508 24878 24517
rect 24570 24506 24576 24508
rect 24632 24506 24656 24508
rect 24712 24506 24736 24508
rect 24792 24506 24816 24508
rect 24872 24506 24878 24508
rect 24632 24454 24634 24506
rect 24814 24454 24816 24506
rect 24570 24452 24576 24454
rect 24632 24452 24656 24454
rect 24712 24452 24736 24454
rect 24792 24452 24816 24454
rect 24872 24452 24878 24454
rect 24570 24443 24878 24452
rect 24570 23420 24878 23429
rect 24570 23418 24576 23420
rect 24632 23418 24656 23420
rect 24712 23418 24736 23420
rect 24792 23418 24816 23420
rect 24872 23418 24878 23420
rect 24632 23366 24634 23418
rect 24814 23366 24816 23418
rect 24570 23364 24576 23366
rect 24632 23364 24656 23366
rect 24712 23364 24736 23366
rect 24792 23364 24816 23366
rect 24872 23364 24878 23366
rect 24570 23355 24878 23364
rect 24570 22332 24878 22341
rect 24570 22330 24576 22332
rect 24632 22330 24656 22332
rect 24712 22330 24736 22332
rect 24792 22330 24816 22332
rect 24872 22330 24878 22332
rect 24632 22278 24634 22330
rect 24814 22278 24816 22330
rect 24570 22276 24576 22278
rect 24632 22276 24656 22278
rect 24712 22276 24736 22278
rect 24792 22276 24816 22278
rect 24872 22276 24878 22278
rect 24570 22267 24878 22276
rect 24400 22092 24452 22098
rect 24400 22034 24452 22040
rect 24570 21244 24878 21253
rect 24570 21242 24576 21244
rect 24632 21242 24656 21244
rect 24712 21242 24736 21244
rect 24792 21242 24816 21244
rect 24872 21242 24878 21244
rect 24632 21190 24634 21242
rect 24814 21190 24816 21242
rect 24570 21188 24576 21190
rect 24632 21188 24656 21190
rect 24712 21188 24736 21190
rect 24792 21188 24816 21190
rect 24872 21188 24878 21190
rect 24570 21179 24878 21188
rect 24570 20156 24878 20165
rect 24570 20154 24576 20156
rect 24632 20154 24656 20156
rect 24712 20154 24736 20156
rect 24792 20154 24816 20156
rect 24872 20154 24878 20156
rect 24632 20102 24634 20154
rect 24814 20102 24816 20154
rect 24570 20100 24576 20102
rect 24632 20100 24656 20102
rect 24712 20100 24736 20102
rect 24792 20100 24816 20102
rect 24872 20100 24878 20102
rect 24570 20091 24878 20100
rect 24570 19068 24878 19077
rect 24570 19066 24576 19068
rect 24632 19066 24656 19068
rect 24712 19066 24736 19068
rect 24792 19066 24816 19068
rect 24872 19066 24878 19068
rect 24632 19014 24634 19066
rect 24814 19014 24816 19066
rect 24570 19012 24576 19014
rect 24632 19012 24656 19014
rect 24712 19012 24736 19014
rect 24792 19012 24816 19014
rect 24872 19012 24878 19014
rect 24570 19003 24878 19012
rect 24492 18760 24544 18766
rect 24492 18702 24544 18708
rect 24504 17678 24532 18702
rect 24570 17980 24878 17989
rect 24570 17978 24576 17980
rect 24632 17978 24656 17980
rect 24712 17978 24736 17980
rect 24792 17978 24816 17980
rect 24872 17978 24878 17980
rect 24632 17926 24634 17978
rect 24814 17926 24816 17978
rect 24570 17924 24576 17926
rect 24632 17924 24656 17926
rect 24712 17924 24736 17926
rect 24792 17924 24816 17926
rect 24872 17924 24878 17926
rect 24570 17915 24878 17924
rect 24492 17672 24544 17678
rect 24492 17614 24544 17620
rect 24570 16892 24878 16901
rect 24570 16890 24576 16892
rect 24632 16890 24656 16892
rect 24712 16890 24736 16892
rect 24792 16890 24816 16892
rect 24872 16890 24878 16892
rect 24632 16838 24634 16890
rect 24814 16838 24816 16890
rect 24570 16836 24576 16838
rect 24632 16836 24656 16838
rect 24712 16836 24736 16838
rect 24792 16836 24816 16838
rect 24872 16836 24878 16838
rect 24570 16827 24878 16836
rect 24492 16040 24544 16046
rect 24492 15982 24544 15988
rect 24308 15972 24360 15978
rect 24308 15914 24360 15920
rect 23664 14476 23716 14482
rect 23664 14418 23716 14424
rect 23676 14074 23704 14418
rect 23664 14068 23716 14074
rect 23664 14010 23716 14016
rect 23572 14000 23624 14006
rect 23572 13942 23624 13948
rect 24320 13462 24348 15914
rect 24504 15434 24532 15982
rect 24570 15804 24878 15813
rect 24570 15802 24576 15804
rect 24632 15802 24656 15804
rect 24712 15802 24736 15804
rect 24792 15802 24816 15804
rect 24872 15802 24878 15804
rect 24632 15750 24634 15802
rect 24814 15750 24816 15802
rect 24570 15748 24576 15750
rect 24632 15748 24656 15750
rect 24712 15748 24736 15750
rect 24792 15748 24816 15750
rect 24872 15748 24878 15750
rect 24570 15739 24878 15748
rect 24964 15706 24992 27338
rect 25044 26240 25096 26246
rect 25044 26182 25096 26188
rect 25056 25906 25084 26182
rect 25044 25900 25096 25906
rect 25044 25842 25096 25848
rect 25320 25832 25372 25838
rect 25320 25774 25372 25780
rect 25332 25294 25360 25774
rect 25320 25288 25372 25294
rect 25320 25230 25372 25236
rect 25424 21894 25452 29990
rect 28184 28082 28212 31214
rect 28276 30938 28304 31758
rect 29012 31482 29040 31962
rect 29294 31580 29602 31589
rect 29294 31578 29300 31580
rect 29356 31578 29380 31580
rect 29436 31578 29460 31580
rect 29516 31578 29540 31580
rect 29596 31578 29602 31580
rect 29356 31526 29358 31578
rect 29538 31526 29540 31578
rect 29294 31524 29300 31526
rect 29356 31524 29380 31526
rect 29436 31524 29460 31526
rect 29516 31524 29540 31526
rect 29596 31524 29602 31526
rect 29294 31515 29602 31524
rect 29000 31476 29052 31482
rect 29000 31418 29052 31424
rect 28264 30932 28316 30938
rect 28264 30874 28316 30880
rect 28816 30728 28868 30734
rect 28816 30670 28868 30676
rect 28828 29850 28856 30670
rect 28816 29844 28868 29850
rect 28816 29786 28868 29792
rect 28908 29640 28960 29646
rect 28908 29582 28960 29588
rect 28920 29170 28948 29582
rect 28908 29164 28960 29170
rect 28908 29106 28960 29112
rect 29012 28218 29040 31418
rect 29552 31340 29604 31346
rect 29552 31282 29604 31288
rect 29564 30938 29592 31282
rect 34018 31036 34326 31045
rect 34018 31034 34024 31036
rect 34080 31034 34104 31036
rect 34160 31034 34184 31036
rect 34240 31034 34264 31036
rect 34320 31034 34326 31036
rect 34080 30982 34082 31034
rect 34262 30982 34264 31034
rect 34018 30980 34024 30982
rect 34080 30980 34104 30982
rect 34160 30980 34184 30982
rect 34240 30980 34264 30982
rect 34320 30980 34326 30982
rect 34018 30971 34326 30980
rect 29552 30932 29604 30938
rect 29552 30874 29604 30880
rect 29736 30728 29788 30734
rect 29736 30670 29788 30676
rect 29294 30492 29602 30501
rect 29294 30490 29300 30492
rect 29356 30490 29380 30492
rect 29436 30490 29460 30492
rect 29516 30490 29540 30492
rect 29596 30490 29602 30492
rect 29356 30438 29358 30490
rect 29538 30438 29540 30490
rect 29294 30436 29300 30438
rect 29356 30436 29380 30438
rect 29436 30436 29460 30438
rect 29516 30436 29540 30438
rect 29596 30436 29602 30438
rect 29294 30427 29602 30436
rect 29294 29404 29602 29413
rect 29294 29402 29300 29404
rect 29356 29402 29380 29404
rect 29436 29402 29460 29404
rect 29516 29402 29540 29404
rect 29596 29402 29602 29404
rect 29356 29350 29358 29402
rect 29538 29350 29540 29402
rect 29294 29348 29300 29350
rect 29356 29348 29380 29350
rect 29436 29348 29460 29350
rect 29516 29348 29540 29350
rect 29596 29348 29602 29350
rect 29294 29339 29602 29348
rect 29748 29306 29776 30670
rect 34018 29948 34326 29957
rect 34018 29946 34024 29948
rect 34080 29946 34104 29948
rect 34160 29946 34184 29948
rect 34240 29946 34264 29948
rect 34320 29946 34326 29948
rect 34080 29894 34082 29946
rect 34262 29894 34264 29946
rect 34018 29892 34024 29894
rect 34080 29892 34104 29894
rect 34160 29892 34184 29894
rect 34240 29892 34264 29894
rect 34320 29892 34326 29894
rect 34018 29883 34326 29892
rect 31392 29572 31444 29578
rect 31392 29514 31444 29520
rect 31404 29306 31432 29514
rect 32680 29504 32732 29510
rect 32680 29446 32732 29452
rect 32692 29306 32720 29446
rect 29736 29300 29788 29306
rect 29736 29242 29788 29248
rect 31392 29300 31444 29306
rect 31392 29242 31444 29248
rect 32680 29300 32732 29306
rect 32680 29242 32732 29248
rect 34796 29300 34848 29306
rect 34796 29242 34848 29248
rect 31300 29164 31352 29170
rect 31300 29106 31352 29112
rect 31208 29096 31260 29102
rect 31208 29038 31260 29044
rect 29294 28316 29602 28325
rect 29294 28314 29300 28316
rect 29356 28314 29380 28316
rect 29436 28314 29460 28316
rect 29516 28314 29540 28316
rect 29596 28314 29602 28316
rect 29356 28262 29358 28314
rect 29538 28262 29540 28314
rect 29294 28260 29300 28262
rect 29356 28260 29380 28262
rect 29436 28260 29460 28262
rect 29516 28260 29540 28262
rect 29596 28260 29602 28262
rect 29294 28251 29602 28260
rect 29000 28212 29052 28218
rect 29000 28154 29052 28160
rect 28172 28076 28224 28082
rect 28172 28018 28224 28024
rect 28448 28076 28500 28082
rect 28448 28018 28500 28024
rect 28460 27130 28488 28018
rect 31220 28014 31248 29038
rect 31312 28490 31340 29106
rect 31300 28484 31352 28490
rect 31300 28426 31352 28432
rect 31208 28008 31260 28014
rect 31208 27950 31260 27956
rect 28540 27464 28592 27470
rect 28540 27406 28592 27412
rect 28448 27124 28500 27130
rect 28448 27066 28500 27072
rect 25964 25900 26016 25906
rect 25964 25842 26016 25848
rect 28448 25900 28500 25906
rect 28448 25842 28500 25848
rect 25976 25226 26004 25842
rect 27712 25764 27764 25770
rect 27712 25706 27764 25712
rect 27724 25226 27752 25706
rect 27804 25696 27856 25702
rect 27804 25638 27856 25644
rect 27816 25294 27844 25638
rect 27804 25288 27856 25294
rect 27804 25230 27856 25236
rect 25964 25220 26016 25226
rect 25964 25162 26016 25168
rect 27712 25220 27764 25226
rect 27712 25162 27764 25168
rect 25976 24818 26004 25162
rect 25964 24812 26016 24818
rect 25964 24754 26016 24760
rect 25872 23860 25924 23866
rect 25872 23802 25924 23808
rect 25688 22636 25740 22642
rect 25688 22578 25740 22584
rect 25412 21888 25464 21894
rect 25412 21830 25464 21836
rect 25136 21548 25188 21554
rect 25136 21490 25188 21496
rect 25044 19780 25096 19786
rect 25044 19722 25096 19728
rect 25056 17678 25084 19722
rect 25044 17672 25096 17678
rect 25044 17614 25096 17620
rect 25148 17338 25176 21490
rect 25424 20874 25452 21830
rect 25700 21690 25728 22578
rect 25884 22030 25912 23802
rect 27724 23662 27752 25162
rect 28460 24954 28488 25842
rect 28448 24948 28500 24954
rect 28448 24890 28500 24896
rect 28552 24274 28580 27406
rect 28724 27328 28776 27334
rect 28724 27270 28776 27276
rect 28736 26994 28764 27270
rect 29294 27228 29602 27237
rect 29294 27226 29300 27228
rect 29356 27226 29380 27228
rect 29436 27226 29460 27228
rect 29516 27226 29540 27228
rect 29596 27226 29602 27228
rect 29356 27174 29358 27226
rect 29538 27174 29540 27226
rect 29294 27172 29300 27174
rect 29356 27172 29380 27174
rect 29436 27172 29460 27174
rect 29516 27172 29540 27174
rect 29596 27172 29602 27174
rect 29294 27163 29602 27172
rect 28724 26988 28776 26994
rect 28724 26930 28776 26936
rect 30656 26988 30708 26994
rect 30656 26930 30708 26936
rect 29294 26140 29602 26149
rect 29294 26138 29300 26140
rect 29356 26138 29380 26140
rect 29436 26138 29460 26140
rect 29516 26138 29540 26140
rect 29596 26138 29602 26140
rect 29356 26086 29358 26138
rect 29538 26086 29540 26138
rect 29294 26084 29300 26086
rect 29356 26084 29380 26086
rect 29436 26084 29460 26086
rect 29516 26084 29540 26086
rect 29596 26084 29602 26086
rect 29294 26075 29602 26084
rect 30668 25838 30696 26930
rect 30656 25832 30708 25838
rect 30656 25774 30708 25780
rect 28724 25152 28776 25158
rect 28724 25094 28776 25100
rect 28632 24812 28684 24818
rect 28632 24754 28684 24760
rect 28540 24268 28592 24274
rect 28540 24210 28592 24216
rect 28644 24206 28672 24754
rect 28632 24200 28684 24206
rect 28632 24142 28684 24148
rect 28540 24132 28592 24138
rect 28540 24074 28592 24080
rect 28552 23866 28580 24074
rect 28736 23866 28764 25094
rect 29294 25052 29602 25061
rect 29294 25050 29300 25052
rect 29356 25050 29380 25052
rect 29436 25050 29460 25052
rect 29516 25050 29540 25052
rect 29596 25050 29602 25052
rect 29356 24998 29358 25050
rect 29538 24998 29540 25050
rect 29294 24996 29300 24998
rect 29356 24996 29380 24998
rect 29436 24996 29460 24998
rect 29516 24996 29540 24998
rect 29596 24996 29602 24998
rect 29294 24987 29602 24996
rect 30564 24676 30616 24682
rect 30564 24618 30616 24624
rect 30576 24070 30604 24618
rect 28816 24064 28868 24070
rect 28816 24006 28868 24012
rect 30564 24064 30616 24070
rect 30564 24006 30616 24012
rect 28540 23860 28592 23866
rect 28540 23802 28592 23808
rect 28724 23860 28776 23866
rect 28724 23802 28776 23808
rect 28828 23730 28856 24006
rect 29294 23964 29602 23973
rect 29294 23962 29300 23964
rect 29356 23962 29380 23964
rect 29436 23962 29460 23964
rect 29516 23962 29540 23964
rect 29596 23962 29602 23964
rect 29356 23910 29358 23962
rect 29538 23910 29540 23962
rect 29294 23908 29300 23910
rect 29356 23908 29380 23910
rect 29436 23908 29460 23910
rect 29516 23908 29540 23910
rect 29596 23908 29602 23910
rect 29294 23899 29602 23908
rect 28816 23724 28868 23730
rect 28816 23666 28868 23672
rect 27712 23656 27764 23662
rect 27712 23598 27764 23604
rect 26240 22432 26292 22438
rect 26240 22374 26292 22380
rect 26252 22030 26280 22374
rect 25872 22024 25924 22030
rect 25872 21966 25924 21972
rect 26240 22024 26292 22030
rect 26240 21966 26292 21972
rect 27068 22024 27120 22030
rect 27068 21966 27120 21972
rect 25688 21684 25740 21690
rect 25688 21626 25740 21632
rect 25412 20868 25464 20874
rect 25412 20810 25464 20816
rect 25412 18760 25464 18766
rect 25412 18702 25464 18708
rect 25228 18624 25280 18630
rect 25228 18566 25280 18572
rect 25240 18290 25268 18566
rect 25424 18426 25452 18702
rect 25412 18420 25464 18426
rect 25412 18362 25464 18368
rect 25228 18284 25280 18290
rect 25228 18226 25280 18232
rect 25136 17332 25188 17338
rect 25136 17274 25188 17280
rect 25884 16250 25912 21966
rect 25964 19372 26016 19378
rect 25964 19314 26016 19320
rect 25976 18698 26004 19314
rect 26240 19236 26292 19242
rect 26240 19178 26292 19184
rect 25964 18692 26016 18698
rect 25964 18634 26016 18640
rect 25872 16244 25924 16250
rect 25872 16186 25924 16192
rect 26252 16182 26280 19178
rect 26332 17672 26384 17678
rect 26332 17614 26384 17620
rect 26976 17672 27028 17678
rect 26976 17614 27028 17620
rect 26240 16176 26292 16182
rect 26240 16118 26292 16124
rect 25136 16108 25188 16114
rect 25136 16050 25188 16056
rect 24952 15700 25004 15706
rect 24952 15642 25004 15648
rect 24492 15428 24544 15434
rect 24492 15370 24544 15376
rect 24504 14890 24532 15370
rect 24492 14884 24544 14890
rect 24492 14826 24544 14832
rect 24308 13456 24360 13462
rect 24308 13398 24360 13404
rect 23756 13184 23808 13190
rect 23756 13126 23808 13132
rect 23768 12850 23796 13126
rect 23756 12844 23808 12850
rect 23756 12786 23808 12792
rect 24504 11082 24532 14826
rect 24570 14716 24878 14725
rect 24570 14714 24576 14716
rect 24632 14714 24656 14716
rect 24712 14714 24736 14716
rect 24792 14714 24816 14716
rect 24872 14714 24878 14716
rect 24632 14662 24634 14714
rect 24814 14662 24816 14714
rect 24570 14660 24576 14662
rect 24632 14660 24656 14662
rect 24712 14660 24736 14662
rect 24792 14660 24816 14662
rect 24872 14660 24878 14662
rect 24570 14651 24878 14660
rect 24570 13628 24878 13637
rect 24570 13626 24576 13628
rect 24632 13626 24656 13628
rect 24712 13626 24736 13628
rect 24792 13626 24816 13628
rect 24872 13626 24878 13628
rect 24632 13574 24634 13626
rect 24814 13574 24816 13626
rect 24570 13572 24576 13574
rect 24632 13572 24656 13574
rect 24712 13572 24736 13574
rect 24792 13572 24816 13574
rect 24872 13572 24878 13574
rect 24570 13563 24878 13572
rect 25148 13326 25176 16050
rect 26252 15570 26280 16118
rect 26344 16114 26372 17614
rect 26988 17338 27016 17614
rect 26976 17332 27028 17338
rect 26976 17274 27028 17280
rect 26332 16108 26384 16114
rect 26332 16050 26384 16056
rect 27080 15638 27108 21966
rect 27528 20460 27580 20466
rect 27528 20402 27580 20408
rect 27540 19786 27568 20402
rect 27528 19780 27580 19786
rect 27528 19722 27580 19728
rect 27068 15632 27120 15638
rect 27068 15574 27120 15580
rect 26240 15564 26292 15570
rect 26240 15506 26292 15512
rect 26056 15428 26108 15434
rect 26056 15370 26108 15376
rect 26068 15026 26096 15370
rect 26056 15020 26108 15026
rect 26056 14962 26108 14968
rect 26068 14346 26096 14962
rect 26056 14340 26108 14346
rect 26056 14282 26108 14288
rect 26068 13462 26096 14282
rect 26252 14006 26280 15506
rect 27724 15162 27752 23598
rect 29294 22876 29602 22885
rect 29294 22874 29300 22876
rect 29356 22874 29380 22876
rect 29436 22874 29460 22876
rect 29516 22874 29540 22876
rect 29596 22874 29602 22876
rect 29356 22822 29358 22874
rect 29538 22822 29540 22874
rect 29294 22820 29300 22822
rect 29356 22820 29380 22822
rect 29436 22820 29460 22822
rect 29516 22820 29540 22822
rect 29596 22820 29602 22822
rect 29294 22811 29602 22820
rect 29294 21788 29602 21797
rect 29294 21786 29300 21788
rect 29356 21786 29380 21788
rect 29436 21786 29460 21788
rect 29516 21786 29540 21788
rect 29596 21786 29602 21788
rect 29356 21734 29358 21786
rect 29538 21734 29540 21786
rect 29294 21732 29300 21734
rect 29356 21732 29380 21734
rect 29436 21732 29460 21734
rect 29516 21732 29540 21734
rect 29596 21732 29602 21734
rect 29294 21723 29602 21732
rect 29736 20936 29788 20942
rect 29736 20878 29788 20884
rect 30472 20936 30524 20942
rect 30472 20878 30524 20884
rect 29294 20700 29602 20709
rect 29294 20698 29300 20700
rect 29356 20698 29380 20700
rect 29436 20698 29460 20700
rect 29516 20698 29540 20700
rect 29596 20698 29602 20700
rect 29356 20646 29358 20698
rect 29538 20646 29540 20698
rect 29294 20644 29300 20646
rect 29356 20644 29380 20646
rect 29436 20644 29460 20646
rect 29516 20644 29540 20646
rect 29596 20644 29602 20646
rect 29294 20635 29602 20644
rect 29748 20602 29776 20878
rect 29920 20800 29972 20806
rect 29920 20742 29972 20748
rect 30380 20800 30432 20806
rect 30380 20742 30432 20748
rect 29736 20596 29788 20602
rect 29736 20538 29788 20544
rect 29932 19854 29960 20742
rect 28908 19848 28960 19854
rect 28908 19790 28960 19796
rect 29920 19848 29972 19854
rect 29920 19790 29972 19796
rect 28920 19514 28948 19790
rect 29294 19612 29602 19621
rect 29294 19610 29300 19612
rect 29356 19610 29380 19612
rect 29436 19610 29460 19612
rect 29516 19610 29540 19612
rect 29596 19610 29602 19612
rect 29356 19558 29358 19610
rect 29538 19558 29540 19610
rect 29294 19556 29300 19558
rect 29356 19556 29380 19558
rect 29436 19556 29460 19558
rect 29516 19556 29540 19558
rect 29596 19556 29602 19558
rect 29294 19547 29602 19556
rect 28908 19508 28960 19514
rect 28908 19450 28960 19456
rect 28920 19378 28948 19450
rect 30392 19378 30420 20742
rect 30484 20398 30512 20878
rect 30472 20392 30524 20398
rect 30472 20334 30524 20340
rect 30472 19712 30524 19718
rect 30472 19654 30524 19660
rect 30484 19514 30512 19654
rect 30472 19508 30524 19514
rect 30472 19450 30524 19456
rect 28908 19372 28960 19378
rect 28908 19314 28960 19320
rect 30380 19372 30432 19378
rect 30380 19314 30432 19320
rect 28920 17270 28948 19314
rect 30484 18970 30512 19450
rect 29828 18964 29880 18970
rect 29828 18906 29880 18912
rect 30472 18964 30524 18970
rect 30472 18906 30524 18912
rect 29294 18524 29602 18533
rect 29294 18522 29300 18524
rect 29356 18522 29380 18524
rect 29436 18522 29460 18524
rect 29516 18522 29540 18524
rect 29596 18522 29602 18524
rect 29356 18470 29358 18522
rect 29538 18470 29540 18522
rect 29294 18468 29300 18470
rect 29356 18468 29380 18470
rect 29436 18468 29460 18470
rect 29516 18468 29540 18470
rect 29596 18468 29602 18470
rect 29294 18459 29602 18468
rect 29092 17536 29144 17542
rect 29092 17478 29144 17484
rect 28908 17264 28960 17270
rect 28908 17206 28960 17212
rect 29104 17202 29132 17478
rect 29294 17436 29602 17445
rect 29294 17434 29300 17436
rect 29356 17434 29380 17436
rect 29436 17434 29460 17436
rect 29516 17434 29540 17436
rect 29596 17434 29602 17436
rect 29356 17382 29358 17434
rect 29538 17382 29540 17434
rect 29294 17380 29300 17382
rect 29356 17380 29380 17382
rect 29436 17380 29460 17382
rect 29516 17380 29540 17382
rect 29596 17380 29602 17382
rect 29294 17371 29602 17380
rect 29092 17196 29144 17202
rect 29092 17138 29144 17144
rect 29840 17066 29868 18906
rect 29828 17060 29880 17066
rect 29828 17002 29880 17008
rect 29294 16348 29602 16357
rect 29294 16346 29300 16348
rect 29356 16346 29380 16348
rect 29436 16346 29460 16348
rect 29516 16346 29540 16348
rect 29596 16346 29602 16348
rect 29356 16294 29358 16346
rect 29538 16294 29540 16346
rect 29294 16292 29300 16294
rect 29356 16292 29380 16294
rect 29436 16292 29460 16294
rect 29516 16292 29540 16294
rect 29596 16292 29602 16294
rect 29294 16283 29602 16292
rect 30196 15904 30248 15910
rect 30196 15846 30248 15852
rect 30012 15496 30064 15502
rect 30012 15438 30064 15444
rect 29294 15260 29602 15269
rect 29294 15258 29300 15260
rect 29356 15258 29380 15260
rect 29436 15258 29460 15260
rect 29516 15258 29540 15260
rect 29596 15258 29602 15260
rect 29356 15206 29358 15258
rect 29538 15206 29540 15258
rect 29294 15204 29300 15206
rect 29356 15204 29380 15206
rect 29436 15204 29460 15206
rect 29516 15204 29540 15206
rect 29596 15204 29602 15206
rect 29294 15195 29602 15204
rect 30024 15162 30052 15438
rect 27712 15156 27764 15162
rect 27712 15098 27764 15104
rect 30012 15156 30064 15162
rect 30012 15098 30064 15104
rect 26424 15088 26476 15094
rect 26424 15030 26476 15036
rect 26240 14000 26292 14006
rect 26240 13942 26292 13948
rect 26332 13864 26384 13870
rect 26332 13806 26384 13812
rect 26344 13530 26372 13806
rect 26332 13524 26384 13530
rect 26332 13466 26384 13472
rect 26056 13456 26108 13462
rect 26056 13398 26108 13404
rect 25136 13320 25188 13326
rect 25136 13262 25188 13268
rect 25044 13252 25096 13258
rect 25044 13194 25096 13200
rect 25056 12714 25084 13194
rect 26240 12980 26292 12986
rect 26240 12922 26292 12928
rect 25044 12708 25096 12714
rect 25044 12650 25096 12656
rect 24570 12540 24878 12549
rect 24570 12538 24576 12540
rect 24632 12538 24656 12540
rect 24712 12538 24736 12540
rect 24792 12538 24816 12540
rect 24872 12538 24878 12540
rect 24632 12486 24634 12538
rect 24814 12486 24816 12538
rect 24570 12484 24576 12486
rect 24632 12484 24656 12486
rect 24712 12484 24736 12486
rect 24792 12484 24816 12486
rect 24872 12484 24878 12486
rect 24570 12475 24878 12484
rect 25056 11830 25084 12650
rect 26252 12628 26280 12922
rect 26436 12646 26464 15030
rect 30208 15026 30236 15846
rect 30196 15020 30248 15026
rect 30196 14962 30248 14968
rect 26976 14952 27028 14958
rect 26976 14894 27028 14900
rect 26988 14414 27016 14894
rect 27252 14612 27304 14618
rect 27252 14554 27304 14560
rect 26976 14408 27028 14414
rect 26976 14350 27028 14356
rect 27264 13734 27292 14554
rect 29294 14172 29602 14181
rect 29294 14170 29300 14172
rect 29356 14170 29380 14172
rect 29436 14170 29460 14172
rect 29516 14170 29540 14172
rect 29596 14170 29602 14172
rect 29356 14118 29358 14170
rect 29538 14118 29540 14170
rect 29294 14116 29300 14118
rect 29356 14116 29380 14118
rect 29436 14116 29460 14118
rect 29516 14116 29540 14118
rect 29596 14116 29602 14118
rect 29294 14107 29602 14116
rect 30288 13864 30340 13870
rect 30288 13806 30340 13812
rect 27252 13728 27304 13734
rect 27252 13670 27304 13676
rect 27436 13728 27488 13734
rect 27436 13670 27488 13676
rect 27160 12980 27212 12986
rect 27264 12968 27292 13670
rect 27212 12940 27292 12968
rect 27160 12922 27212 12928
rect 26424 12640 26476 12646
rect 26252 12600 26424 12628
rect 26252 12238 26280 12600
rect 26424 12582 26476 12588
rect 27344 12640 27396 12646
rect 27344 12582 27396 12588
rect 27356 12238 27384 12582
rect 26240 12232 26292 12238
rect 26240 12174 26292 12180
rect 27344 12232 27396 12238
rect 27344 12174 27396 12180
rect 25228 12096 25280 12102
rect 25228 12038 25280 12044
rect 27252 12096 27304 12102
rect 27252 12038 27304 12044
rect 25044 11824 25096 11830
rect 25044 11766 25096 11772
rect 24570 11452 24878 11461
rect 24570 11450 24576 11452
rect 24632 11450 24656 11452
rect 24712 11450 24736 11452
rect 24792 11450 24816 11452
rect 24872 11450 24878 11452
rect 24632 11398 24634 11450
rect 24814 11398 24816 11450
rect 24570 11396 24576 11398
rect 24632 11396 24656 11398
rect 24712 11396 24736 11398
rect 24792 11396 24816 11398
rect 24872 11396 24878 11398
rect 24570 11387 24878 11396
rect 25240 11354 25268 12038
rect 27264 11762 27292 12038
rect 27252 11756 27304 11762
rect 27252 11698 27304 11704
rect 25228 11348 25280 11354
rect 25228 11290 25280 11296
rect 23572 11076 23624 11082
rect 23572 11018 23624 11024
rect 23756 11076 23808 11082
rect 23756 11018 23808 11024
rect 24492 11076 24544 11082
rect 24492 11018 24544 11024
rect 22928 10804 22980 10810
rect 22928 10746 22980 10752
rect 22468 10736 22520 10742
rect 22468 10678 22520 10684
rect 20812 9988 20864 9994
rect 20812 9930 20864 9936
rect 19846 9820 20154 9829
rect 19846 9818 19852 9820
rect 19908 9818 19932 9820
rect 19988 9818 20012 9820
rect 20068 9818 20092 9820
rect 20148 9818 20154 9820
rect 19908 9766 19910 9818
rect 20090 9766 20092 9818
rect 19846 9764 19852 9766
rect 19908 9764 19932 9766
rect 19988 9764 20012 9766
rect 20068 9764 20092 9766
rect 20148 9764 20154 9766
rect 19846 9755 20154 9764
rect 22480 9654 22508 10678
rect 22468 9648 22520 9654
rect 22468 9590 22520 9596
rect 22008 9580 22060 9586
rect 22008 9522 22060 9528
rect 20260 9512 20312 9518
rect 20260 9454 20312 9460
rect 19846 8732 20154 8741
rect 19846 8730 19852 8732
rect 19908 8730 19932 8732
rect 19988 8730 20012 8732
rect 20068 8730 20092 8732
rect 20148 8730 20154 8732
rect 19908 8678 19910 8730
rect 20090 8678 20092 8730
rect 19846 8676 19852 8678
rect 19908 8676 19932 8678
rect 19988 8676 20012 8678
rect 20068 8676 20092 8678
rect 20148 8676 20154 8678
rect 19846 8667 20154 8676
rect 20272 8430 20300 9454
rect 20628 9376 20680 9382
rect 20628 9318 20680 9324
rect 20640 8838 20668 9318
rect 22020 9178 22048 9522
rect 22480 9178 22508 9590
rect 22940 9586 22968 10746
rect 22928 9580 22980 9586
rect 22928 9522 22980 9528
rect 22008 9172 22060 9178
rect 22008 9114 22060 9120
rect 22468 9172 22520 9178
rect 22468 9114 22520 9120
rect 22480 9042 22508 9114
rect 21088 9036 21140 9042
rect 21088 8978 21140 8984
rect 22468 9036 22520 9042
rect 22468 8978 22520 8984
rect 20812 8968 20864 8974
rect 20812 8910 20864 8916
rect 20628 8832 20680 8838
rect 20628 8774 20680 8780
rect 20640 8566 20668 8774
rect 20824 8566 20852 8910
rect 21100 8566 21128 8978
rect 22284 8968 22336 8974
rect 22284 8910 22336 8916
rect 20628 8560 20680 8566
rect 20628 8502 20680 8508
rect 20812 8560 20864 8566
rect 20812 8502 20864 8508
rect 21088 8560 21140 8566
rect 21088 8502 21140 8508
rect 22296 8498 22324 8910
rect 23480 8560 23532 8566
rect 23480 8502 23532 8508
rect 22284 8492 22336 8498
rect 22284 8434 22336 8440
rect 22468 8492 22520 8498
rect 22468 8434 22520 8440
rect 20260 8424 20312 8430
rect 20260 8366 20312 8372
rect 19846 7644 20154 7653
rect 19846 7642 19852 7644
rect 19908 7642 19932 7644
rect 19988 7642 20012 7644
rect 20068 7642 20092 7644
rect 20148 7642 20154 7644
rect 19908 7590 19910 7642
rect 20090 7590 20092 7642
rect 19846 7588 19852 7590
rect 19908 7588 19932 7590
rect 19988 7588 20012 7590
rect 20068 7588 20092 7590
rect 20148 7588 20154 7590
rect 19846 7579 20154 7588
rect 19708 6928 19760 6934
rect 19708 6870 19760 6876
rect 19720 5846 19748 6870
rect 19846 6556 20154 6565
rect 19846 6554 19852 6556
rect 19908 6554 19932 6556
rect 19988 6554 20012 6556
rect 20068 6554 20092 6556
rect 20148 6554 20154 6556
rect 19908 6502 19910 6554
rect 20090 6502 20092 6554
rect 19846 6500 19852 6502
rect 19908 6500 19932 6502
rect 19988 6500 20012 6502
rect 20068 6500 20092 6502
rect 20148 6500 20154 6502
rect 19846 6491 20154 6500
rect 19708 5840 19760 5846
rect 19708 5782 19760 5788
rect 20272 5710 20300 8366
rect 22008 7336 22060 7342
rect 22008 7278 22060 7284
rect 20536 6180 20588 6186
rect 20536 6122 20588 6128
rect 20260 5704 20312 5710
rect 20260 5646 20312 5652
rect 19846 5468 20154 5477
rect 19846 5466 19852 5468
rect 19908 5466 19932 5468
rect 19988 5466 20012 5468
rect 20068 5466 20092 5468
rect 20148 5466 20154 5468
rect 19908 5414 19910 5466
rect 20090 5414 20092 5466
rect 19846 5412 19852 5414
rect 19908 5412 19932 5414
rect 19988 5412 20012 5414
rect 20068 5412 20092 5414
rect 20148 5412 20154 5414
rect 19846 5403 20154 5412
rect 20272 5302 20300 5646
rect 20260 5296 20312 5302
rect 20260 5238 20312 5244
rect 20548 5234 20576 6122
rect 22020 5778 22048 7278
rect 22008 5772 22060 5778
rect 22008 5714 22060 5720
rect 22376 5704 22428 5710
rect 22376 5646 22428 5652
rect 22388 5234 22416 5646
rect 22480 5370 22508 8434
rect 23020 8356 23072 8362
rect 23020 8298 23072 8304
rect 23032 7478 23060 8298
rect 23492 8090 23520 8502
rect 23480 8084 23532 8090
rect 23480 8026 23532 8032
rect 23020 7472 23072 7478
rect 23020 7414 23072 7420
rect 23204 5840 23256 5846
rect 23204 5782 23256 5788
rect 22468 5364 22520 5370
rect 22468 5306 22520 5312
rect 20076 5228 20128 5234
rect 20076 5170 20128 5176
rect 20536 5228 20588 5234
rect 20536 5170 20588 5176
rect 22376 5228 22428 5234
rect 22376 5170 22428 5176
rect 22560 5228 22612 5234
rect 22560 5170 22612 5176
rect 20088 4554 20116 5170
rect 20260 5160 20312 5166
rect 20260 5102 20312 5108
rect 20168 5024 20220 5030
rect 20168 4966 20220 4972
rect 20180 4622 20208 4966
rect 20272 4826 20300 5102
rect 20260 4820 20312 4826
rect 20260 4762 20312 4768
rect 20168 4616 20220 4622
rect 20168 4558 20220 4564
rect 20076 4548 20128 4554
rect 20076 4490 20128 4496
rect 19628 4406 19748 4434
rect 18328 4140 18380 4146
rect 18328 4082 18380 4088
rect 19720 3942 19748 4406
rect 19846 4380 20154 4389
rect 19846 4378 19852 4380
rect 19908 4378 19932 4380
rect 19988 4378 20012 4380
rect 20068 4378 20092 4380
rect 20148 4378 20154 4380
rect 19908 4326 19910 4378
rect 20090 4326 20092 4378
rect 19846 4324 19852 4326
rect 19908 4324 19932 4326
rect 19988 4324 20012 4326
rect 20068 4324 20092 4326
rect 20148 4324 20154 4326
rect 19846 4315 20154 4324
rect 20272 4146 20300 4762
rect 20548 4622 20576 5170
rect 20536 4616 20588 4622
rect 20536 4558 20588 4564
rect 22388 4554 22416 5170
rect 22572 4826 22600 5170
rect 22560 4820 22612 4826
rect 22560 4762 22612 4768
rect 23216 4690 23244 5782
rect 23204 4684 23256 4690
rect 23204 4626 23256 4632
rect 20444 4548 20496 4554
rect 20444 4490 20496 4496
rect 22376 4548 22428 4554
rect 22376 4490 22428 4496
rect 20456 4146 20484 4490
rect 23480 4480 23532 4486
rect 23480 4422 23532 4428
rect 23492 4146 23520 4422
rect 20260 4140 20312 4146
rect 20260 4082 20312 4088
rect 20444 4140 20496 4146
rect 20444 4082 20496 4088
rect 23480 4140 23532 4146
rect 23480 4082 23532 4088
rect 19708 3936 19760 3942
rect 19708 3878 19760 3884
rect 20260 3936 20312 3942
rect 20260 3878 20312 3884
rect 19248 3528 19300 3534
rect 19248 3470 19300 3476
rect 17592 2984 17644 2990
rect 17592 2926 17644 2932
rect 17592 2848 17644 2854
rect 17592 2790 17644 2796
rect 16856 2644 16908 2650
rect 16856 2586 16908 2592
rect 14832 2576 14884 2582
rect 14832 2518 14884 2524
rect 16764 2576 16816 2582
rect 16764 2518 16816 2524
rect 17604 2446 17632 2790
rect 19260 2650 19288 3470
rect 19248 2644 19300 2650
rect 19248 2586 19300 2592
rect 2228 2440 2280 2446
rect 2228 2382 2280 2388
rect 5540 2440 5592 2446
rect 5540 2382 5592 2388
rect 6276 2440 6328 2446
rect 6276 2382 6328 2388
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 8392 2440 8444 2446
rect 8392 2382 8444 2388
rect 12440 2440 12492 2446
rect 12440 2382 12492 2388
rect 12808 2440 12860 2446
rect 12808 2382 12860 2388
rect 14004 2440 14056 2446
rect 14004 2382 14056 2388
rect 15200 2440 15252 2446
rect 15200 2382 15252 2388
rect 16396 2440 16448 2446
rect 16396 2382 16448 2388
rect 17592 2440 17644 2446
rect 17592 2382 17644 2388
rect 18788 2440 18840 2446
rect 18788 2382 18840 2388
rect 1492 2304 1544 2310
rect 1492 2246 1544 2252
rect 2044 2304 2096 2310
rect 2044 2246 2096 2252
rect 3240 2304 3292 2310
rect 3240 2246 3292 2252
rect 4436 2304 4488 2310
rect 4436 2246 4488 2252
rect 5632 2304 5684 2310
rect 5632 2246 5684 2252
rect 6828 2304 6880 2310
rect 6828 2246 6880 2252
rect 8024 2304 8076 2310
rect 8024 2246 8076 2252
rect 9220 2304 9272 2310
rect 9220 2246 9272 2252
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 1504 1737 1532 2246
rect 1490 1728 1546 1737
rect 1490 1663 1546 1672
rect 2056 800 2084 2246
rect 3252 800 3280 2246
rect 4448 800 4476 2246
rect 5644 800 5672 2246
rect 6840 800 6868 2246
rect 8036 800 8064 2246
rect 9232 800 9260 2246
rect 10398 2204 10706 2213
rect 10398 2202 10404 2204
rect 10460 2202 10484 2204
rect 10540 2202 10564 2204
rect 10620 2202 10644 2204
rect 10700 2202 10706 2204
rect 10460 2150 10462 2202
rect 10642 2150 10644 2202
rect 10398 2148 10404 2150
rect 10460 2148 10484 2150
rect 10540 2148 10564 2150
rect 10620 2148 10644 2150
rect 10700 2148 10706 2150
rect 10398 2139 10706 2148
rect 11624 800 11652 2246
rect 12820 800 12848 2382
rect 14016 800 14044 2382
rect 15212 800 15240 2382
rect 16408 800 16436 2382
rect 17604 800 17632 2382
rect 18800 2310 18828 2382
rect 19720 2378 19748 3878
rect 20272 3602 20300 3878
rect 20720 3732 20772 3738
rect 20720 3674 20772 3680
rect 20260 3596 20312 3602
rect 20260 3538 20312 3544
rect 19846 3292 20154 3301
rect 19846 3290 19852 3292
rect 19908 3290 19932 3292
rect 19988 3290 20012 3292
rect 20068 3290 20092 3292
rect 20148 3290 20154 3292
rect 19908 3238 19910 3290
rect 20090 3238 20092 3290
rect 19846 3236 19852 3238
rect 19908 3236 19932 3238
rect 19988 3236 20012 3238
rect 20068 3236 20092 3238
rect 20148 3236 20154 3238
rect 19846 3227 20154 3236
rect 20260 2848 20312 2854
rect 20260 2790 20312 2796
rect 20272 2446 20300 2790
rect 20732 2650 20760 3674
rect 22928 3596 22980 3602
rect 22928 3538 22980 3544
rect 21364 3528 21416 3534
rect 21364 3470 21416 3476
rect 21376 2650 21404 3470
rect 22468 3460 22520 3466
rect 22468 3402 22520 3408
rect 22480 2650 22508 3402
rect 22940 2650 22968 3538
rect 23480 3392 23532 3398
rect 23480 3334 23532 3340
rect 20720 2644 20772 2650
rect 20720 2586 20772 2592
rect 21364 2644 21416 2650
rect 21364 2586 21416 2592
rect 22468 2644 22520 2650
rect 22468 2586 22520 2592
rect 22928 2644 22980 2650
rect 22928 2586 22980 2592
rect 20260 2440 20312 2446
rect 20260 2382 20312 2388
rect 22376 2440 22428 2446
rect 23492 2428 23520 3334
rect 23584 3058 23612 11018
rect 23768 8294 23796 11018
rect 24570 10364 24878 10373
rect 24570 10362 24576 10364
rect 24632 10362 24656 10364
rect 24712 10362 24736 10364
rect 24792 10362 24816 10364
rect 24872 10362 24878 10364
rect 24632 10310 24634 10362
rect 24814 10310 24816 10362
rect 24570 10308 24576 10310
rect 24632 10308 24656 10310
rect 24712 10308 24736 10310
rect 24792 10308 24816 10310
rect 24872 10308 24878 10310
rect 24570 10299 24878 10308
rect 27448 10062 27476 13670
rect 29294 13084 29602 13093
rect 29294 13082 29300 13084
rect 29356 13082 29380 13084
rect 29436 13082 29460 13084
rect 29516 13082 29540 13084
rect 29596 13082 29602 13084
rect 29356 13030 29358 13082
rect 29538 13030 29540 13082
rect 29294 13028 29300 13030
rect 29356 13028 29380 13030
rect 29436 13028 29460 13030
rect 29516 13028 29540 13030
rect 29596 13028 29602 13030
rect 29294 13019 29602 13028
rect 30300 12850 30328 13806
rect 30576 12986 30604 24006
rect 30668 17338 30696 25774
rect 31220 24750 31248 27950
rect 31404 27606 31432 29242
rect 32312 29164 32364 29170
rect 32312 29106 32364 29112
rect 31576 28484 31628 28490
rect 31576 28426 31628 28432
rect 31392 27600 31444 27606
rect 31392 27542 31444 27548
rect 31300 26988 31352 26994
rect 31404 26976 31432 27542
rect 31352 26948 31432 26976
rect 31300 26930 31352 26936
rect 31208 24744 31260 24750
rect 31208 24686 31260 24692
rect 31220 24070 31248 24686
rect 31300 24268 31352 24274
rect 31300 24210 31352 24216
rect 31208 24064 31260 24070
rect 31208 24006 31260 24012
rect 30932 23112 30984 23118
rect 30932 23054 30984 23060
rect 30944 21554 30972 23054
rect 30932 21548 30984 21554
rect 30932 21490 30984 21496
rect 31220 20330 31248 24006
rect 31312 23730 31340 24210
rect 31300 23724 31352 23730
rect 31300 23666 31352 23672
rect 31312 23526 31340 23666
rect 31300 23520 31352 23526
rect 31300 23462 31352 23468
rect 31312 20466 31340 23462
rect 31588 22094 31616 28426
rect 32324 28422 32352 29106
rect 34018 28860 34326 28869
rect 34018 28858 34024 28860
rect 34080 28858 34104 28860
rect 34160 28858 34184 28860
rect 34240 28858 34264 28860
rect 34320 28858 34326 28860
rect 34080 28806 34082 28858
rect 34262 28806 34264 28858
rect 34018 28804 34024 28806
rect 34080 28804 34104 28806
rect 34160 28804 34184 28806
rect 34240 28804 34264 28806
rect 34320 28804 34326 28806
rect 34018 28795 34326 28804
rect 34808 28762 34836 29242
rect 34796 28756 34848 28762
rect 34796 28698 34848 28704
rect 32312 28416 32364 28422
rect 32312 28358 32364 28364
rect 32324 28150 32352 28358
rect 32312 28144 32364 28150
rect 32312 28086 32364 28092
rect 31852 28076 31904 28082
rect 31852 28018 31904 28024
rect 31864 26994 31892 28018
rect 31852 26988 31904 26994
rect 31852 26930 31904 26936
rect 31668 26784 31720 26790
rect 31668 26726 31720 26732
rect 31680 26382 31708 26726
rect 31668 26376 31720 26382
rect 31668 26318 31720 26324
rect 31864 23730 31892 26930
rect 32324 26234 32352 28086
rect 34808 28014 34836 28698
rect 34520 28008 34572 28014
rect 34520 27950 34572 27956
rect 34796 28008 34848 28014
rect 34796 27950 34848 27956
rect 34018 27772 34326 27781
rect 34018 27770 34024 27772
rect 34080 27770 34104 27772
rect 34160 27770 34184 27772
rect 34240 27770 34264 27772
rect 34320 27770 34326 27772
rect 34080 27718 34082 27770
rect 34262 27718 34264 27770
rect 34018 27716 34024 27718
rect 34080 27716 34104 27718
rect 34160 27716 34184 27718
rect 34240 27716 34264 27718
rect 34320 27716 34326 27718
rect 34018 27707 34326 27716
rect 32956 26988 33008 26994
rect 32956 26930 33008 26936
rect 32968 26586 32996 26930
rect 33784 26920 33836 26926
rect 33784 26862 33836 26868
rect 32956 26580 33008 26586
rect 32956 26522 33008 26528
rect 32232 26206 32352 26234
rect 31852 23724 31904 23730
rect 31852 23666 31904 23672
rect 31864 23186 31892 23666
rect 32036 23656 32088 23662
rect 32036 23598 32088 23604
rect 31852 23180 31904 23186
rect 31852 23122 31904 23128
rect 31588 22066 31708 22094
rect 31300 20460 31352 20466
rect 31300 20402 31352 20408
rect 31208 20324 31260 20330
rect 31208 20266 31260 20272
rect 30656 17332 30708 17338
rect 30656 17274 30708 17280
rect 30748 17060 30800 17066
rect 30748 17002 30800 17008
rect 30760 15706 30788 17002
rect 30748 15700 30800 15706
rect 30748 15642 30800 15648
rect 31484 15020 31536 15026
rect 31484 14962 31536 14968
rect 31496 14618 31524 14962
rect 31300 14612 31352 14618
rect 31300 14554 31352 14560
rect 31484 14612 31536 14618
rect 31484 14554 31536 14560
rect 30656 14476 30708 14482
rect 30656 14418 30708 14424
rect 30564 12980 30616 12986
rect 30564 12922 30616 12928
rect 30288 12844 30340 12850
rect 30288 12786 30340 12792
rect 29294 11996 29602 12005
rect 29294 11994 29300 11996
rect 29356 11994 29380 11996
rect 29436 11994 29460 11996
rect 29516 11994 29540 11996
rect 29596 11994 29602 11996
rect 29356 11942 29358 11994
rect 29538 11942 29540 11994
rect 29294 11940 29300 11942
rect 29356 11940 29380 11942
rect 29436 11940 29460 11942
rect 29516 11940 29540 11942
rect 29596 11940 29602 11942
rect 29294 11931 29602 11940
rect 28724 11756 28776 11762
rect 28724 11698 28776 11704
rect 28736 11354 28764 11698
rect 28724 11348 28776 11354
rect 28724 11290 28776 11296
rect 29294 10908 29602 10917
rect 29294 10906 29300 10908
rect 29356 10906 29380 10908
rect 29436 10906 29460 10908
rect 29516 10906 29540 10908
rect 29596 10906 29602 10908
rect 29356 10854 29358 10906
rect 29538 10854 29540 10906
rect 29294 10852 29300 10854
rect 29356 10852 29380 10854
rect 29436 10852 29460 10854
rect 29516 10852 29540 10854
rect 29596 10852 29602 10854
rect 29294 10843 29602 10852
rect 27436 10056 27488 10062
rect 27436 9998 27488 10004
rect 27436 9920 27488 9926
rect 27436 9862 27488 9868
rect 24400 9580 24452 9586
rect 24400 9522 24452 9528
rect 24412 9178 24440 9522
rect 26792 9512 26844 9518
rect 26792 9454 26844 9460
rect 24570 9276 24878 9285
rect 24570 9274 24576 9276
rect 24632 9274 24656 9276
rect 24712 9274 24736 9276
rect 24792 9274 24816 9276
rect 24872 9274 24878 9276
rect 24632 9222 24634 9274
rect 24814 9222 24816 9274
rect 24570 9220 24576 9222
rect 24632 9220 24656 9222
rect 24712 9220 24736 9222
rect 24792 9220 24816 9222
rect 24872 9220 24878 9222
rect 24570 9211 24878 9220
rect 26804 9178 26832 9454
rect 27160 9376 27212 9382
rect 27160 9318 27212 9324
rect 24400 9172 24452 9178
rect 24400 9114 24452 9120
rect 26792 9172 26844 9178
rect 26792 9114 26844 9120
rect 27172 8974 27200 9318
rect 27448 9042 27476 9862
rect 29294 9820 29602 9829
rect 29294 9818 29300 9820
rect 29356 9818 29380 9820
rect 29436 9818 29460 9820
rect 29516 9818 29540 9820
rect 29596 9818 29602 9820
rect 29356 9766 29358 9818
rect 29538 9766 29540 9818
rect 29294 9764 29300 9766
rect 29356 9764 29380 9766
rect 29436 9764 29460 9766
rect 29516 9764 29540 9766
rect 29596 9764 29602 9766
rect 29294 9755 29602 9764
rect 30668 9518 30696 14418
rect 31116 12980 31168 12986
rect 31116 12922 31168 12928
rect 30656 9512 30708 9518
rect 30656 9454 30708 9460
rect 30380 9444 30432 9450
rect 30380 9386 30432 9392
rect 27436 9036 27488 9042
rect 27436 8978 27488 8984
rect 24768 8968 24820 8974
rect 24768 8910 24820 8916
rect 27160 8968 27212 8974
rect 27160 8910 27212 8916
rect 24780 8498 24808 8910
rect 24860 8900 24912 8906
rect 24860 8842 24912 8848
rect 24768 8492 24820 8498
rect 24768 8434 24820 8440
rect 24872 8430 24900 8842
rect 27448 8430 27476 8978
rect 28724 8832 28776 8838
rect 28724 8774 28776 8780
rect 28736 8430 28764 8774
rect 29294 8732 29602 8741
rect 29294 8730 29300 8732
rect 29356 8730 29380 8732
rect 29436 8730 29460 8732
rect 29516 8730 29540 8732
rect 29596 8730 29602 8732
rect 29356 8678 29358 8730
rect 29538 8678 29540 8730
rect 29294 8676 29300 8678
rect 29356 8676 29380 8678
rect 29436 8676 29460 8678
rect 29516 8676 29540 8678
rect 29596 8676 29602 8678
rect 29294 8667 29602 8676
rect 30288 8628 30340 8634
rect 30288 8570 30340 8576
rect 24860 8424 24912 8430
rect 24860 8366 24912 8372
rect 27436 8424 27488 8430
rect 27436 8366 27488 8372
rect 27620 8424 27672 8430
rect 27620 8366 27672 8372
rect 28724 8424 28776 8430
rect 28724 8366 28776 8372
rect 23756 8288 23808 8294
rect 23756 8230 23808 8236
rect 23768 4214 23796 8230
rect 24570 8188 24878 8197
rect 24570 8186 24576 8188
rect 24632 8186 24656 8188
rect 24712 8186 24736 8188
rect 24792 8186 24816 8188
rect 24872 8186 24878 8188
rect 24632 8134 24634 8186
rect 24814 8134 24816 8186
rect 24570 8132 24576 8134
rect 24632 8132 24656 8134
rect 24712 8132 24736 8134
rect 24792 8132 24816 8134
rect 24872 8132 24878 8134
rect 24570 8123 24878 8132
rect 27632 7886 27660 8366
rect 30300 8362 30328 8570
rect 30392 8566 30420 9386
rect 30472 9376 30524 9382
rect 30472 9318 30524 9324
rect 30484 8906 30512 9318
rect 30668 8974 30696 9454
rect 30656 8968 30708 8974
rect 30656 8910 30708 8916
rect 30472 8900 30524 8906
rect 30472 8842 30524 8848
rect 30484 8634 30512 8842
rect 30748 8832 30800 8838
rect 30748 8774 30800 8780
rect 30472 8628 30524 8634
rect 30472 8570 30524 8576
rect 30380 8560 30432 8566
rect 30380 8502 30432 8508
rect 30288 8356 30340 8362
rect 30288 8298 30340 8304
rect 27620 7880 27672 7886
rect 27620 7822 27672 7828
rect 30104 7744 30156 7750
rect 30104 7686 30156 7692
rect 29294 7644 29602 7653
rect 29294 7642 29300 7644
rect 29356 7642 29380 7644
rect 29436 7642 29460 7644
rect 29516 7642 29540 7644
rect 29596 7642 29602 7644
rect 29356 7590 29358 7642
rect 29538 7590 29540 7642
rect 29294 7588 29300 7590
rect 29356 7588 29380 7590
rect 29436 7588 29460 7590
rect 29516 7588 29540 7590
rect 29596 7588 29602 7590
rect 29294 7579 29602 7588
rect 30116 7206 30144 7686
rect 30392 7478 30420 8502
rect 30484 8294 30512 8570
rect 30760 8498 30788 8774
rect 30748 8492 30800 8498
rect 30748 8434 30800 8440
rect 30472 8288 30524 8294
rect 30472 8230 30524 8236
rect 30760 7546 30788 8434
rect 31128 8090 31156 12922
rect 31312 12918 31340 14554
rect 31680 12918 31708 22066
rect 32048 16574 32076 23598
rect 31956 16546 32076 16574
rect 32128 16584 32180 16590
rect 31956 13002 31984 16546
rect 32128 16526 32180 16532
rect 32140 16402 32168 16526
rect 32048 16374 32168 16402
rect 32048 14278 32076 16374
rect 32036 14272 32088 14278
rect 32036 14214 32088 14220
rect 32048 13938 32076 14214
rect 32036 13932 32088 13938
rect 32036 13874 32088 13880
rect 31956 12974 32076 13002
rect 31300 12912 31352 12918
rect 31300 12854 31352 12860
rect 31668 12912 31720 12918
rect 31668 12854 31720 12860
rect 31944 12912 31996 12918
rect 31944 12854 31996 12860
rect 31760 12640 31812 12646
rect 31760 12582 31812 12588
rect 31772 12170 31800 12582
rect 31956 12442 31984 12854
rect 31944 12436 31996 12442
rect 31944 12378 31996 12384
rect 31760 12164 31812 12170
rect 31760 12106 31812 12112
rect 31772 11354 31800 12106
rect 31760 11348 31812 11354
rect 31760 11290 31812 11296
rect 31484 11212 31536 11218
rect 31484 11154 31536 11160
rect 31496 11082 31524 11154
rect 31484 11076 31536 11082
rect 31484 11018 31536 11024
rect 31116 8084 31168 8090
rect 31116 8026 31168 8032
rect 30748 7540 30800 7546
rect 30748 7482 30800 7488
rect 30380 7472 30432 7478
rect 30380 7414 30432 7420
rect 30104 7200 30156 7206
rect 30104 7142 30156 7148
rect 24570 7100 24878 7109
rect 24570 7098 24576 7100
rect 24632 7098 24656 7100
rect 24712 7098 24736 7100
rect 24792 7098 24816 7100
rect 24872 7098 24878 7100
rect 24632 7046 24634 7098
rect 24814 7046 24816 7098
rect 24570 7044 24576 7046
rect 24632 7044 24656 7046
rect 24712 7044 24736 7046
rect 24792 7044 24816 7046
rect 24872 7044 24878 7046
rect 24570 7035 24878 7044
rect 26516 6792 26568 6798
rect 26516 6734 26568 6740
rect 26884 6792 26936 6798
rect 26884 6734 26936 6740
rect 24570 6012 24878 6021
rect 24570 6010 24576 6012
rect 24632 6010 24656 6012
rect 24712 6010 24736 6012
rect 24792 6010 24816 6012
rect 24872 6010 24878 6012
rect 24632 5958 24634 6010
rect 24814 5958 24816 6010
rect 24570 5956 24576 5958
rect 24632 5956 24656 5958
rect 24712 5956 24736 5958
rect 24792 5956 24816 5958
rect 24872 5956 24878 5958
rect 24570 5947 24878 5956
rect 26528 5370 26556 6734
rect 26896 5710 26924 6734
rect 29294 6556 29602 6565
rect 29294 6554 29300 6556
rect 29356 6554 29380 6556
rect 29436 6554 29460 6556
rect 29516 6554 29540 6556
rect 29596 6554 29602 6556
rect 29356 6502 29358 6554
rect 29538 6502 29540 6554
rect 29294 6500 29300 6502
rect 29356 6500 29380 6502
rect 29436 6500 29460 6502
rect 29516 6500 29540 6502
rect 29596 6500 29602 6502
rect 29294 6491 29602 6500
rect 30116 5914 30144 7142
rect 30392 7002 30420 7414
rect 30380 6996 30432 7002
rect 30380 6938 30432 6944
rect 30760 6662 30788 7482
rect 31496 7002 31524 11018
rect 31852 11008 31904 11014
rect 31852 10950 31904 10956
rect 31864 10674 31892 10950
rect 31852 10668 31904 10674
rect 31852 10610 31904 10616
rect 31956 9178 31984 12378
rect 32048 11082 32076 12974
rect 32232 11218 32260 26206
rect 32956 24812 33008 24818
rect 32956 24754 33008 24760
rect 32864 24744 32916 24750
rect 32864 24686 32916 24692
rect 32876 24206 32904 24686
rect 32864 24200 32916 24206
rect 32864 24142 32916 24148
rect 32968 23866 32996 24754
rect 33796 24614 33824 26862
rect 33876 26784 33928 26790
rect 33876 26726 33928 26732
rect 33140 24608 33192 24614
rect 33140 24550 33192 24556
rect 33784 24608 33836 24614
rect 33784 24550 33836 24556
rect 33152 24206 33180 24550
rect 33140 24200 33192 24206
rect 33140 24142 33192 24148
rect 32956 23860 33008 23866
rect 32956 23802 33008 23808
rect 33796 23798 33824 24550
rect 33888 24206 33916 26726
rect 34018 26684 34326 26693
rect 34018 26682 34024 26684
rect 34080 26682 34104 26684
rect 34160 26682 34184 26684
rect 34240 26682 34264 26684
rect 34320 26682 34326 26684
rect 34080 26630 34082 26682
rect 34262 26630 34264 26682
rect 34018 26628 34024 26630
rect 34080 26628 34104 26630
rect 34160 26628 34184 26630
rect 34240 26628 34264 26630
rect 34320 26628 34326 26630
rect 34018 26619 34326 26628
rect 34018 25596 34326 25605
rect 34018 25594 34024 25596
rect 34080 25594 34104 25596
rect 34160 25594 34184 25596
rect 34240 25594 34264 25596
rect 34320 25594 34326 25596
rect 34080 25542 34082 25594
rect 34262 25542 34264 25594
rect 34018 25540 34024 25542
rect 34080 25540 34104 25542
rect 34160 25540 34184 25542
rect 34240 25540 34264 25542
rect 34320 25540 34326 25542
rect 34018 25531 34326 25540
rect 34018 24508 34326 24517
rect 34018 24506 34024 24508
rect 34080 24506 34104 24508
rect 34160 24506 34184 24508
rect 34240 24506 34264 24508
rect 34320 24506 34326 24508
rect 34080 24454 34082 24506
rect 34262 24454 34264 24506
rect 34018 24452 34024 24454
rect 34080 24452 34104 24454
rect 34160 24452 34184 24454
rect 34240 24452 34264 24454
rect 34320 24452 34326 24454
rect 34018 24443 34326 24452
rect 33876 24200 33928 24206
rect 33876 24142 33928 24148
rect 33888 23866 33916 24142
rect 33876 23860 33928 23866
rect 33876 23802 33928 23808
rect 33784 23792 33836 23798
rect 33784 23734 33836 23740
rect 33888 22030 33916 23802
rect 34018 23420 34326 23429
rect 34018 23418 34024 23420
rect 34080 23418 34104 23420
rect 34160 23418 34184 23420
rect 34240 23418 34264 23420
rect 34320 23418 34326 23420
rect 34080 23366 34082 23418
rect 34262 23366 34264 23418
rect 34018 23364 34024 23366
rect 34080 23364 34104 23366
rect 34160 23364 34184 23366
rect 34240 23364 34264 23366
rect 34320 23364 34326 23366
rect 34018 23355 34326 23364
rect 34018 22332 34326 22341
rect 34018 22330 34024 22332
rect 34080 22330 34104 22332
rect 34160 22330 34184 22332
rect 34240 22330 34264 22332
rect 34320 22330 34326 22332
rect 34080 22278 34082 22330
rect 34262 22278 34264 22330
rect 34018 22276 34024 22278
rect 34080 22276 34104 22278
rect 34160 22276 34184 22278
rect 34240 22276 34264 22278
rect 34320 22276 34326 22278
rect 34018 22267 34326 22276
rect 33876 22024 33928 22030
rect 33876 21966 33928 21972
rect 34532 21554 34560 27950
rect 34980 27872 35032 27878
rect 34980 27814 35032 27820
rect 35900 27872 35952 27878
rect 35900 27814 35952 27820
rect 34992 27470 35020 27814
rect 34980 27464 35032 27470
rect 34980 27406 35032 27412
rect 35624 27464 35676 27470
rect 35624 27406 35676 27412
rect 35636 26926 35664 27406
rect 35912 26994 35940 27814
rect 36728 27464 36780 27470
rect 36728 27406 36780 27412
rect 36740 26994 36768 27406
rect 35900 26988 35952 26994
rect 35900 26930 35952 26936
rect 36728 26988 36780 26994
rect 36728 26930 36780 26936
rect 35624 26920 35676 26926
rect 35624 26862 35676 26868
rect 36740 23866 36768 26930
rect 36728 23860 36780 23866
rect 36728 23802 36780 23808
rect 36740 23730 36768 23802
rect 35900 23724 35952 23730
rect 35900 23666 35952 23672
rect 36728 23724 36780 23730
rect 36728 23666 36780 23672
rect 34612 23656 34664 23662
rect 34612 23598 34664 23604
rect 34520 21548 34572 21554
rect 34520 21490 34572 21496
rect 34428 21480 34480 21486
rect 34428 21422 34480 21428
rect 34018 21244 34326 21253
rect 34018 21242 34024 21244
rect 34080 21242 34104 21244
rect 34160 21242 34184 21244
rect 34240 21242 34264 21244
rect 34320 21242 34326 21244
rect 34080 21190 34082 21242
rect 34262 21190 34264 21242
rect 34018 21188 34024 21190
rect 34080 21188 34104 21190
rect 34160 21188 34184 21190
rect 34240 21188 34264 21190
rect 34320 21188 34326 21190
rect 34018 21179 34326 21188
rect 34440 20482 34468 21422
rect 34348 20466 34468 20482
rect 33232 20460 33284 20466
rect 33232 20402 33284 20408
rect 34336 20460 34468 20466
rect 34388 20454 34468 20460
rect 34336 20402 34388 20408
rect 33244 17202 33272 20402
rect 33876 20256 33928 20262
rect 33876 20198 33928 20204
rect 33888 19854 33916 20198
rect 34018 20156 34326 20165
rect 34018 20154 34024 20156
rect 34080 20154 34104 20156
rect 34160 20154 34184 20156
rect 34240 20154 34264 20156
rect 34320 20154 34326 20156
rect 34080 20102 34082 20154
rect 34262 20102 34264 20154
rect 34018 20100 34024 20102
rect 34080 20100 34104 20102
rect 34160 20100 34184 20102
rect 34240 20100 34264 20102
rect 34320 20100 34326 20102
rect 34018 20091 34326 20100
rect 33876 19848 33928 19854
rect 33876 19790 33928 19796
rect 34018 19068 34326 19077
rect 34018 19066 34024 19068
rect 34080 19066 34104 19068
rect 34160 19066 34184 19068
rect 34240 19066 34264 19068
rect 34320 19066 34326 19068
rect 34080 19014 34082 19066
rect 34262 19014 34264 19066
rect 34018 19012 34024 19014
rect 34080 19012 34104 19014
rect 34160 19012 34184 19014
rect 34240 19012 34264 19014
rect 34320 19012 34326 19014
rect 34018 19003 34326 19012
rect 34018 17980 34326 17989
rect 34018 17978 34024 17980
rect 34080 17978 34104 17980
rect 34160 17978 34184 17980
rect 34240 17978 34264 17980
rect 34320 17978 34326 17980
rect 34080 17926 34082 17978
rect 34262 17926 34264 17978
rect 34018 17924 34024 17926
rect 34080 17924 34104 17926
rect 34160 17924 34184 17926
rect 34240 17924 34264 17926
rect 34320 17924 34326 17926
rect 34018 17915 34326 17924
rect 33232 17196 33284 17202
rect 33232 17138 33284 17144
rect 33244 16658 33272 17138
rect 33416 16992 33468 16998
rect 33416 16934 33468 16940
rect 33232 16652 33284 16658
rect 33232 16594 33284 16600
rect 33244 16454 33272 16594
rect 33428 16590 33456 16934
rect 34018 16892 34326 16901
rect 34018 16890 34024 16892
rect 34080 16890 34104 16892
rect 34160 16890 34184 16892
rect 34240 16890 34264 16892
rect 34320 16890 34326 16892
rect 34080 16838 34082 16890
rect 34262 16838 34264 16890
rect 34018 16836 34024 16838
rect 34080 16836 34104 16838
rect 34160 16836 34184 16838
rect 34240 16836 34264 16838
rect 34320 16836 34326 16838
rect 34018 16827 34326 16836
rect 34624 16590 34652 23598
rect 35532 23520 35584 23526
rect 35532 23462 35584 23468
rect 35544 23118 35572 23462
rect 35912 23322 35940 23666
rect 35900 23316 35952 23322
rect 35900 23258 35952 23264
rect 35532 23112 35584 23118
rect 35532 23054 35584 23060
rect 35992 21344 36044 21350
rect 35992 21286 36044 21292
rect 36004 20942 36032 21286
rect 35992 20936 36044 20942
rect 35992 20878 36044 20884
rect 36912 20800 36964 20806
rect 36912 20742 36964 20748
rect 35992 20256 36044 20262
rect 35992 20198 36044 20204
rect 36004 19854 36032 20198
rect 35992 19848 36044 19854
rect 35992 19790 36044 19796
rect 35900 19780 35952 19786
rect 35900 19722 35952 19728
rect 34704 19712 34756 19718
rect 34704 19654 34756 19660
rect 34716 19378 34744 19654
rect 35912 19378 35940 19722
rect 34704 19372 34756 19378
rect 34704 19314 34756 19320
rect 35900 19372 35952 19378
rect 35900 19314 35952 19320
rect 36636 19372 36688 19378
rect 36636 19314 36688 19320
rect 36648 18766 36676 19314
rect 36924 18766 36952 20742
rect 37464 19712 37516 19718
rect 37464 19654 37516 19660
rect 37476 19514 37504 19654
rect 37464 19508 37516 19514
rect 37464 19450 37516 19456
rect 36636 18760 36688 18766
rect 36636 18702 36688 18708
rect 36912 18760 36964 18766
rect 36912 18702 36964 18708
rect 35072 17196 35124 17202
rect 35072 17138 35124 17144
rect 35084 16794 35112 17138
rect 35072 16788 35124 16794
rect 35072 16730 35124 16736
rect 33416 16584 33468 16590
rect 33416 16526 33468 16532
rect 34612 16584 34664 16590
rect 34612 16526 34664 16532
rect 35716 16584 35768 16590
rect 35716 16526 35768 16532
rect 33232 16448 33284 16454
rect 33232 16390 33284 16396
rect 34520 16108 34572 16114
rect 34520 16050 34572 16056
rect 34018 15804 34326 15813
rect 34018 15802 34024 15804
rect 34080 15802 34104 15804
rect 34160 15802 34184 15804
rect 34240 15802 34264 15804
rect 34320 15802 34326 15804
rect 34080 15750 34082 15802
rect 34262 15750 34264 15802
rect 34018 15748 34024 15750
rect 34080 15748 34104 15750
rect 34160 15748 34184 15750
rect 34240 15748 34264 15750
rect 34320 15748 34326 15750
rect 34018 15739 34326 15748
rect 33692 15020 33744 15026
rect 33692 14962 33744 14968
rect 33704 14618 33732 14962
rect 34532 14958 34560 16050
rect 34624 15978 34652 16526
rect 35728 16114 35756 16526
rect 36648 16250 36676 18702
rect 37476 18630 37504 19450
rect 37464 18624 37516 18630
rect 37464 18566 37516 18572
rect 36728 16992 36780 16998
rect 36728 16934 36780 16940
rect 36452 16244 36504 16250
rect 36452 16186 36504 16192
rect 36636 16244 36688 16250
rect 36636 16186 36688 16192
rect 35716 16108 35768 16114
rect 35716 16050 35768 16056
rect 34612 15972 34664 15978
rect 34612 15914 34664 15920
rect 36464 15570 36492 16186
rect 36452 15564 36504 15570
rect 36452 15506 36504 15512
rect 36740 15502 36768 16934
rect 37476 16726 37504 18566
rect 37464 16720 37516 16726
rect 37464 16662 37516 16668
rect 37476 15706 37504 16662
rect 37464 15700 37516 15706
rect 37464 15642 37516 15648
rect 36728 15496 36780 15502
rect 36728 15438 36780 15444
rect 37476 15162 37504 15642
rect 37464 15156 37516 15162
rect 37464 15098 37516 15104
rect 34520 14952 34572 14958
rect 34520 14894 34572 14900
rect 34018 14716 34326 14725
rect 34018 14714 34024 14716
rect 34080 14714 34104 14716
rect 34160 14714 34184 14716
rect 34240 14714 34264 14716
rect 34320 14714 34326 14716
rect 34080 14662 34082 14714
rect 34262 14662 34264 14714
rect 34018 14660 34024 14662
rect 34080 14660 34104 14662
rect 34160 14660 34184 14662
rect 34240 14660 34264 14662
rect 34320 14660 34326 14662
rect 34018 14651 34326 14660
rect 33692 14612 33744 14618
rect 33692 14554 33744 14560
rect 32496 14408 32548 14414
rect 32496 14350 32548 14356
rect 32508 14074 32536 14350
rect 35348 14272 35400 14278
rect 35348 14214 35400 14220
rect 32496 14068 32548 14074
rect 32496 14010 32548 14016
rect 34018 13628 34326 13637
rect 34018 13626 34024 13628
rect 34080 13626 34104 13628
rect 34160 13626 34184 13628
rect 34240 13626 34264 13628
rect 34320 13626 34326 13628
rect 34080 13574 34082 13626
rect 34262 13574 34264 13626
rect 34018 13572 34024 13574
rect 34080 13572 34104 13574
rect 34160 13572 34184 13574
rect 34240 13572 34264 13574
rect 34320 13572 34326 13574
rect 34018 13563 34326 13572
rect 35360 12850 35388 14214
rect 35348 12844 35400 12850
rect 35348 12786 35400 12792
rect 34018 12540 34326 12549
rect 34018 12538 34024 12540
rect 34080 12538 34104 12540
rect 34160 12538 34184 12540
rect 34240 12538 34264 12540
rect 34320 12538 34326 12540
rect 34080 12486 34082 12538
rect 34262 12486 34264 12538
rect 34018 12484 34024 12486
rect 34080 12484 34104 12486
rect 34160 12484 34184 12486
rect 34240 12484 34264 12486
rect 34320 12484 34326 12486
rect 34018 12475 34326 12484
rect 35360 12306 35388 12786
rect 36084 12640 36136 12646
rect 36084 12582 36136 12588
rect 36360 12640 36412 12646
rect 36360 12582 36412 12588
rect 34796 12300 34848 12306
rect 34796 12242 34848 12248
rect 35348 12300 35400 12306
rect 35348 12242 35400 12248
rect 34520 12096 34572 12102
rect 34520 12038 34572 12044
rect 34532 11558 34560 12038
rect 34520 11552 34572 11558
rect 34520 11494 34572 11500
rect 34018 11452 34326 11461
rect 34018 11450 34024 11452
rect 34080 11450 34104 11452
rect 34160 11450 34184 11452
rect 34240 11450 34264 11452
rect 34320 11450 34326 11452
rect 34080 11398 34082 11450
rect 34262 11398 34264 11450
rect 34018 11396 34024 11398
rect 34080 11396 34104 11398
rect 34160 11396 34184 11398
rect 34240 11396 34264 11398
rect 34320 11396 34326 11398
rect 34018 11387 34326 11396
rect 33692 11280 33744 11286
rect 33692 11222 33744 11228
rect 32220 11212 32272 11218
rect 32220 11154 32272 11160
rect 32036 11076 32088 11082
rect 32036 11018 32088 11024
rect 32048 10810 32076 11018
rect 32036 10804 32088 10810
rect 32036 10746 32088 10752
rect 31944 9172 31996 9178
rect 31944 9114 31996 9120
rect 31668 9104 31720 9110
rect 31668 9046 31720 9052
rect 31680 8566 31708 9046
rect 31668 8560 31720 8566
rect 31668 8502 31720 8508
rect 30840 6996 30892 7002
rect 30840 6938 30892 6944
rect 31484 6996 31536 7002
rect 31484 6938 31536 6944
rect 30748 6656 30800 6662
rect 30748 6598 30800 6604
rect 30852 6118 30880 6938
rect 31680 6798 31708 8502
rect 32048 8294 32076 10746
rect 33704 10674 33732 11222
rect 34808 10674 34836 12242
rect 36096 12238 36124 12582
rect 36084 12232 36136 12238
rect 36084 12174 36136 12180
rect 36372 12102 36400 12582
rect 35808 12096 35860 12102
rect 35808 12038 35860 12044
rect 36360 12096 36412 12102
rect 36360 12038 36412 12044
rect 35820 10810 35848 12038
rect 35808 10804 35860 10810
rect 35808 10746 35860 10752
rect 33692 10668 33744 10674
rect 33692 10610 33744 10616
rect 34796 10668 34848 10674
rect 34796 10610 34848 10616
rect 34018 10364 34326 10373
rect 34018 10362 34024 10364
rect 34080 10362 34104 10364
rect 34160 10362 34184 10364
rect 34240 10362 34264 10364
rect 34320 10362 34326 10364
rect 34080 10310 34082 10362
rect 34262 10310 34264 10362
rect 34018 10308 34024 10310
rect 34080 10308 34104 10310
rect 34160 10308 34184 10310
rect 34240 10308 34264 10310
rect 34320 10308 34326 10310
rect 34018 10299 34326 10308
rect 34808 10130 34836 10610
rect 35716 10464 35768 10470
rect 35716 10406 35768 10412
rect 34796 10124 34848 10130
rect 34796 10066 34848 10072
rect 35728 10062 35756 10406
rect 35820 10266 35848 10746
rect 35808 10260 35860 10266
rect 35808 10202 35860 10208
rect 35716 10056 35768 10062
rect 35716 9998 35768 10004
rect 34018 9276 34326 9285
rect 34018 9274 34024 9276
rect 34080 9274 34104 9276
rect 34160 9274 34184 9276
rect 34240 9274 34264 9276
rect 34320 9274 34326 9276
rect 34080 9222 34082 9274
rect 34262 9222 34264 9274
rect 34018 9220 34024 9222
rect 34080 9220 34104 9222
rect 34160 9220 34184 9222
rect 34240 9220 34264 9222
rect 34320 9220 34326 9222
rect 34018 9211 34326 9220
rect 34428 8628 34480 8634
rect 34428 8570 34480 8576
rect 33140 8424 33192 8430
rect 33140 8366 33192 8372
rect 32036 8288 32088 8294
rect 32036 8230 32088 8236
rect 32048 8090 32076 8230
rect 32036 8084 32088 8090
rect 32036 8026 32088 8032
rect 32128 8016 32180 8022
rect 32128 7958 32180 7964
rect 32036 7200 32088 7206
rect 32036 7142 32088 7148
rect 32048 6798 32076 7142
rect 31668 6792 31720 6798
rect 31668 6734 31720 6740
rect 32036 6792 32088 6798
rect 32036 6734 32088 6740
rect 31680 6458 31708 6734
rect 31668 6452 31720 6458
rect 31668 6394 31720 6400
rect 32140 6322 32168 7958
rect 32404 6656 32456 6662
rect 32404 6598 32456 6604
rect 32416 6322 32444 6598
rect 33152 6458 33180 8366
rect 33784 8356 33836 8362
rect 33784 8298 33836 8304
rect 33796 7886 33824 8298
rect 34018 8188 34326 8197
rect 34018 8186 34024 8188
rect 34080 8186 34104 8188
rect 34160 8186 34184 8188
rect 34240 8186 34264 8188
rect 34320 8186 34326 8188
rect 34080 8134 34082 8186
rect 34262 8134 34264 8186
rect 34018 8132 34024 8134
rect 34080 8132 34104 8134
rect 34160 8132 34184 8134
rect 34240 8132 34264 8134
rect 34320 8132 34326 8134
rect 34018 8123 34326 8132
rect 34440 7886 34468 8570
rect 33784 7880 33836 7886
rect 33784 7822 33836 7828
rect 34428 7880 34480 7886
rect 34428 7822 34480 7828
rect 35440 7880 35492 7886
rect 35440 7822 35492 7828
rect 33968 7744 34020 7750
rect 33968 7686 34020 7692
rect 33980 7410 34008 7686
rect 33968 7404 34020 7410
rect 33968 7346 34020 7352
rect 35452 7342 35480 7822
rect 36728 7744 36780 7750
rect 36728 7686 36780 7692
rect 36740 7546 36768 7686
rect 36452 7540 36504 7546
rect 36452 7482 36504 7488
rect 36728 7540 36780 7546
rect 36728 7482 36780 7488
rect 35440 7336 35492 7342
rect 35440 7278 35492 7284
rect 34018 7100 34326 7109
rect 34018 7098 34024 7100
rect 34080 7098 34104 7100
rect 34160 7098 34184 7100
rect 34240 7098 34264 7100
rect 34320 7098 34326 7100
rect 34080 7046 34082 7098
rect 34262 7046 34264 7098
rect 34018 7044 34024 7046
rect 34080 7044 34104 7046
rect 34160 7044 34184 7046
rect 34240 7044 34264 7046
rect 34320 7044 34326 7046
rect 34018 7035 34326 7044
rect 34888 6656 34940 6662
rect 34888 6598 34940 6604
rect 33140 6452 33192 6458
rect 33140 6394 33192 6400
rect 34900 6322 34928 6598
rect 32128 6316 32180 6322
rect 32128 6258 32180 6264
rect 32404 6316 32456 6322
rect 32404 6258 32456 6264
rect 34888 6316 34940 6322
rect 34888 6258 34940 6264
rect 35452 6254 35480 7278
rect 36464 6458 36492 7482
rect 36452 6452 36504 6458
rect 36452 6394 36504 6400
rect 35440 6248 35492 6254
rect 35440 6190 35492 6196
rect 30840 6112 30892 6118
rect 30840 6054 30892 6060
rect 30104 5908 30156 5914
rect 30104 5850 30156 5856
rect 26884 5704 26936 5710
rect 26884 5646 26936 5652
rect 27620 5704 27672 5710
rect 27620 5646 27672 5652
rect 26516 5364 26568 5370
rect 26516 5306 26568 5312
rect 24400 5092 24452 5098
rect 24400 5034 24452 5040
rect 23756 4208 23808 4214
rect 23756 4150 23808 4156
rect 24308 3936 24360 3942
rect 24308 3878 24360 3884
rect 24320 3058 24348 3878
rect 24412 3602 24440 5034
rect 24570 4924 24878 4933
rect 24570 4922 24576 4924
rect 24632 4922 24656 4924
rect 24712 4922 24736 4924
rect 24792 4922 24816 4924
rect 24872 4922 24878 4924
rect 24632 4870 24634 4922
rect 24814 4870 24816 4922
rect 24570 4868 24576 4870
rect 24632 4868 24656 4870
rect 24712 4868 24736 4870
rect 24792 4868 24816 4870
rect 24872 4868 24878 4870
rect 24570 4859 24878 4868
rect 24570 3836 24878 3845
rect 24570 3834 24576 3836
rect 24632 3834 24656 3836
rect 24712 3834 24736 3836
rect 24792 3834 24816 3836
rect 24872 3834 24878 3836
rect 24632 3782 24634 3834
rect 24814 3782 24816 3834
rect 24570 3780 24576 3782
rect 24632 3780 24656 3782
rect 24712 3780 24736 3782
rect 24792 3780 24816 3782
rect 24872 3780 24878 3782
rect 24570 3771 24878 3780
rect 26896 3602 26924 5646
rect 27160 5228 27212 5234
rect 27160 5170 27212 5176
rect 27172 4282 27200 5170
rect 27632 4622 27660 5646
rect 28540 5568 28592 5574
rect 28540 5510 28592 5516
rect 28552 4622 28580 5510
rect 29294 5468 29602 5477
rect 29294 5466 29300 5468
rect 29356 5466 29380 5468
rect 29436 5466 29460 5468
rect 29516 5466 29540 5468
rect 29596 5466 29602 5468
rect 29356 5414 29358 5466
rect 29538 5414 29540 5466
rect 29294 5412 29300 5414
rect 29356 5412 29380 5414
rect 29436 5412 29460 5414
rect 29516 5412 29540 5414
rect 29596 5412 29602 5414
rect 29294 5403 29602 5412
rect 27620 4616 27672 4622
rect 27620 4558 27672 4564
rect 28540 4616 28592 4622
rect 28540 4558 28592 4564
rect 27344 4548 27396 4554
rect 27344 4490 27396 4496
rect 27160 4276 27212 4282
rect 27160 4218 27212 4224
rect 24400 3596 24452 3602
rect 24400 3538 24452 3544
rect 26884 3596 26936 3602
rect 26884 3538 26936 3544
rect 24412 3058 24440 3538
rect 27356 3534 27384 4490
rect 27620 4480 27672 4486
rect 27620 4422 27672 4428
rect 27528 4276 27580 4282
rect 27528 4218 27580 4224
rect 27344 3528 27396 3534
rect 27344 3470 27396 3476
rect 23572 3052 23624 3058
rect 23572 2994 23624 3000
rect 24308 3052 24360 3058
rect 24308 2994 24360 3000
rect 24400 3052 24452 3058
rect 24400 2994 24452 3000
rect 27540 2922 27568 4218
rect 27632 4214 27660 4422
rect 27620 4208 27672 4214
rect 27620 4150 27672 4156
rect 27988 4140 28040 4146
rect 27988 4082 28040 4088
rect 28000 3534 28028 4082
rect 28552 3942 28580 4558
rect 29294 4380 29602 4389
rect 29294 4378 29300 4380
rect 29356 4378 29380 4380
rect 29436 4378 29460 4380
rect 29516 4378 29540 4380
rect 29596 4378 29602 4380
rect 29356 4326 29358 4378
rect 29538 4326 29540 4378
rect 29294 4324 29300 4326
rect 29356 4324 29380 4326
rect 29436 4324 29460 4326
rect 29516 4324 29540 4326
rect 29596 4324 29602 4326
rect 29294 4315 29602 4324
rect 30852 4146 30880 6054
rect 34018 6012 34326 6021
rect 34018 6010 34024 6012
rect 34080 6010 34104 6012
rect 34160 6010 34184 6012
rect 34240 6010 34264 6012
rect 34320 6010 34326 6012
rect 34080 5958 34082 6010
rect 34262 5958 34264 6010
rect 34018 5956 34024 5958
rect 34080 5956 34104 5958
rect 34160 5956 34184 5958
rect 34240 5956 34264 5958
rect 34320 5956 34326 5958
rect 34018 5947 34326 5956
rect 34018 4924 34326 4933
rect 34018 4922 34024 4924
rect 34080 4922 34104 4924
rect 34160 4922 34184 4924
rect 34240 4922 34264 4924
rect 34320 4922 34326 4924
rect 34080 4870 34082 4922
rect 34262 4870 34264 4922
rect 34018 4868 34024 4870
rect 34080 4868 34104 4870
rect 34160 4868 34184 4870
rect 34240 4868 34264 4870
rect 34320 4868 34326 4870
rect 34018 4859 34326 4868
rect 31852 4752 31904 4758
rect 31852 4694 31904 4700
rect 30840 4140 30892 4146
rect 30840 4082 30892 4088
rect 28540 3936 28592 3942
rect 28540 3878 28592 3884
rect 28552 3534 28580 3878
rect 31760 3732 31812 3738
rect 31760 3674 31812 3680
rect 31300 3664 31352 3670
rect 31300 3606 31352 3612
rect 27988 3528 28040 3534
rect 27988 3470 28040 3476
rect 28540 3528 28592 3534
rect 28540 3470 28592 3476
rect 27528 2916 27580 2922
rect 27528 2858 27580 2864
rect 24570 2748 24878 2757
rect 24570 2746 24576 2748
rect 24632 2746 24656 2748
rect 24712 2746 24736 2748
rect 24792 2746 24816 2748
rect 24872 2746 24878 2748
rect 24632 2694 24634 2746
rect 24814 2694 24816 2746
rect 24570 2692 24576 2694
rect 24632 2692 24656 2694
rect 24712 2692 24736 2694
rect 24792 2692 24816 2694
rect 24872 2692 24878 2694
rect 24570 2683 24878 2692
rect 27540 2446 27568 2858
rect 28000 2514 28028 3470
rect 29000 3460 29052 3466
rect 29000 3402 29052 3408
rect 30012 3460 30064 3466
rect 30012 3402 30064 3408
rect 28356 2848 28408 2854
rect 28356 2790 28408 2796
rect 27988 2508 28040 2514
rect 27988 2450 28040 2456
rect 28368 2446 28396 2790
rect 29012 2650 29040 3402
rect 29294 3292 29602 3301
rect 29294 3290 29300 3292
rect 29356 3290 29380 3292
rect 29436 3290 29460 3292
rect 29516 3290 29540 3292
rect 29596 3290 29602 3292
rect 29356 3238 29358 3290
rect 29538 3238 29540 3290
rect 29294 3236 29300 3238
rect 29356 3236 29380 3238
rect 29436 3236 29460 3238
rect 29516 3236 29540 3238
rect 29596 3236 29602 3238
rect 29294 3227 29602 3236
rect 30024 2650 30052 3402
rect 31024 3392 31076 3398
rect 31024 3334 31076 3340
rect 31036 3126 31064 3334
rect 31024 3120 31076 3126
rect 31024 3062 31076 3068
rect 31312 3058 31340 3606
rect 31576 3596 31628 3602
rect 31576 3538 31628 3544
rect 31392 3528 31444 3534
rect 31392 3470 31444 3476
rect 31404 3058 31432 3470
rect 31588 3126 31616 3538
rect 31576 3120 31628 3126
rect 31576 3062 31628 3068
rect 31300 3052 31352 3058
rect 31300 2994 31352 3000
rect 31392 3052 31444 3058
rect 31392 2994 31444 3000
rect 31772 2650 31800 3674
rect 31864 3534 31892 4694
rect 34018 3836 34326 3845
rect 34018 3834 34024 3836
rect 34080 3834 34104 3836
rect 34160 3834 34184 3836
rect 34240 3834 34264 3836
rect 34320 3834 34326 3836
rect 34080 3782 34082 3834
rect 34262 3782 34264 3834
rect 34018 3780 34024 3782
rect 34080 3780 34104 3782
rect 34160 3780 34184 3782
rect 34240 3780 34264 3782
rect 34320 3780 34326 3782
rect 34018 3771 34326 3780
rect 36820 3732 36872 3738
rect 36820 3674 36872 3680
rect 33692 3596 33744 3602
rect 33692 3538 33744 3544
rect 31852 3528 31904 3534
rect 31852 3470 31904 3476
rect 32404 3528 32456 3534
rect 32404 3470 32456 3476
rect 31944 2848 31996 2854
rect 31944 2790 31996 2796
rect 29000 2644 29052 2650
rect 29000 2586 29052 2592
rect 30012 2644 30064 2650
rect 30012 2586 30064 2592
rect 31760 2644 31812 2650
rect 31760 2586 31812 2592
rect 31956 2446 31984 2790
rect 32416 2650 32444 3470
rect 33232 3460 33284 3466
rect 33232 3402 33284 3408
rect 33244 2650 33272 3402
rect 33704 2650 33732 3538
rect 34520 2848 34572 2854
rect 34520 2790 34572 2796
rect 36728 2848 36780 2854
rect 36728 2790 36780 2796
rect 34018 2748 34326 2757
rect 34018 2746 34024 2748
rect 34080 2746 34104 2748
rect 34160 2746 34184 2748
rect 34240 2746 34264 2748
rect 34320 2746 34326 2748
rect 34080 2694 34082 2746
rect 34262 2694 34264 2746
rect 34018 2692 34024 2694
rect 34080 2692 34104 2694
rect 34160 2692 34184 2694
rect 34240 2692 34264 2694
rect 34320 2692 34326 2694
rect 34018 2683 34326 2692
rect 32404 2644 32456 2650
rect 32404 2586 32456 2592
rect 33232 2644 33284 2650
rect 33232 2586 33284 2592
rect 33692 2644 33744 2650
rect 33692 2586 33744 2592
rect 34532 2446 34560 2790
rect 23572 2440 23624 2446
rect 23492 2400 23572 2428
rect 22376 2382 22428 2388
rect 23572 2382 23624 2388
rect 27528 2440 27580 2446
rect 27528 2382 27580 2388
rect 28356 2440 28408 2446
rect 28356 2382 28408 2388
rect 29644 2440 29696 2446
rect 29644 2382 29696 2388
rect 30748 2440 30800 2446
rect 30748 2382 30800 2388
rect 31944 2440 31996 2446
rect 31944 2382 31996 2388
rect 33140 2440 33192 2446
rect 34520 2440 34572 2446
rect 33140 2382 33192 2388
rect 34348 2388 34520 2394
rect 34348 2382 34572 2388
rect 35532 2440 35584 2446
rect 35532 2382 35584 2388
rect 19708 2372 19760 2378
rect 19708 2314 19760 2320
rect 18788 2304 18840 2310
rect 18788 2246 18840 2252
rect 18800 800 18828 2246
rect 19846 2204 20154 2213
rect 19846 2202 19852 2204
rect 19908 2202 19932 2204
rect 19988 2202 20012 2204
rect 20068 2202 20092 2204
rect 20148 2202 20154 2204
rect 19908 2150 19910 2202
rect 20090 2150 20092 2202
rect 19846 2148 19852 2150
rect 19908 2148 19932 2150
rect 19988 2148 20012 2150
rect 20068 2148 20092 2150
rect 20148 2148 20154 2150
rect 19846 2139 20154 2148
rect 19996 870 20116 898
rect 19996 800 20024 870
rect 846 0 902 800
rect 2042 0 2098 800
rect 3238 0 3294 800
rect 4434 0 4490 800
rect 5630 0 5686 800
rect 6826 0 6882 800
rect 8022 0 8078 800
rect 9218 0 9274 800
rect 10414 0 10470 800
rect 11610 0 11666 800
rect 12806 0 12862 800
rect 14002 0 14058 800
rect 15198 0 15254 800
rect 16394 0 16450 800
rect 17590 0 17646 800
rect 18786 0 18842 800
rect 19982 0 20038 800
rect 20088 762 20116 870
rect 20272 762 20300 2382
rect 21180 2304 21232 2310
rect 21180 2246 21232 2252
rect 21192 800 21220 2246
rect 22388 800 22416 2382
rect 23584 800 23612 2382
rect 24768 2304 24820 2310
rect 24768 2246 24820 2252
rect 27160 2304 27212 2310
rect 27160 2246 27212 2252
rect 24780 800 24808 2246
rect 27172 800 27200 2246
rect 28368 800 28396 2382
rect 29294 2204 29602 2213
rect 29294 2202 29300 2204
rect 29356 2202 29380 2204
rect 29436 2202 29460 2204
rect 29516 2202 29540 2204
rect 29596 2202 29602 2204
rect 29356 2150 29358 2202
rect 29538 2150 29540 2202
rect 29294 2148 29300 2150
rect 29356 2148 29380 2150
rect 29436 2148 29460 2150
rect 29516 2148 29540 2150
rect 29596 2148 29602 2150
rect 29294 2139 29602 2148
rect 29656 1578 29684 2382
rect 29564 1550 29684 1578
rect 29564 800 29592 1550
rect 30760 800 30788 2382
rect 31956 800 31984 2382
rect 33152 800 33180 2382
rect 34348 2366 34560 2382
rect 34348 800 34376 2366
rect 35544 800 35572 2382
rect 36740 800 36768 2790
rect 36832 2650 36860 3674
rect 37924 3528 37976 3534
rect 37924 3470 37976 3476
rect 37648 3460 37700 3466
rect 37648 3402 37700 3408
rect 37280 3392 37332 3398
rect 37280 3334 37332 3340
rect 37292 2650 37320 3334
rect 37464 2848 37516 2854
rect 37464 2790 37516 2796
rect 36820 2644 36872 2650
rect 36820 2586 36872 2592
rect 37280 2644 37332 2650
rect 37280 2586 37332 2592
rect 37476 2446 37504 2790
rect 37660 2650 37688 3402
rect 37936 3194 37964 3470
rect 38108 3392 38160 3398
rect 38108 3334 38160 3340
rect 37924 3188 37976 3194
rect 37924 3130 37976 3136
rect 38120 3058 38148 3334
rect 38108 3052 38160 3058
rect 38108 2994 38160 3000
rect 39120 3052 39172 3058
rect 39120 2994 39172 3000
rect 38016 2984 38068 2990
rect 38016 2926 38068 2932
rect 37648 2644 37700 2650
rect 37648 2586 37700 2592
rect 38028 2446 38056 2926
rect 37464 2440 37516 2446
rect 38016 2440 38068 2446
rect 37464 2382 37516 2388
rect 37936 2400 38016 2428
rect 37936 800 37964 2400
rect 38016 2382 38068 2388
rect 39132 800 39160 2994
rect 20088 734 20300 762
rect 21178 0 21234 800
rect 22374 0 22430 800
rect 23570 0 23626 800
rect 24766 0 24822 800
rect 25962 0 26018 800
rect 27158 0 27214 800
rect 28354 0 28410 800
rect 29550 0 29606 800
rect 30746 0 30802 800
rect 31942 0 31998 800
rect 33138 0 33194 800
rect 34334 0 34390 800
rect 35530 0 35586 800
rect 36726 0 36782 800
rect 37922 0 37978 800
rect 39118 0 39174 800
<< via2 >>
rect 1398 34312 1454 34368
rect 1490 32952 1546 33008
rect 1490 31628 1492 31648
rect 1492 31628 1544 31648
rect 1544 31628 1546 31648
rect 1490 31592 1546 31628
rect 1490 30232 1546 30288
rect 1490 28872 1546 28928
rect 1490 27512 1546 27568
rect 10404 33754 10460 33756
rect 10484 33754 10540 33756
rect 10564 33754 10620 33756
rect 10644 33754 10700 33756
rect 10404 33702 10450 33754
rect 10450 33702 10460 33754
rect 10484 33702 10514 33754
rect 10514 33702 10526 33754
rect 10526 33702 10540 33754
rect 10564 33702 10578 33754
rect 10578 33702 10590 33754
rect 10590 33702 10620 33754
rect 10644 33702 10654 33754
rect 10654 33702 10700 33754
rect 10404 33700 10460 33702
rect 10484 33700 10540 33702
rect 10564 33700 10620 33702
rect 10644 33700 10700 33702
rect 19852 33754 19908 33756
rect 19932 33754 19988 33756
rect 20012 33754 20068 33756
rect 20092 33754 20148 33756
rect 19852 33702 19898 33754
rect 19898 33702 19908 33754
rect 19932 33702 19962 33754
rect 19962 33702 19974 33754
rect 19974 33702 19988 33754
rect 20012 33702 20026 33754
rect 20026 33702 20038 33754
rect 20038 33702 20068 33754
rect 20092 33702 20102 33754
rect 20102 33702 20148 33754
rect 19852 33700 19908 33702
rect 19932 33700 19988 33702
rect 20012 33700 20068 33702
rect 20092 33700 20148 33702
rect 5680 33210 5736 33212
rect 5760 33210 5816 33212
rect 5840 33210 5896 33212
rect 5920 33210 5976 33212
rect 5680 33158 5726 33210
rect 5726 33158 5736 33210
rect 5760 33158 5790 33210
rect 5790 33158 5802 33210
rect 5802 33158 5816 33210
rect 5840 33158 5854 33210
rect 5854 33158 5866 33210
rect 5866 33158 5896 33210
rect 5920 33158 5930 33210
rect 5930 33158 5976 33210
rect 5680 33156 5736 33158
rect 5760 33156 5816 33158
rect 5840 33156 5896 33158
rect 5920 33156 5976 33158
rect 29300 33754 29356 33756
rect 29380 33754 29436 33756
rect 29460 33754 29516 33756
rect 29540 33754 29596 33756
rect 29300 33702 29346 33754
rect 29346 33702 29356 33754
rect 29380 33702 29410 33754
rect 29410 33702 29422 33754
rect 29422 33702 29436 33754
rect 29460 33702 29474 33754
rect 29474 33702 29486 33754
rect 29486 33702 29516 33754
rect 29540 33702 29550 33754
rect 29550 33702 29596 33754
rect 29300 33700 29356 33702
rect 29380 33700 29436 33702
rect 29460 33700 29516 33702
rect 29540 33700 29596 33702
rect 1490 26188 1492 26208
rect 1492 26188 1544 26208
rect 1544 26188 1546 26208
rect 1490 26152 1546 26188
rect 1490 24792 1546 24848
rect 1490 23468 1492 23488
rect 1492 23468 1544 23488
rect 1544 23468 1546 23488
rect 1490 23432 1546 23468
rect 1398 22072 1454 22128
rect 1490 20748 1492 20768
rect 1492 20748 1544 20768
rect 1544 20748 1546 20768
rect 1490 20712 1546 20748
rect 1490 19352 1546 19408
rect 1490 18028 1492 18048
rect 1492 18028 1544 18048
rect 1544 18028 1546 18048
rect 1490 17992 1546 18028
rect 1490 16632 1546 16688
rect 1490 15308 1492 15328
rect 1492 15308 1544 15328
rect 1544 15308 1546 15328
rect 1490 15272 1546 15308
rect 1490 13912 1546 13968
rect 1490 12588 1492 12608
rect 1492 12588 1544 12608
rect 1544 12588 1546 12608
rect 1490 12552 1546 12588
rect 1490 11192 1546 11248
rect 1490 9868 1492 9888
rect 1492 9868 1544 9888
rect 1544 9868 1546 9888
rect 1490 9832 1546 9868
rect 1490 8472 1546 8528
rect 1490 7148 1492 7168
rect 1492 7148 1544 7168
rect 1544 7148 1546 7168
rect 1490 7112 1546 7148
rect 5680 32122 5736 32124
rect 5760 32122 5816 32124
rect 5840 32122 5896 32124
rect 5920 32122 5976 32124
rect 5680 32070 5726 32122
rect 5726 32070 5736 32122
rect 5760 32070 5790 32122
rect 5790 32070 5802 32122
rect 5802 32070 5816 32122
rect 5840 32070 5854 32122
rect 5854 32070 5866 32122
rect 5866 32070 5896 32122
rect 5920 32070 5930 32122
rect 5930 32070 5976 32122
rect 5680 32068 5736 32070
rect 5760 32068 5816 32070
rect 5840 32068 5896 32070
rect 5920 32068 5976 32070
rect 5680 31034 5736 31036
rect 5760 31034 5816 31036
rect 5840 31034 5896 31036
rect 5920 31034 5976 31036
rect 5680 30982 5726 31034
rect 5726 30982 5736 31034
rect 5760 30982 5790 31034
rect 5790 30982 5802 31034
rect 5802 30982 5816 31034
rect 5840 30982 5854 31034
rect 5854 30982 5866 31034
rect 5866 30982 5896 31034
rect 5920 30982 5930 31034
rect 5930 30982 5976 31034
rect 5680 30980 5736 30982
rect 5760 30980 5816 30982
rect 5840 30980 5896 30982
rect 5920 30980 5976 30982
rect 5680 29946 5736 29948
rect 5760 29946 5816 29948
rect 5840 29946 5896 29948
rect 5920 29946 5976 29948
rect 5680 29894 5726 29946
rect 5726 29894 5736 29946
rect 5760 29894 5790 29946
rect 5790 29894 5802 29946
rect 5802 29894 5816 29946
rect 5840 29894 5854 29946
rect 5854 29894 5866 29946
rect 5866 29894 5896 29946
rect 5920 29894 5930 29946
rect 5930 29894 5976 29946
rect 5680 29892 5736 29894
rect 5760 29892 5816 29894
rect 5840 29892 5896 29894
rect 5920 29892 5976 29894
rect 1490 5752 1546 5808
rect 1490 4428 1492 4448
rect 1492 4428 1544 4448
rect 1544 4428 1546 4448
rect 1490 4392 1546 4428
rect 5680 28858 5736 28860
rect 5760 28858 5816 28860
rect 5840 28858 5896 28860
rect 5920 28858 5976 28860
rect 5680 28806 5726 28858
rect 5726 28806 5736 28858
rect 5760 28806 5790 28858
rect 5790 28806 5802 28858
rect 5802 28806 5816 28858
rect 5840 28806 5854 28858
rect 5854 28806 5866 28858
rect 5866 28806 5896 28858
rect 5920 28806 5930 28858
rect 5930 28806 5976 28858
rect 5680 28804 5736 28806
rect 5760 28804 5816 28806
rect 5840 28804 5896 28806
rect 5920 28804 5976 28806
rect 5680 27770 5736 27772
rect 5760 27770 5816 27772
rect 5840 27770 5896 27772
rect 5920 27770 5976 27772
rect 5680 27718 5726 27770
rect 5726 27718 5736 27770
rect 5760 27718 5790 27770
rect 5790 27718 5802 27770
rect 5802 27718 5816 27770
rect 5840 27718 5854 27770
rect 5854 27718 5866 27770
rect 5866 27718 5896 27770
rect 5920 27718 5930 27770
rect 5930 27718 5976 27770
rect 5680 27716 5736 27718
rect 5760 27716 5816 27718
rect 5840 27716 5896 27718
rect 5920 27716 5976 27718
rect 5680 26682 5736 26684
rect 5760 26682 5816 26684
rect 5840 26682 5896 26684
rect 5920 26682 5976 26684
rect 5680 26630 5726 26682
rect 5726 26630 5736 26682
rect 5760 26630 5790 26682
rect 5790 26630 5802 26682
rect 5802 26630 5816 26682
rect 5840 26630 5854 26682
rect 5854 26630 5866 26682
rect 5866 26630 5896 26682
rect 5920 26630 5930 26682
rect 5930 26630 5976 26682
rect 5680 26628 5736 26630
rect 5760 26628 5816 26630
rect 5840 26628 5896 26630
rect 5920 26628 5976 26630
rect 5680 25594 5736 25596
rect 5760 25594 5816 25596
rect 5840 25594 5896 25596
rect 5920 25594 5976 25596
rect 5680 25542 5726 25594
rect 5726 25542 5736 25594
rect 5760 25542 5790 25594
rect 5790 25542 5802 25594
rect 5802 25542 5816 25594
rect 5840 25542 5854 25594
rect 5854 25542 5866 25594
rect 5866 25542 5896 25594
rect 5920 25542 5930 25594
rect 5930 25542 5976 25594
rect 5680 25540 5736 25542
rect 5760 25540 5816 25542
rect 5840 25540 5896 25542
rect 5920 25540 5976 25542
rect 5680 24506 5736 24508
rect 5760 24506 5816 24508
rect 5840 24506 5896 24508
rect 5920 24506 5976 24508
rect 5680 24454 5726 24506
rect 5726 24454 5736 24506
rect 5760 24454 5790 24506
rect 5790 24454 5802 24506
rect 5802 24454 5816 24506
rect 5840 24454 5854 24506
rect 5854 24454 5866 24506
rect 5866 24454 5896 24506
rect 5920 24454 5930 24506
rect 5930 24454 5976 24506
rect 5680 24452 5736 24454
rect 5760 24452 5816 24454
rect 5840 24452 5896 24454
rect 5920 24452 5976 24454
rect 5680 23418 5736 23420
rect 5760 23418 5816 23420
rect 5840 23418 5896 23420
rect 5920 23418 5976 23420
rect 5680 23366 5726 23418
rect 5726 23366 5736 23418
rect 5760 23366 5790 23418
rect 5790 23366 5802 23418
rect 5802 23366 5816 23418
rect 5840 23366 5854 23418
rect 5854 23366 5866 23418
rect 5866 23366 5896 23418
rect 5920 23366 5930 23418
rect 5930 23366 5976 23418
rect 5680 23364 5736 23366
rect 5760 23364 5816 23366
rect 5840 23364 5896 23366
rect 5920 23364 5976 23366
rect 5680 22330 5736 22332
rect 5760 22330 5816 22332
rect 5840 22330 5896 22332
rect 5920 22330 5976 22332
rect 5680 22278 5726 22330
rect 5726 22278 5736 22330
rect 5760 22278 5790 22330
rect 5790 22278 5802 22330
rect 5802 22278 5816 22330
rect 5840 22278 5854 22330
rect 5854 22278 5866 22330
rect 5866 22278 5896 22330
rect 5920 22278 5930 22330
rect 5930 22278 5976 22330
rect 5680 22276 5736 22278
rect 5760 22276 5816 22278
rect 5840 22276 5896 22278
rect 5920 22276 5976 22278
rect 5680 21242 5736 21244
rect 5760 21242 5816 21244
rect 5840 21242 5896 21244
rect 5920 21242 5976 21244
rect 5680 21190 5726 21242
rect 5726 21190 5736 21242
rect 5760 21190 5790 21242
rect 5790 21190 5802 21242
rect 5802 21190 5816 21242
rect 5840 21190 5854 21242
rect 5854 21190 5866 21242
rect 5866 21190 5896 21242
rect 5920 21190 5930 21242
rect 5930 21190 5976 21242
rect 5680 21188 5736 21190
rect 5760 21188 5816 21190
rect 5840 21188 5896 21190
rect 5920 21188 5976 21190
rect 5680 20154 5736 20156
rect 5760 20154 5816 20156
rect 5840 20154 5896 20156
rect 5920 20154 5976 20156
rect 5680 20102 5726 20154
rect 5726 20102 5736 20154
rect 5760 20102 5790 20154
rect 5790 20102 5802 20154
rect 5802 20102 5816 20154
rect 5840 20102 5854 20154
rect 5854 20102 5866 20154
rect 5866 20102 5896 20154
rect 5920 20102 5930 20154
rect 5930 20102 5976 20154
rect 5680 20100 5736 20102
rect 5760 20100 5816 20102
rect 5840 20100 5896 20102
rect 5920 20100 5976 20102
rect 5680 19066 5736 19068
rect 5760 19066 5816 19068
rect 5840 19066 5896 19068
rect 5920 19066 5976 19068
rect 5680 19014 5726 19066
rect 5726 19014 5736 19066
rect 5760 19014 5790 19066
rect 5790 19014 5802 19066
rect 5802 19014 5816 19066
rect 5840 19014 5854 19066
rect 5854 19014 5866 19066
rect 5866 19014 5896 19066
rect 5920 19014 5930 19066
rect 5930 19014 5976 19066
rect 5680 19012 5736 19014
rect 5760 19012 5816 19014
rect 5840 19012 5896 19014
rect 5920 19012 5976 19014
rect 5680 17978 5736 17980
rect 5760 17978 5816 17980
rect 5840 17978 5896 17980
rect 5920 17978 5976 17980
rect 5680 17926 5726 17978
rect 5726 17926 5736 17978
rect 5760 17926 5790 17978
rect 5790 17926 5802 17978
rect 5802 17926 5816 17978
rect 5840 17926 5854 17978
rect 5854 17926 5866 17978
rect 5866 17926 5896 17978
rect 5920 17926 5930 17978
rect 5930 17926 5976 17978
rect 5680 17924 5736 17926
rect 5760 17924 5816 17926
rect 5840 17924 5896 17926
rect 5920 17924 5976 17926
rect 5680 16890 5736 16892
rect 5760 16890 5816 16892
rect 5840 16890 5896 16892
rect 5920 16890 5976 16892
rect 5680 16838 5726 16890
rect 5726 16838 5736 16890
rect 5760 16838 5790 16890
rect 5790 16838 5802 16890
rect 5802 16838 5816 16890
rect 5840 16838 5854 16890
rect 5854 16838 5866 16890
rect 5866 16838 5896 16890
rect 5920 16838 5930 16890
rect 5930 16838 5976 16890
rect 5680 16836 5736 16838
rect 5760 16836 5816 16838
rect 5840 16836 5896 16838
rect 5920 16836 5976 16838
rect 5680 15802 5736 15804
rect 5760 15802 5816 15804
rect 5840 15802 5896 15804
rect 5920 15802 5976 15804
rect 5680 15750 5726 15802
rect 5726 15750 5736 15802
rect 5760 15750 5790 15802
rect 5790 15750 5802 15802
rect 5802 15750 5816 15802
rect 5840 15750 5854 15802
rect 5854 15750 5866 15802
rect 5866 15750 5896 15802
rect 5920 15750 5930 15802
rect 5930 15750 5976 15802
rect 5680 15748 5736 15750
rect 5760 15748 5816 15750
rect 5840 15748 5896 15750
rect 5920 15748 5976 15750
rect 5680 14714 5736 14716
rect 5760 14714 5816 14716
rect 5840 14714 5896 14716
rect 5920 14714 5976 14716
rect 5680 14662 5726 14714
rect 5726 14662 5736 14714
rect 5760 14662 5790 14714
rect 5790 14662 5802 14714
rect 5802 14662 5816 14714
rect 5840 14662 5854 14714
rect 5854 14662 5866 14714
rect 5866 14662 5896 14714
rect 5920 14662 5930 14714
rect 5930 14662 5976 14714
rect 5680 14660 5736 14662
rect 5760 14660 5816 14662
rect 5840 14660 5896 14662
rect 5920 14660 5976 14662
rect 5680 13626 5736 13628
rect 5760 13626 5816 13628
rect 5840 13626 5896 13628
rect 5920 13626 5976 13628
rect 5680 13574 5726 13626
rect 5726 13574 5736 13626
rect 5760 13574 5790 13626
rect 5790 13574 5802 13626
rect 5802 13574 5816 13626
rect 5840 13574 5854 13626
rect 5854 13574 5866 13626
rect 5866 13574 5896 13626
rect 5920 13574 5930 13626
rect 5930 13574 5976 13626
rect 5680 13572 5736 13574
rect 5760 13572 5816 13574
rect 5840 13572 5896 13574
rect 5920 13572 5976 13574
rect 5680 12538 5736 12540
rect 5760 12538 5816 12540
rect 5840 12538 5896 12540
rect 5920 12538 5976 12540
rect 5680 12486 5726 12538
rect 5726 12486 5736 12538
rect 5760 12486 5790 12538
rect 5790 12486 5802 12538
rect 5802 12486 5816 12538
rect 5840 12486 5854 12538
rect 5854 12486 5866 12538
rect 5866 12486 5896 12538
rect 5920 12486 5930 12538
rect 5930 12486 5976 12538
rect 5680 12484 5736 12486
rect 5760 12484 5816 12486
rect 5840 12484 5896 12486
rect 5920 12484 5976 12486
rect 1490 3032 1546 3088
rect 5680 11450 5736 11452
rect 5760 11450 5816 11452
rect 5840 11450 5896 11452
rect 5920 11450 5976 11452
rect 5680 11398 5726 11450
rect 5726 11398 5736 11450
rect 5760 11398 5790 11450
rect 5790 11398 5802 11450
rect 5802 11398 5816 11450
rect 5840 11398 5854 11450
rect 5854 11398 5866 11450
rect 5866 11398 5896 11450
rect 5920 11398 5930 11450
rect 5930 11398 5976 11450
rect 5680 11396 5736 11398
rect 5760 11396 5816 11398
rect 5840 11396 5896 11398
rect 5920 11396 5976 11398
rect 5680 10362 5736 10364
rect 5760 10362 5816 10364
rect 5840 10362 5896 10364
rect 5920 10362 5976 10364
rect 5680 10310 5726 10362
rect 5726 10310 5736 10362
rect 5760 10310 5790 10362
rect 5790 10310 5802 10362
rect 5802 10310 5816 10362
rect 5840 10310 5854 10362
rect 5854 10310 5866 10362
rect 5866 10310 5896 10362
rect 5920 10310 5930 10362
rect 5930 10310 5976 10362
rect 5680 10308 5736 10310
rect 5760 10308 5816 10310
rect 5840 10308 5896 10310
rect 5920 10308 5976 10310
rect 5680 9274 5736 9276
rect 5760 9274 5816 9276
rect 5840 9274 5896 9276
rect 5920 9274 5976 9276
rect 5680 9222 5726 9274
rect 5726 9222 5736 9274
rect 5760 9222 5790 9274
rect 5790 9222 5802 9274
rect 5802 9222 5816 9274
rect 5840 9222 5854 9274
rect 5854 9222 5866 9274
rect 5866 9222 5896 9274
rect 5920 9222 5930 9274
rect 5930 9222 5976 9274
rect 5680 9220 5736 9222
rect 5760 9220 5816 9222
rect 5840 9220 5896 9222
rect 5920 9220 5976 9222
rect 5680 8186 5736 8188
rect 5760 8186 5816 8188
rect 5840 8186 5896 8188
rect 5920 8186 5976 8188
rect 5680 8134 5726 8186
rect 5726 8134 5736 8186
rect 5760 8134 5790 8186
rect 5790 8134 5802 8186
rect 5802 8134 5816 8186
rect 5840 8134 5854 8186
rect 5854 8134 5866 8186
rect 5866 8134 5896 8186
rect 5920 8134 5930 8186
rect 5930 8134 5976 8186
rect 5680 8132 5736 8134
rect 5760 8132 5816 8134
rect 5840 8132 5896 8134
rect 5920 8132 5976 8134
rect 5680 7098 5736 7100
rect 5760 7098 5816 7100
rect 5840 7098 5896 7100
rect 5920 7098 5976 7100
rect 5680 7046 5726 7098
rect 5726 7046 5736 7098
rect 5760 7046 5790 7098
rect 5790 7046 5802 7098
rect 5802 7046 5816 7098
rect 5840 7046 5854 7098
rect 5854 7046 5866 7098
rect 5866 7046 5896 7098
rect 5920 7046 5930 7098
rect 5930 7046 5976 7098
rect 5680 7044 5736 7046
rect 5760 7044 5816 7046
rect 5840 7044 5896 7046
rect 5920 7044 5976 7046
rect 5680 6010 5736 6012
rect 5760 6010 5816 6012
rect 5840 6010 5896 6012
rect 5920 6010 5976 6012
rect 5680 5958 5726 6010
rect 5726 5958 5736 6010
rect 5760 5958 5790 6010
rect 5790 5958 5802 6010
rect 5802 5958 5816 6010
rect 5840 5958 5854 6010
rect 5854 5958 5866 6010
rect 5866 5958 5896 6010
rect 5920 5958 5930 6010
rect 5930 5958 5976 6010
rect 5680 5956 5736 5958
rect 5760 5956 5816 5958
rect 5840 5956 5896 5958
rect 5920 5956 5976 5958
rect 5680 4922 5736 4924
rect 5760 4922 5816 4924
rect 5840 4922 5896 4924
rect 5920 4922 5976 4924
rect 5680 4870 5726 4922
rect 5726 4870 5736 4922
rect 5760 4870 5790 4922
rect 5790 4870 5802 4922
rect 5802 4870 5816 4922
rect 5840 4870 5854 4922
rect 5854 4870 5866 4922
rect 5866 4870 5896 4922
rect 5920 4870 5930 4922
rect 5930 4870 5976 4922
rect 5680 4868 5736 4870
rect 5760 4868 5816 4870
rect 5840 4868 5896 4870
rect 5920 4868 5976 4870
rect 5680 3834 5736 3836
rect 5760 3834 5816 3836
rect 5840 3834 5896 3836
rect 5920 3834 5976 3836
rect 5680 3782 5726 3834
rect 5726 3782 5736 3834
rect 5760 3782 5790 3834
rect 5790 3782 5802 3834
rect 5802 3782 5816 3834
rect 5840 3782 5854 3834
rect 5854 3782 5866 3834
rect 5866 3782 5896 3834
rect 5920 3782 5930 3834
rect 5930 3782 5976 3834
rect 5680 3780 5736 3782
rect 5760 3780 5816 3782
rect 5840 3780 5896 3782
rect 5920 3780 5976 3782
rect 5680 2746 5736 2748
rect 5760 2746 5816 2748
rect 5840 2746 5896 2748
rect 5920 2746 5976 2748
rect 5680 2694 5726 2746
rect 5726 2694 5736 2746
rect 5760 2694 5790 2746
rect 5790 2694 5802 2746
rect 5802 2694 5816 2746
rect 5840 2694 5854 2746
rect 5854 2694 5866 2746
rect 5866 2694 5896 2746
rect 5920 2694 5930 2746
rect 5930 2694 5976 2746
rect 5680 2692 5736 2694
rect 5760 2692 5816 2694
rect 5840 2692 5896 2694
rect 5920 2692 5976 2694
rect 10404 32666 10460 32668
rect 10484 32666 10540 32668
rect 10564 32666 10620 32668
rect 10644 32666 10700 32668
rect 10404 32614 10450 32666
rect 10450 32614 10460 32666
rect 10484 32614 10514 32666
rect 10514 32614 10526 32666
rect 10526 32614 10540 32666
rect 10564 32614 10578 32666
rect 10578 32614 10590 32666
rect 10590 32614 10620 32666
rect 10644 32614 10654 32666
rect 10654 32614 10700 32666
rect 10404 32612 10460 32614
rect 10484 32612 10540 32614
rect 10564 32612 10620 32614
rect 10644 32612 10700 32614
rect 10404 31578 10460 31580
rect 10484 31578 10540 31580
rect 10564 31578 10620 31580
rect 10644 31578 10700 31580
rect 10404 31526 10450 31578
rect 10450 31526 10460 31578
rect 10484 31526 10514 31578
rect 10514 31526 10526 31578
rect 10526 31526 10540 31578
rect 10564 31526 10578 31578
rect 10578 31526 10590 31578
rect 10590 31526 10620 31578
rect 10644 31526 10654 31578
rect 10654 31526 10700 31578
rect 10404 31524 10460 31526
rect 10484 31524 10540 31526
rect 10564 31524 10620 31526
rect 10644 31524 10700 31526
rect 10404 30490 10460 30492
rect 10484 30490 10540 30492
rect 10564 30490 10620 30492
rect 10644 30490 10700 30492
rect 10404 30438 10450 30490
rect 10450 30438 10460 30490
rect 10484 30438 10514 30490
rect 10514 30438 10526 30490
rect 10526 30438 10540 30490
rect 10564 30438 10578 30490
rect 10578 30438 10590 30490
rect 10590 30438 10620 30490
rect 10644 30438 10654 30490
rect 10654 30438 10700 30490
rect 10404 30436 10460 30438
rect 10484 30436 10540 30438
rect 10564 30436 10620 30438
rect 10644 30436 10700 30438
rect 10404 29402 10460 29404
rect 10484 29402 10540 29404
rect 10564 29402 10620 29404
rect 10644 29402 10700 29404
rect 10404 29350 10450 29402
rect 10450 29350 10460 29402
rect 10484 29350 10514 29402
rect 10514 29350 10526 29402
rect 10526 29350 10540 29402
rect 10564 29350 10578 29402
rect 10578 29350 10590 29402
rect 10590 29350 10620 29402
rect 10644 29350 10654 29402
rect 10654 29350 10700 29402
rect 10404 29348 10460 29350
rect 10484 29348 10540 29350
rect 10564 29348 10620 29350
rect 10644 29348 10700 29350
rect 10404 28314 10460 28316
rect 10484 28314 10540 28316
rect 10564 28314 10620 28316
rect 10644 28314 10700 28316
rect 10404 28262 10450 28314
rect 10450 28262 10460 28314
rect 10484 28262 10514 28314
rect 10514 28262 10526 28314
rect 10526 28262 10540 28314
rect 10564 28262 10578 28314
rect 10578 28262 10590 28314
rect 10590 28262 10620 28314
rect 10644 28262 10654 28314
rect 10654 28262 10700 28314
rect 10404 28260 10460 28262
rect 10484 28260 10540 28262
rect 10564 28260 10620 28262
rect 10644 28260 10700 28262
rect 10404 27226 10460 27228
rect 10484 27226 10540 27228
rect 10564 27226 10620 27228
rect 10644 27226 10700 27228
rect 10404 27174 10450 27226
rect 10450 27174 10460 27226
rect 10484 27174 10514 27226
rect 10514 27174 10526 27226
rect 10526 27174 10540 27226
rect 10564 27174 10578 27226
rect 10578 27174 10590 27226
rect 10590 27174 10620 27226
rect 10644 27174 10654 27226
rect 10654 27174 10700 27226
rect 10404 27172 10460 27174
rect 10484 27172 10540 27174
rect 10564 27172 10620 27174
rect 10644 27172 10700 27174
rect 10404 26138 10460 26140
rect 10484 26138 10540 26140
rect 10564 26138 10620 26140
rect 10644 26138 10700 26140
rect 10404 26086 10450 26138
rect 10450 26086 10460 26138
rect 10484 26086 10514 26138
rect 10514 26086 10526 26138
rect 10526 26086 10540 26138
rect 10564 26086 10578 26138
rect 10578 26086 10590 26138
rect 10590 26086 10620 26138
rect 10644 26086 10654 26138
rect 10654 26086 10700 26138
rect 10404 26084 10460 26086
rect 10484 26084 10540 26086
rect 10564 26084 10620 26086
rect 10644 26084 10700 26086
rect 10404 25050 10460 25052
rect 10484 25050 10540 25052
rect 10564 25050 10620 25052
rect 10644 25050 10700 25052
rect 10404 24998 10450 25050
rect 10450 24998 10460 25050
rect 10484 24998 10514 25050
rect 10514 24998 10526 25050
rect 10526 24998 10540 25050
rect 10564 24998 10578 25050
rect 10578 24998 10590 25050
rect 10590 24998 10620 25050
rect 10644 24998 10654 25050
rect 10654 24998 10700 25050
rect 10404 24996 10460 24998
rect 10484 24996 10540 24998
rect 10564 24996 10620 24998
rect 10644 24996 10700 24998
rect 10404 23962 10460 23964
rect 10484 23962 10540 23964
rect 10564 23962 10620 23964
rect 10644 23962 10700 23964
rect 10404 23910 10450 23962
rect 10450 23910 10460 23962
rect 10484 23910 10514 23962
rect 10514 23910 10526 23962
rect 10526 23910 10540 23962
rect 10564 23910 10578 23962
rect 10578 23910 10590 23962
rect 10590 23910 10620 23962
rect 10644 23910 10654 23962
rect 10654 23910 10700 23962
rect 10404 23908 10460 23910
rect 10484 23908 10540 23910
rect 10564 23908 10620 23910
rect 10644 23908 10700 23910
rect 10404 22874 10460 22876
rect 10484 22874 10540 22876
rect 10564 22874 10620 22876
rect 10644 22874 10700 22876
rect 10404 22822 10450 22874
rect 10450 22822 10460 22874
rect 10484 22822 10514 22874
rect 10514 22822 10526 22874
rect 10526 22822 10540 22874
rect 10564 22822 10578 22874
rect 10578 22822 10590 22874
rect 10590 22822 10620 22874
rect 10644 22822 10654 22874
rect 10654 22822 10700 22874
rect 10404 22820 10460 22822
rect 10484 22820 10540 22822
rect 10564 22820 10620 22822
rect 10644 22820 10700 22822
rect 10404 21786 10460 21788
rect 10484 21786 10540 21788
rect 10564 21786 10620 21788
rect 10644 21786 10700 21788
rect 10404 21734 10450 21786
rect 10450 21734 10460 21786
rect 10484 21734 10514 21786
rect 10514 21734 10526 21786
rect 10526 21734 10540 21786
rect 10564 21734 10578 21786
rect 10578 21734 10590 21786
rect 10590 21734 10620 21786
rect 10644 21734 10654 21786
rect 10654 21734 10700 21786
rect 10404 21732 10460 21734
rect 10484 21732 10540 21734
rect 10564 21732 10620 21734
rect 10644 21732 10700 21734
rect 10404 20698 10460 20700
rect 10484 20698 10540 20700
rect 10564 20698 10620 20700
rect 10644 20698 10700 20700
rect 10404 20646 10450 20698
rect 10450 20646 10460 20698
rect 10484 20646 10514 20698
rect 10514 20646 10526 20698
rect 10526 20646 10540 20698
rect 10564 20646 10578 20698
rect 10578 20646 10590 20698
rect 10590 20646 10620 20698
rect 10644 20646 10654 20698
rect 10654 20646 10700 20698
rect 10404 20644 10460 20646
rect 10484 20644 10540 20646
rect 10564 20644 10620 20646
rect 10644 20644 10700 20646
rect 10404 19610 10460 19612
rect 10484 19610 10540 19612
rect 10564 19610 10620 19612
rect 10644 19610 10700 19612
rect 10404 19558 10450 19610
rect 10450 19558 10460 19610
rect 10484 19558 10514 19610
rect 10514 19558 10526 19610
rect 10526 19558 10540 19610
rect 10564 19558 10578 19610
rect 10578 19558 10590 19610
rect 10590 19558 10620 19610
rect 10644 19558 10654 19610
rect 10654 19558 10700 19610
rect 10404 19556 10460 19558
rect 10484 19556 10540 19558
rect 10564 19556 10620 19558
rect 10644 19556 10700 19558
rect 10404 18522 10460 18524
rect 10484 18522 10540 18524
rect 10564 18522 10620 18524
rect 10644 18522 10700 18524
rect 10404 18470 10450 18522
rect 10450 18470 10460 18522
rect 10484 18470 10514 18522
rect 10514 18470 10526 18522
rect 10526 18470 10540 18522
rect 10564 18470 10578 18522
rect 10578 18470 10590 18522
rect 10590 18470 10620 18522
rect 10644 18470 10654 18522
rect 10654 18470 10700 18522
rect 10404 18468 10460 18470
rect 10484 18468 10540 18470
rect 10564 18468 10620 18470
rect 10644 18468 10700 18470
rect 10404 17434 10460 17436
rect 10484 17434 10540 17436
rect 10564 17434 10620 17436
rect 10644 17434 10700 17436
rect 10404 17382 10450 17434
rect 10450 17382 10460 17434
rect 10484 17382 10514 17434
rect 10514 17382 10526 17434
rect 10526 17382 10540 17434
rect 10564 17382 10578 17434
rect 10578 17382 10590 17434
rect 10590 17382 10620 17434
rect 10644 17382 10654 17434
rect 10654 17382 10700 17434
rect 10404 17380 10460 17382
rect 10484 17380 10540 17382
rect 10564 17380 10620 17382
rect 10644 17380 10700 17382
rect 10404 16346 10460 16348
rect 10484 16346 10540 16348
rect 10564 16346 10620 16348
rect 10644 16346 10700 16348
rect 10404 16294 10450 16346
rect 10450 16294 10460 16346
rect 10484 16294 10514 16346
rect 10514 16294 10526 16346
rect 10526 16294 10540 16346
rect 10564 16294 10578 16346
rect 10578 16294 10590 16346
rect 10590 16294 10620 16346
rect 10644 16294 10654 16346
rect 10654 16294 10700 16346
rect 10404 16292 10460 16294
rect 10484 16292 10540 16294
rect 10564 16292 10620 16294
rect 10644 16292 10700 16294
rect 10404 15258 10460 15260
rect 10484 15258 10540 15260
rect 10564 15258 10620 15260
rect 10644 15258 10700 15260
rect 10404 15206 10450 15258
rect 10450 15206 10460 15258
rect 10484 15206 10514 15258
rect 10514 15206 10526 15258
rect 10526 15206 10540 15258
rect 10564 15206 10578 15258
rect 10578 15206 10590 15258
rect 10590 15206 10620 15258
rect 10644 15206 10654 15258
rect 10654 15206 10700 15258
rect 10404 15204 10460 15206
rect 10484 15204 10540 15206
rect 10564 15204 10620 15206
rect 10644 15204 10700 15206
rect 10404 14170 10460 14172
rect 10484 14170 10540 14172
rect 10564 14170 10620 14172
rect 10644 14170 10700 14172
rect 10404 14118 10450 14170
rect 10450 14118 10460 14170
rect 10484 14118 10514 14170
rect 10514 14118 10526 14170
rect 10526 14118 10540 14170
rect 10564 14118 10578 14170
rect 10578 14118 10590 14170
rect 10590 14118 10620 14170
rect 10644 14118 10654 14170
rect 10654 14118 10700 14170
rect 10404 14116 10460 14118
rect 10484 14116 10540 14118
rect 10564 14116 10620 14118
rect 10644 14116 10700 14118
rect 10404 13082 10460 13084
rect 10484 13082 10540 13084
rect 10564 13082 10620 13084
rect 10644 13082 10700 13084
rect 10404 13030 10450 13082
rect 10450 13030 10460 13082
rect 10484 13030 10514 13082
rect 10514 13030 10526 13082
rect 10526 13030 10540 13082
rect 10564 13030 10578 13082
rect 10578 13030 10590 13082
rect 10590 13030 10620 13082
rect 10644 13030 10654 13082
rect 10654 13030 10700 13082
rect 10404 13028 10460 13030
rect 10484 13028 10540 13030
rect 10564 13028 10620 13030
rect 10644 13028 10700 13030
rect 10404 11994 10460 11996
rect 10484 11994 10540 11996
rect 10564 11994 10620 11996
rect 10644 11994 10700 11996
rect 10404 11942 10450 11994
rect 10450 11942 10460 11994
rect 10484 11942 10514 11994
rect 10514 11942 10526 11994
rect 10526 11942 10540 11994
rect 10564 11942 10578 11994
rect 10578 11942 10590 11994
rect 10590 11942 10620 11994
rect 10644 11942 10654 11994
rect 10654 11942 10700 11994
rect 10404 11940 10460 11942
rect 10484 11940 10540 11942
rect 10564 11940 10620 11942
rect 10644 11940 10700 11942
rect 10404 10906 10460 10908
rect 10484 10906 10540 10908
rect 10564 10906 10620 10908
rect 10644 10906 10700 10908
rect 10404 10854 10450 10906
rect 10450 10854 10460 10906
rect 10484 10854 10514 10906
rect 10514 10854 10526 10906
rect 10526 10854 10540 10906
rect 10564 10854 10578 10906
rect 10578 10854 10590 10906
rect 10590 10854 10620 10906
rect 10644 10854 10654 10906
rect 10654 10854 10700 10906
rect 10404 10852 10460 10854
rect 10484 10852 10540 10854
rect 10564 10852 10620 10854
rect 10644 10852 10700 10854
rect 10404 9818 10460 9820
rect 10484 9818 10540 9820
rect 10564 9818 10620 9820
rect 10644 9818 10700 9820
rect 10404 9766 10450 9818
rect 10450 9766 10460 9818
rect 10484 9766 10514 9818
rect 10514 9766 10526 9818
rect 10526 9766 10540 9818
rect 10564 9766 10578 9818
rect 10578 9766 10590 9818
rect 10590 9766 10620 9818
rect 10644 9766 10654 9818
rect 10654 9766 10700 9818
rect 10404 9764 10460 9766
rect 10484 9764 10540 9766
rect 10564 9764 10620 9766
rect 10644 9764 10700 9766
rect 10404 8730 10460 8732
rect 10484 8730 10540 8732
rect 10564 8730 10620 8732
rect 10644 8730 10700 8732
rect 10404 8678 10450 8730
rect 10450 8678 10460 8730
rect 10484 8678 10514 8730
rect 10514 8678 10526 8730
rect 10526 8678 10540 8730
rect 10564 8678 10578 8730
rect 10578 8678 10590 8730
rect 10590 8678 10620 8730
rect 10644 8678 10654 8730
rect 10654 8678 10700 8730
rect 10404 8676 10460 8678
rect 10484 8676 10540 8678
rect 10564 8676 10620 8678
rect 10644 8676 10700 8678
rect 10404 7642 10460 7644
rect 10484 7642 10540 7644
rect 10564 7642 10620 7644
rect 10644 7642 10700 7644
rect 10404 7590 10450 7642
rect 10450 7590 10460 7642
rect 10484 7590 10514 7642
rect 10514 7590 10526 7642
rect 10526 7590 10540 7642
rect 10564 7590 10578 7642
rect 10578 7590 10590 7642
rect 10590 7590 10620 7642
rect 10644 7590 10654 7642
rect 10654 7590 10700 7642
rect 10404 7588 10460 7590
rect 10484 7588 10540 7590
rect 10564 7588 10620 7590
rect 10644 7588 10700 7590
rect 10404 6554 10460 6556
rect 10484 6554 10540 6556
rect 10564 6554 10620 6556
rect 10644 6554 10700 6556
rect 10404 6502 10450 6554
rect 10450 6502 10460 6554
rect 10484 6502 10514 6554
rect 10514 6502 10526 6554
rect 10526 6502 10540 6554
rect 10564 6502 10578 6554
rect 10578 6502 10590 6554
rect 10590 6502 10620 6554
rect 10644 6502 10654 6554
rect 10654 6502 10700 6554
rect 10404 6500 10460 6502
rect 10484 6500 10540 6502
rect 10564 6500 10620 6502
rect 10644 6500 10700 6502
rect 10404 5466 10460 5468
rect 10484 5466 10540 5468
rect 10564 5466 10620 5468
rect 10644 5466 10700 5468
rect 10404 5414 10450 5466
rect 10450 5414 10460 5466
rect 10484 5414 10514 5466
rect 10514 5414 10526 5466
rect 10526 5414 10540 5466
rect 10564 5414 10578 5466
rect 10578 5414 10590 5466
rect 10590 5414 10620 5466
rect 10644 5414 10654 5466
rect 10654 5414 10700 5466
rect 10404 5412 10460 5414
rect 10484 5412 10540 5414
rect 10564 5412 10620 5414
rect 10644 5412 10700 5414
rect 10404 4378 10460 4380
rect 10484 4378 10540 4380
rect 10564 4378 10620 4380
rect 10644 4378 10700 4380
rect 10404 4326 10450 4378
rect 10450 4326 10460 4378
rect 10484 4326 10514 4378
rect 10514 4326 10526 4378
rect 10526 4326 10540 4378
rect 10564 4326 10578 4378
rect 10578 4326 10590 4378
rect 10590 4326 10620 4378
rect 10644 4326 10654 4378
rect 10654 4326 10700 4378
rect 10404 4324 10460 4326
rect 10484 4324 10540 4326
rect 10564 4324 10620 4326
rect 10644 4324 10700 4326
rect 15128 33210 15184 33212
rect 15208 33210 15264 33212
rect 15288 33210 15344 33212
rect 15368 33210 15424 33212
rect 15128 33158 15174 33210
rect 15174 33158 15184 33210
rect 15208 33158 15238 33210
rect 15238 33158 15250 33210
rect 15250 33158 15264 33210
rect 15288 33158 15302 33210
rect 15302 33158 15314 33210
rect 15314 33158 15344 33210
rect 15368 33158 15378 33210
rect 15378 33158 15424 33210
rect 15128 33156 15184 33158
rect 15208 33156 15264 33158
rect 15288 33156 15344 33158
rect 15368 33156 15424 33158
rect 24576 33210 24632 33212
rect 24656 33210 24712 33212
rect 24736 33210 24792 33212
rect 24816 33210 24872 33212
rect 24576 33158 24622 33210
rect 24622 33158 24632 33210
rect 24656 33158 24686 33210
rect 24686 33158 24698 33210
rect 24698 33158 24712 33210
rect 24736 33158 24750 33210
rect 24750 33158 24762 33210
rect 24762 33158 24792 33210
rect 24816 33158 24826 33210
rect 24826 33158 24872 33210
rect 24576 33156 24632 33158
rect 24656 33156 24712 33158
rect 24736 33156 24792 33158
rect 24816 33156 24872 33158
rect 34024 33210 34080 33212
rect 34104 33210 34160 33212
rect 34184 33210 34240 33212
rect 34264 33210 34320 33212
rect 34024 33158 34070 33210
rect 34070 33158 34080 33210
rect 34104 33158 34134 33210
rect 34134 33158 34146 33210
rect 34146 33158 34160 33210
rect 34184 33158 34198 33210
rect 34198 33158 34210 33210
rect 34210 33158 34240 33210
rect 34264 33158 34274 33210
rect 34274 33158 34320 33210
rect 34024 33156 34080 33158
rect 34104 33156 34160 33158
rect 34184 33156 34240 33158
rect 34264 33156 34320 33158
rect 19852 32666 19908 32668
rect 19932 32666 19988 32668
rect 20012 32666 20068 32668
rect 20092 32666 20148 32668
rect 19852 32614 19898 32666
rect 19898 32614 19908 32666
rect 19932 32614 19962 32666
rect 19962 32614 19974 32666
rect 19974 32614 19988 32666
rect 20012 32614 20026 32666
rect 20026 32614 20038 32666
rect 20038 32614 20068 32666
rect 20092 32614 20102 32666
rect 20102 32614 20148 32666
rect 19852 32612 19908 32614
rect 19932 32612 19988 32614
rect 20012 32612 20068 32614
rect 20092 32612 20148 32614
rect 29300 32666 29356 32668
rect 29380 32666 29436 32668
rect 29460 32666 29516 32668
rect 29540 32666 29596 32668
rect 29300 32614 29346 32666
rect 29346 32614 29356 32666
rect 29380 32614 29410 32666
rect 29410 32614 29422 32666
rect 29422 32614 29436 32666
rect 29460 32614 29474 32666
rect 29474 32614 29486 32666
rect 29486 32614 29516 32666
rect 29540 32614 29550 32666
rect 29550 32614 29596 32666
rect 29300 32612 29356 32614
rect 29380 32612 29436 32614
rect 29460 32612 29516 32614
rect 29540 32612 29596 32614
rect 15128 32122 15184 32124
rect 15208 32122 15264 32124
rect 15288 32122 15344 32124
rect 15368 32122 15424 32124
rect 15128 32070 15174 32122
rect 15174 32070 15184 32122
rect 15208 32070 15238 32122
rect 15238 32070 15250 32122
rect 15250 32070 15264 32122
rect 15288 32070 15302 32122
rect 15302 32070 15314 32122
rect 15314 32070 15344 32122
rect 15368 32070 15378 32122
rect 15378 32070 15424 32122
rect 15128 32068 15184 32070
rect 15208 32068 15264 32070
rect 15288 32068 15344 32070
rect 15368 32068 15424 32070
rect 15128 31034 15184 31036
rect 15208 31034 15264 31036
rect 15288 31034 15344 31036
rect 15368 31034 15424 31036
rect 15128 30982 15174 31034
rect 15174 30982 15184 31034
rect 15208 30982 15238 31034
rect 15238 30982 15250 31034
rect 15250 30982 15264 31034
rect 15288 30982 15302 31034
rect 15302 30982 15314 31034
rect 15314 30982 15344 31034
rect 15368 30982 15378 31034
rect 15378 30982 15424 31034
rect 15128 30980 15184 30982
rect 15208 30980 15264 30982
rect 15288 30980 15344 30982
rect 15368 30980 15424 30982
rect 15128 29946 15184 29948
rect 15208 29946 15264 29948
rect 15288 29946 15344 29948
rect 15368 29946 15424 29948
rect 15128 29894 15174 29946
rect 15174 29894 15184 29946
rect 15208 29894 15238 29946
rect 15238 29894 15250 29946
rect 15250 29894 15264 29946
rect 15288 29894 15302 29946
rect 15302 29894 15314 29946
rect 15314 29894 15344 29946
rect 15368 29894 15378 29946
rect 15378 29894 15424 29946
rect 15128 29892 15184 29894
rect 15208 29892 15264 29894
rect 15288 29892 15344 29894
rect 15368 29892 15424 29894
rect 15128 28858 15184 28860
rect 15208 28858 15264 28860
rect 15288 28858 15344 28860
rect 15368 28858 15424 28860
rect 15128 28806 15174 28858
rect 15174 28806 15184 28858
rect 15208 28806 15238 28858
rect 15238 28806 15250 28858
rect 15250 28806 15264 28858
rect 15288 28806 15302 28858
rect 15302 28806 15314 28858
rect 15314 28806 15344 28858
rect 15368 28806 15378 28858
rect 15378 28806 15424 28858
rect 15128 28804 15184 28806
rect 15208 28804 15264 28806
rect 15288 28804 15344 28806
rect 15368 28804 15424 28806
rect 15128 27770 15184 27772
rect 15208 27770 15264 27772
rect 15288 27770 15344 27772
rect 15368 27770 15424 27772
rect 15128 27718 15174 27770
rect 15174 27718 15184 27770
rect 15208 27718 15238 27770
rect 15238 27718 15250 27770
rect 15250 27718 15264 27770
rect 15288 27718 15302 27770
rect 15302 27718 15314 27770
rect 15314 27718 15344 27770
rect 15368 27718 15378 27770
rect 15378 27718 15424 27770
rect 15128 27716 15184 27718
rect 15208 27716 15264 27718
rect 15288 27716 15344 27718
rect 15368 27716 15424 27718
rect 15128 26682 15184 26684
rect 15208 26682 15264 26684
rect 15288 26682 15344 26684
rect 15368 26682 15424 26684
rect 15128 26630 15174 26682
rect 15174 26630 15184 26682
rect 15208 26630 15238 26682
rect 15238 26630 15250 26682
rect 15250 26630 15264 26682
rect 15288 26630 15302 26682
rect 15302 26630 15314 26682
rect 15314 26630 15344 26682
rect 15368 26630 15378 26682
rect 15378 26630 15424 26682
rect 15128 26628 15184 26630
rect 15208 26628 15264 26630
rect 15288 26628 15344 26630
rect 15368 26628 15424 26630
rect 15128 25594 15184 25596
rect 15208 25594 15264 25596
rect 15288 25594 15344 25596
rect 15368 25594 15424 25596
rect 15128 25542 15174 25594
rect 15174 25542 15184 25594
rect 15208 25542 15238 25594
rect 15238 25542 15250 25594
rect 15250 25542 15264 25594
rect 15288 25542 15302 25594
rect 15302 25542 15314 25594
rect 15314 25542 15344 25594
rect 15368 25542 15378 25594
rect 15378 25542 15424 25594
rect 15128 25540 15184 25542
rect 15208 25540 15264 25542
rect 15288 25540 15344 25542
rect 15368 25540 15424 25542
rect 15128 24506 15184 24508
rect 15208 24506 15264 24508
rect 15288 24506 15344 24508
rect 15368 24506 15424 24508
rect 15128 24454 15174 24506
rect 15174 24454 15184 24506
rect 15208 24454 15238 24506
rect 15238 24454 15250 24506
rect 15250 24454 15264 24506
rect 15288 24454 15302 24506
rect 15302 24454 15314 24506
rect 15314 24454 15344 24506
rect 15368 24454 15378 24506
rect 15378 24454 15424 24506
rect 15128 24452 15184 24454
rect 15208 24452 15264 24454
rect 15288 24452 15344 24454
rect 15368 24452 15424 24454
rect 15128 23418 15184 23420
rect 15208 23418 15264 23420
rect 15288 23418 15344 23420
rect 15368 23418 15424 23420
rect 15128 23366 15174 23418
rect 15174 23366 15184 23418
rect 15208 23366 15238 23418
rect 15238 23366 15250 23418
rect 15250 23366 15264 23418
rect 15288 23366 15302 23418
rect 15302 23366 15314 23418
rect 15314 23366 15344 23418
rect 15368 23366 15378 23418
rect 15378 23366 15424 23418
rect 15128 23364 15184 23366
rect 15208 23364 15264 23366
rect 15288 23364 15344 23366
rect 15368 23364 15424 23366
rect 15128 22330 15184 22332
rect 15208 22330 15264 22332
rect 15288 22330 15344 22332
rect 15368 22330 15424 22332
rect 15128 22278 15174 22330
rect 15174 22278 15184 22330
rect 15208 22278 15238 22330
rect 15238 22278 15250 22330
rect 15250 22278 15264 22330
rect 15288 22278 15302 22330
rect 15302 22278 15314 22330
rect 15314 22278 15344 22330
rect 15368 22278 15378 22330
rect 15378 22278 15424 22330
rect 15128 22276 15184 22278
rect 15208 22276 15264 22278
rect 15288 22276 15344 22278
rect 15368 22276 15424 22278
rect 15128 21242 15184 21244
rect 15208 21242 15264 21244
rect 15288 21242 15344 21244
rect 15368 21242 15424 21244
rect 15128 21190 15174 21242
rect 15174 21190 15184 21242
rect 15208 21190 15238 21242
rect 15238 21190 15250 21242
rect 15250 21190 15264 21242
rect 15288 21190 15302 21242
rect 15302 21190 15314 21242
rect 15314 21190 15344 21242
rect 15368 21190 15378 21242
rect 15378 21190 15424 21242
rect 15128 21188 15184 21190
rect 15208 21188 15264 21190
rect 15288 21188 15344 21190
rect 15368 21188 15424 21190
rect 15128 20154 15184 20156
rect 15208 20154 15264 20156
rect 15288 20154 15344 20156
rect 15368 20154 15424 20156
rect 15128 20102 15174 20154
rect 15174 20102 15184 20154
rect 15208 20102 15238 20154
rect 15238 20102 15250 20154
rect 15250 20102 15264 20154
rect 15288 20102 15302 20154
rect 15302 20102 15314 20154
rect 15314 20102 15344 20154
rect 15368 20102 15378 20154
rect 15378 20102 15424 20154
rect 15128 20100 15184 20102
rect 15208 20100 15264 20102
rect 15288 20100 15344 20102
rect 15368 20100 15424 20102
rect 24576 32122 24632 32124
rect 24656 32122 24712 32124
rect 24736 32122 24792 32124
rect 24816 32122 24872 32124
rect 24576 32070 24622 32122
rect 24622 32070 24632 32122
rect 24656 32070 24686 32122
rect 24686 32070 24698 32122
rect 24698 32070 24712 32122
rect 24736 32070 24750 32122
rect 24750 32070 24762 32122
rect 24762 32070 24792 32122
rect 24816 32070 24826 32122
rect 24826 32070 24872 32122
rect 24576 32068 24632 32070
rect 24656 32068 24712 32070
rect 24736 32068 24792 32070
rect 24816 32068 24872 32070
rect 34024 32122 34080 32124
rect 34104 32122 34160 32124
rect 34184 32122 34240 32124
rect 34264 32122 34320 32124
rect 34024 32070 34070 32122
rect 34070 32070 34080 32122
rect 34104 32070 34134 32122
rect 34134 32070 34146 32122
rect 34146 32070 34160 32122
rect 34184 32070 34198 32122
rect 34198 32070 34210 32122
rect 34210 32070 34240 32122
rect 34264 32070 34274 32122
rect 34274 32070 34320 32122
rect 34024 32068 34080 32070
rect 34104 32068 34160 32070
rect 34184 32068 34240 32070
rect 34264 32068 34320 32070
rect 19852 31578 19908 31580
rect 19932 31578 19988 31580
rect 20012 31578 20068 31580
rect 20092 31578 20148 31580
rect 19852 31526 19898 31578
rect 19898 31526 19908 31578
rect 19932 31526 19962 31578
rect 19962 31526 19974 31578
rect 19974 31526 19988 31578
rect 20012 31526 20026 31578
rect 20026 31526 20038 31578
rect 20038 31526 20068 31578
rect 20092 31526 20102 31578
rect 20102 31526 20148 31578
rect 19852 31524 19908 31526
rect 19932 31524 19988 31526
rect 20012 31524 20068 31526
rect 20092 31524 20148 31526
rect 15128 19066 15184 19068
rect 15208 19066 15264 19068
rect 15288 19066 15344 19068
rect 15368 19066 15424 19068
rect 15128 19014 15174 19066
rect 15174 19014 15184 19066
rect 15208 19014 15238 19066
rect 15238 19014 15250 19066
rect 15250 19014 15264 19066
rect 15288 19014 15302 19066
rect 15302 19014 15314 19066
rect 15314 19014 15344 19066
rect 15368 19014 15378 19066
rect 15378 19014 15424 19066
rect 15128 19012 15184 19014
rect 15208 19012 15264 19014
rect 15288 19012 15344 19014
rect 15368 19012 15424 19014
rect 15128 17978 15184 17980
rect 15208 17978 15264 17980
rect 15288 17978 15344 17980
rect 15368 17978 15424 17980
rect 15128 17926 15174 17978
rect 15174 17926 15184 17978
rect 15208 17926 15238 17978
rect 15238 17926 15250 17978
rect 15250 17926 15264 17978
rect 15288 17926 15302 17978
rect 15302 17926 15314 17978
rect 15314 17926 15344 17978
rect 15368 17926 15378 17978
rect 15378 17926 15424 17978
rect 15128 17924 15184 17926
rect 15208 17924 15264 17926
rect 15288 17924 15344 17926
rect 15368 17924 15424 17926
rect 15128 16890 15184 16892
rect 15208 16890 15264 16892
rect 15288 16890 15344 16892
rect 15368 16890 15424 16892
rect 15128 16838 15174 16890
rect 15174 16838 15184 16890
rect 15208 16838 15238 16890
rect 15238 16838 15250 16890
rect 15250 16838 15264 16890
rect 15288 16838 15302 16890
rect 15302 16838 15314 16890
rect 15314 16838 15344 16890
rect 15368 16838 15378 16890
rect 15378 16838 15424 16890
rect 15128 16836 15184 16838
rect 15208 16836 15264 16838
rect 15288 16836 15344 16838
rect 15368 16836 15424 16838
rect 15128 15802 15184 15804
rect 15208 15802 15264 15804
rect 15288 15802 15344 15804
rect 15368 15802 15424 15804
rect 15128 15750 15174 15802
rect 15174 15750 15184 15802
rect 15208 15750 15238 15802
rect 15238 15750 15250 15802
rect 15250 15750 15264 15802
rect 15288 15750 15302 15802
rect 15302 15750 15314 15802
rect 15314 15750 15344 15802
rect 15368 15750 15378 15802
rect 15378 15750 15424 15802
rect 15128 15748 15184 15750
rect 15208 15748 15264 15750
rect 15288 15748 15344 15750
rect 15368 15748 15424 15750
rect 15128 14714 15184 14716
rect 15208 14714 15264 14716
rect 15288 14714 15344 14716
rect 15368 14714 15424 14716
rect 15128 14662 15174 14714
rect 15174 14662 15184 14714
rect 15208 14662 15238 14714
rect 15238 14662 15250 14714
rect 15250 14662 15264 14714
rect 15288 14662 15302 14714
rect 15302 14662 15314 14714
rect 15314 14662 15344 14714
rect 15368 14662 15378 14714
rect 15378 14662 15424 14714
rect 15128 14660 15184 14662
rect 15208 14660 15264 14662
rect 15288 14660 15344 14662
rect 15368 14660 15424 14662
rect 19852 30490 19908 30492
rect 19932 30490 19988 30492
rect 20012 30490 20068 30492
rect 20092 30490 20148 30492
rect 19852 30438 19898 30490
rect 19898 30438 19908 30490
rect 19932 30438 19962 30490
rect 19962 30438 19974 30490
rect 19974 30438 19988 30490
rect 20012 30438 20026 30490
rect 20026 30438 20038 30490
rect 20038 30438 20068 30490
rect 20092 30438 20102 30490
rect 20102 30438 20148 30490
rect 19852 30436 19908 30438
rect 19932 30436 19988 30438
rect 20012 30436 20068 30438
rect 20092 30436 20148 30438
rect 19852 29402 19908 29404
rect 19932 29402 19988 29404
rect 20012 29402 20068 29404
rect 20092 29402 20148 29404
rect 19852 29350 19898 29402
rect 19898 29350 19908 29402
rect 19932 29350 19962 29402
rect 19962 29350 19974 29402
rect 19974 29350 19988 29402
rect 20012 29350 20026 29402
rect 20026 29350 20038 29402
rect 20038 29350 20068 29402
rect 20092 29350 20102 29402
rect 20102 29350 20148 29402
rect 19852 29348 19908 29350
rect 19932 29348 19988 29350
rect 20012 29348 20068 29350
rect 20092 29348 20148 29350
rect 19852 28314 19908 28316
rect 19932 28314 19988 28316
rect 20012 28314 20068 28316
rect 20092 28314 20148 28316
rect 19852 28262 19898 28314
rect 19898 28262 19908 28314
rect 19932 28262 19962 28314
rect 19962 28262 19974 28314
rect 19974 28262 19988 28314
rect 20012 28262 20026 28314
rect 20026 28262 20038 28314
rect 20038 28262 20068 28314
rect 20092 28262 20102 28314
rect 20102 28262 20148 28314
rect 19852 28260 19908 28262
rect 19932 28260 19988 28262
rect 20012 28260 20068 28262
rect 20092 28260 20148 28262
rect 19852 27226 19908 27228
rect 19932 27226 19988 27228
rect 20012 27226 20068 27228
rect 20092 27226 20148 27228
rect 19852 27174 19898 27226
rect 19898 27174 19908 27226
rect 19932 27174 19962 27226
rect 19962 27174 19974 27226
rect 19974 27174 19988 27226
rect 20012 27174 20026 27226
rect 20026 27174 20038 27226
rect 20038 27174 20068 27226
rect 20092 27174 20102 27226
rect 20102 27174 20148 27226
rect 19852 27172 19908 27174
rect 19932 27172 19988 27174
rect 20012 27172 20068 27174
rect 20092 27172 20148 27174
rect 19852 26138 19908 26140
rect 19932 26138 19988 26140
rect 20012 26138 20068 26140
rect 20092 26138 20148 26140
rect 19852 26086 19898 26138
rect 19898 26086 19908 26138
rect 19932 26086 19962 26138
rect 19962 26086 19974 26138
rect 19974 26086 19988 26138
rect 20012 26086 20026 26138
rect 20026 26086 20038 26138
rect 20038 26086 20068 26138
rect 20092 26086 20102 26138
rect 20102 26086 20148 26138
rect 19852 26084 19908 26086
rect 19932 26084 19988 26086
rect 20012 26084 20068 26086
rect 20092 26084 20148 26086
rect 15128 13626 15184 13628
rect 15208 13626 15264 13628
rect 15288 13626 15344 13628
rect 15368 13626 15424 13628
rect 15128 13574 15174 13626
rect 15174 13574 15184 13626
rect 15208 13574 15238 13626
rect 15238 13574 15250 13626
rect 15250 13574 15264 13626
rect 15288 13574 15302 13626
rect 15302 13574 15314 13626
rect 15314 13574 15344 13626
rect 15368 13574 15378 13626
rect 15378 13574 15424 13626
rect 15128 13572 15184 13574
rect 15208 13572 15264 13574
rect 15288 13572 15344 13574
rect 15368 13572 15424 13574
rect 15128 12538 15184 12540
rect 15208 12538 15264 12540
rect 15288 12538 15344 12540
rect 15368 12538 15424 12540
rect 15128 12486 15174 12538
rect 15174 12486 15184 12538
rect 15208 12486 15238 12538
rect 15238 12486 15250 12538
rect 15250 12486 15264 12538
rect 15288 12486 15302 12538
rect 15302 12486 15314 12538
rect 15314 12486 15344 12538
rect 15368 12486 15378 12538
rect 15378 12486 15424 12538
rect 15128 12484 15184 12486
rect 15208 12484 15264 12486
rect 15288 12484 15344 12486
rect 15368 12484 15424 12486
rect 15128 11450 15184 11452
rect 15208 11450 15264 11452
rect 15288 11450 15344 11452
rect 15368 11450 15424 11452
rect 15128 11398 15174 11450
rect 15174 11398 15184 11450
rect 15208 11398 15238 11450
rect 15238 11398 15250 11450
rect 15250 11398 15264 11450
rect 15288 11398 15302 11450
rect 15302 11398 15314 11450
rect 15314 11398 15344 11450
rect 15368 11398 15378 11450
rect 15378 11398 15424 11450
rect 15128 11396 15184 11398
rect 15208 11396 15264 11398
rect 15288 11396 15344 11398
rect 15368 11396 15424 11398
rect 19852 25050 19908 25052
rect 19932 25050 19988 25052
rect 20012 25050 20068 25052
rect 20092 25050 20148 25052
rect 19852 24998 19898 25050
rect 19898 24998 19908 25050
rect 19932 24998 19962 25050
rect 19962 24998 19974 25050
rect 19974 24998 19988 25050
rect 20012 24998 20026 25050
rect 20026 24998 20038 25050
rect 20038 24998 20068 25050
rect 20092 24998 20102 25050
rect 20102 24998 20148 25050
rect 19852 24996 19908 24998
rect 19932 24996 19988 24998
rect 20012 24996 20068 24998
rect 20092 24996 20148 24998
rect 19852 23962 19908 23964
rect 19932 23962 19988 23964
rect 20012 23962 20068 23964
rect 20092 23962 20148 23964
rect 19852 23910 19898 23962
rect 19898 23910 19908 23962
rect 19932 23910 19962 23962
rect 19962 23910 19974 23962
rect 19974 23910 19988 23962
rect 20012 23910 20026 23962
rect 20026 23910 20038 23962
rect 20038 23910 20068 23962
rect 20092 23910 20102 23962
rect 20102 23910 20148 23962
rect 19852 23908 19908 23910
rect 19932 23908 19988 23910
rect 20012 23908 20068 23910
rect 20092 23908 20148 23910
rect 19852 22874 19908 22876
rect 19932 22874 19988 22876
rect 20012 22874 20068 22876
rect 20092 22874 20148 22876
rect 19852 22822 19898 22874
rect 19898 22822 19908 22874
rect 19932 22822 19962 22874
rect 19962 22822 19974 22874
rect 19974 22822 19988 22874
rect 20012 22822 20026 22874
rect 20026 22822 20038 22874
rect 20038 22822 20068 22874
rect 20092 22822 20102 22874
rect 20102 22822 20148 22874
rect 19852 22820 19908 22822
rect 19932 22820 19988 22822
rect 20012 22820 20068 22822
rect 20092 22820 20148 22822
rect 19852 21786 19908 21788
rect 19932 21786 19988 21788
rect 20012 21786 20068 21788
rect 20092 21786 20148 21788
rect 19852 21734 19898 21786
rect 19898 21734 19908 21786
rect 19932 21734 19962 21786
rect 19962 21734 19974 21786
rect 19974 21734 19988 21786
rect 20012 21734 20026 21786
rect 20026 21734 20038 21786
rect 20038 21734 20068 21786
rect 20092 21734 20102 21786
rect 20102 21734 20148 21786
rect 19852 21732 19908 21734
rect 19932 21732 19988 21734
rect 20012 21732 20068 21734
rect 20092 21732 20148 21734
rect 19852 20698 19908 20700
rect 19932 20698 19988 20700
rect 20012 20698 20068 20700
rect 20092 20698 20148 20700
rect 19852 20646 19898 20698
rect 19898 20646 19908 20698
rect 19932 20646 19962 20698
rect 19962 20646 19974 20698
rect 19974 20646 19988 20698
rect 20012 20646 20026 20698
rect 20026 20646 20038 20698
rect 20038 20646 20068 20698
rect 20092 20646 20102 20698
rect 20102 20646 20148 20698
rect 19852 20644 19908 20646
rect 19932 20644 19988 20646
rect 20012 20644 20068 20646
rect 20092 20644 20148 20646
rect 24576 31034 24632 31036
rect 24656 31034 24712 31036
rect 24736 31034 24792 31036
rect 24816 31034 24872 31036
rect 24576 30982 24622 31034
rect 24622 30982 24632 31034
rect 24656 30982 24686 31034
rect 24686 30982 24698 31034
rect 24698 30982 24712 31034
rect 24736 30982 24750 31034
rect 24750 30982 24762 31034
rect 24762 30982 24792 31034
rect 24816 30982 24826 31034
rect 24826 30982 24872 31034
rect 24576 30980 24632 30982
rect 24656 30980 24712 30982
rect 24736 30980 24792 30982
rect 24816 30980 24872 30982
rect 19852 19610 19908 19612
rect 19932 19610 19988 19612
rect 20012 19610 20068 19612
rect 20092 19610 20148 19612
rect 19852 19558 19898 19610
rect 19898 19558 19908 19610
rect 19932 19558 19962 19610
rect 19962 19558 19974 19610
rect 19974 19558 19988 19610
rect 20012 19558 20026 19610
rect 20026 19558 20038 19610
rect 20038 19558 20068 19610
rect 20092 19558 20102 19610
rect 20102 19558 20148 19610
rect 19852 19556 19908 19558
rect 19932 19556 19988 19558
rect 20012 19556 20068 19558
rect 20092 19556 20148 19558
rect 19852 18522 19908 18524
rect 19932 18522 19988 18524
rect 20012 18522 20068 18524
rect 20092 18522 20148 18524
rect 19852 18470 19898 18522
rect 19898 18470 19908 18522
rect 19932 18470 19962 18522
rect 19962 18470 19974 18522
rect 19974 18470 19988 18522
rect 20012 18470 20026 18522
rect 20026 18470 20038 18522
rect 20038 18470 20068 18522
rect 20092 18470 20102 18522
rect 20102 18470 20148 18522
rect 19852 18468 19908 18470
rect 19932 18468 19988 18470
rect 20012 18468 20068 18470
rect 20092 18468 20148 18470
rect 19852 17434 19908 17436
rect 19932 17434 19988 17436
rect 20012 17434 20068 17436
rect 20092 17434 20148 17436
rect 19852 17382 19898 17434
rect 19898 17382 19908 17434
rect 19932 17382 19962 17434
rect 19962 17382 19974 17434
rect 19974 17382 19988 17434
rect 20012 17382 20026 17434
rect 20026 17382 20038 17434
rect 20038 17382 20068 17434
rect 20092 17382 20102 17434
rect 20102 17382 20148 17434
rect 19852 17380 19908 17382
rect 19932 17380 19988 17382
rect 20012 17380 20068 17382
rect 20092 17380 20148 17382
rect 15128 10362 15184 10364
rect 15208 10362 15264 10364
rect 15288 10362 15344 10364
rect 15368 10362 15424 10364
rect 15128 10310 15174 10362
rect 15174 10310 15184 10362
rect 15208 10310 15238 10362
rect 15238 10310 15250 10362
rect 15250 10310 15264 10362
rect 15288 10310 15302 10362
rect 15302 10310 15314 10362
rect 15314 10310 15344 10362
rect 15368 10310 15378 10362
rect 15378 10310 15424 10362
rect 15128 10308 15184 10310
rect 15208 10308 15264 10310
rect 15288 10308 15344 10310
rect 15368 10308 15424 10310
rect 19852 16346 19908 16348
rect 19932 16346 19988 16348
rect 20012 16346 20068 16348
rect 20092 16346 20148 16348
rect 19852 16294 19898 16346
rect 19898 16294 19908 16346
rect 19932 16294 19962 16346
rect 19962 16294 19974 16346
rect 19974 16294 19988 16346
rect 20012 16294 20026 16346
rect 20026 16294 20038 16346
rect 20038 16294 20068 16346
rect 20092 16294 20102 16346
rect 20102 16294 20148 16346
rect 19852 16292 19908 16294
rect 19932 16292 19988 16294
rect 20012 16292 20068 16294
rect 20092 16292 20148 16294
rect 19852 15258 19908 15260
rect 19932 15258 19988 15260
rect 20012 15258 20068 15260
rect 20092 15258 20148 15260
rect 19852 15206 19898 15258
rect 19898 15206 19908 15258
rect 19932 15206 19962 15258
rect 19962 15206 19974 15258
rect 19974 15206 19988 15258
rect 20012 15206 20026 15258
rect 20026 15206 20038 15258
rect 20038 15206 20068 15258
rect 20092 15206 20102 15258
rect 20102 15206 20148 15258
rect 19852 15204 19908 15206
rect 19932 15204 19988 15206
rect 20012 15204 20068 15206
rect 20092 15204 20148 15206
rect 19852 14170 19908 14172
rect 19932 14170 19988 14172
rect 20012 14170 20068 14172
rect 20092 14170 20148 14172
rect 19852 14118 19898 14170
rect 19898 14118 19908 14170
rect 19932 14118 19962 14170
rect 19962 14118 19974 14170
rect 19974 14118 19988 14170
rect 20012 14118 20026 14170
rect 20026 14118 20038 14170
rect 20038 14118 20068 14170
rect 20092 14118 20102 14170
rect 20102 14118 20148 14170
rect 19852 14116 19908 14118
rect 19932 14116 19988 14118
rect 20012 14116 20068 14118
rect 20092 14116 20148 14118
rect 19852 13082 19908 13084
rect 19932 13082 19988 13084
rect 20012 13082 20068 13084
rect 20092 13082 20148 13084
rect 19852 13030 19898 13082
rect 19898 13030 19908 13082
rect 19932 13030 19962 13082
rect 19962 13030 19974 13082
rect 19974 13030 19988 13082
rect 20012 13030 20026 13082
rect 20026 13030 20038 13082
rect 20038 13030 20068 13082
rect 20092 13030 20102 13082
rect 20102 13030 20148 13082
rect 19852 13028 19908 13030
rect 19932 13028 19988 13030
rect 20012 13028 20068 13030
rect 20092 13028 20148 13030
rect 15128 9274 15184 9276
rect 15208 9274 15264 9276
rect 15288 9274 15344 9276
rect 15368 9274 15424 9276
rect 15128 9222 15174 9274
rect 15174 9222 15184 9274
rect 15208 9222 15238 9274
rect 15238 9222 15250 9274
rect 15250 9222 15264 9274
rect 15288 9222 15302 9274
rect 15302 9222 15314 9274
rect 15314 9222 15344 9274
rect 15368 9222 15378 9274
rect 15378 9222 15424 9274
rect 15128 9220 15184 9222
rect 15208 9220 15264 9222
rect 15288 9220 15344 9222
rect 15368 9220 15424 9222
rect 15128 8186 15184 8188
rect 15208 8186 15264 8188
rect 15288 8186 15344 8188
rect 15368 8186 15424 8188
rect 15128 8134 15174 8186
rect 15174 8134 15184 8186
rect 15208 8134 15238 8186
rect 15238 8134 15250 8186
rect 15250 8134 15264 8186
rect 15288 8134 15302 8186
rect 15302 8134 15314 8186
rect 15314 8134 15344 8186
rect 15368 8134 15378 8186
rect 15378 8134 15424 8186
rect 15128 8132 15184 8134
rect 15208 8132 15264 8134
rect 15288 8132 15344 8134
rect 15368 8132 15424 8134
rect 15128 7098 15184 7100
rect 15208 7098 15264 7100
rect 15288 7098 15344 7100
rect 15368 7098 15424 7100
rect 15128 7046 15174 7098
rect 15174 7046 15184 7098
rect 15208 7046 15238 7098
rect 15238 7046 15250 7098
rect 15250 7046 15264 7098
rect 15288 7046 15302 7098
rect 15302 7046 15314 7098
rect 15314 7046 15344 7098
rect 15368 7046 15378 7098
rect 15378 7046 15424 7098
rect 15128 7044 15184 7046
rect 15208 7044 15264 7046
rect 15288 7044 15344 7046
rect 15368 7044 15424 7046
rect 15128 6010 15184 6012
rect 15208 6010 15264 6012
rect 15288 6010 15344 6012
rect 15368 6010 15424 6012
rect 15128 5958 15174 6010
rect 15174 5958 15184 6010
rect 15208 5958 15238 6010
rect 15238 5958 15250 6010
rect 15250 5958 15264 6010
rect 15288 5958 15302 6010
rect 15302 5958 15314 6010
rect 15314 5958 15344 6010
rect 15368 5958 15378 6010
rect 15378 5958 15424 6010
rect 15128 5956 15184 5958
rect 15208 5956 15264 5958
rect 15288 5956 15344 5958
rect 15368 5956 15424 5958
rect 15128 4922 15184 4924
rect 15208 4922 15264 4924
rect 15288 4922 15344 4924
rect 15368 4922 15424 4924
rect 15128 4870 15174 4922
rect 15174 4870 15184 4922
rect 15208 4870 15238 4922
rect 15238 4870 15250 4922
rect 15250 4870 15264 4922
rect 15288 4870 15302 4922
rect 15302 4870 15314 4922
rect 15314 4870 15344 4922
rect 15368 4870 15378 4922
rect 15378 4870 15424 4922
rect 15128 4868 15184 4870
rect 15208 4868 15264 4870
rect 15288 4868 15344 4870
rect 15368 4868 15424 4870
rect 10404 3290 10460 3292
rect 10484 3290 10540 3292
rect 10564 3290 10620 3292
rect 10644 3290 10700 3292
rect 10404 3238 10450 3290
rect 10450 3238 10460 3290
rect 10484 3238 10514 3290
rect 10514 3238 10526 3290
rect 10526 3238 10540 3290
rect 10564 3238 10578 3290
rect 10578 3238 10590 3290
rect 10590 3238 10620 3290
rect 10644 3238 10654 3290
rect 10654 3238 10700 3290
rect 10404 3236 10460 3238
rect 10484 3236 10540 3238
rect 10564 3236 10620 3238
rect 10644 3236 10700 3238
rect 15128 3834 15184 3836
rect 15208 3834 15264 3836
rect 15288 3834 15344 3836
rect 15368 3834 15424 3836
rect 15128 3782 15174 3834
rect 15174 3782 15184 3834
rect 15208 3782 15238 3834
rect 15238 3782 15250 3834
rect 15250 3782 15264 3834
rect 15288 3782 15302 3834
rect 15302 3782 15314 3834
rect 15314 3782 15344 3834
rect 15368 3782 15378 3834
rect 15378 3782 15424 3834
rect 15128 3780 15184 3782
rect 15208 3780 15264 3782
rect 15288 3780 15344 3782
rect 15368 3780 15424 3782
rect 15128 2746 15184 2748
rect 15208 2746 15264 2748
rect 15288 2746 15344 2748
rect 15368 2746 15424 2748
rect 15128 2694 15174 2746
rect 15174 2694 15184 2746
rect 15208 2694 15238 2746
rect 15238 2694 15250 2746
rect 15250 2694 15264 2746
rect 15288 2694 15302 2746
rect 15302 2694 15314 2746
rect 15314 2694 15344 2746
rect 15368 2694 15378 2746
rect 15378 2694 15424 2746
rect 15128 2692 15184 2694
rect 15208 2692 15264 2694
rect 15288 2692 15344 2694
rect 15368 2692 15424 2694
rect 19852 11994 19908 11996
rect 19932 11994 19988 11996
rect 20012 11994 20068 11996
rect 20092 11994 20148 11996
rect 19852 11942 19898 11994
rect 19898 11942 19908 11994
rect 19932 11942 19962 11994
rect 19962 11942 19974 11994
rect 19974 11942 19988 11994
rect 20012 11942 20026 11994
rect 20026 11942 20038 11994
rect 20038 11942 20068 11994
rect 20092 11942 20102 11994
rect 20102 11942 20148 11994
rect 19852 11940 19908 11942
rect 19932 11940 19988 11942
rect 20012 11940 20068 11942
rect 20092 11940 20148 11942
rect 19852 10906 19908 10908
rect 19932 10906 19988 10908
rect 20012 10906 20068 10908
rect 20092 10906 20148 10908
rect 19852 10854 19898 10906
rect 19898 10854 19908 10906
rect 19932 10854 19962 10906
rect 19962 10854 19974 10906
rect 19974 10854 19988 10906
rect 20012 10854 20026 10906
rect 20026 10854 20038 10906
rect 20038 10854 20068 10906
rect 20092 10854 20102 10906
rect 20102 10854 20148 10906
rect 19852 10852 19908 10854
rect 19932 10852 19988 10854
rect 20012 10852 20068 10854
rect 20092 10852 20148 10854
rect 24576 29946 24632 29948
rect 24656 29946 24712 29948
rect 24736 29946 24792 29948
rect 24816 29946 24872 29948
rect 24576 29894 24622 29946
rect 24622 29894 24632 29946
rect 24656 29894 24686 29946
rect 24686 29894 24698 29946
rect 24698 29894 24712 29946
rect 24736 29894 24750 29946
rect 24750 29894 24762 29946
rect 24762 29894 24792 29946
rect 24816 29894 24826 29946
rect 24826 29894 24872 29946
rect 24576 29892 24632 29894
rect 24656 29892 24712 29894
rect 24736 29892 24792 29894
rect 24816 29892 24872 29894
rect 24576 28858 24632 28860
rect 24656 28858 24712 28860
rect 24736 28858 24792 28860
rect 24816 28858 24872 28860
rect 24576 28806 24622 28858
rect 24622 28806 24632 28858
rect 24656 28806 24686 28858
rect 24686 28806 24698 28858
rect 24698 28806 24712 28858
rect 24736 28806 24750 28858
rect 24750 28806 24762 28858
rect 24762 28806 24792 28858
rect 24816 28806 24826 28858
rect 24826 28806 24872 28858
rect 24576 28804 24632 28806
rect 24656 28804 24712 28806
rect 24736 28804 24792 28806
rect 24816 28804 24872 28806
rect 24576 27770 24632 27772
rect 24656 27770 24712 27772
rect 24736 27770 24792 27772
rect 24816 27770 24872 27772
rect 24576 27718 24622 27770
rect 24622 27718 24632 27770
rect 24656 27718 24686 27770
rect 24686 27718 24698 27770
rect 24698 27718 24712 27770
rect 24736 27718 24750 27770
rect 24750 27718 24762 27770
rect 24762 27718 24792 27770
rect 24816 27718 24826 27770
rect 24826 27718 24872 27770
rect 24576 27716 24632 27718
rect 24656 27716 24712 27718
rect 24736 27716 24792 27718
rect 24816 27716 24872 27718
rect 24576 26682 24632 26684
rect 24656 26682 24712 26684
rect 24736 26682 24792 26684
rect 24816 26682 24872 26684
rect 24576 26630 24622 26682
rect 24622 26630 24632 26682
rect 24656 26630 24686 26682
rect 24686 26630 24698 26682
rect 24698 26630 24712 26682
rect 24736 26630 24750 26682
rect 24750 26630 24762 26682
rect 24762 26630 24792 26682
rect 24816 26630 24826 26682
rect 24826 26630 24872 26682
rect 24576 26628 24632 26630
rect 24656 26628 24712 26630
rect 24736 26628 24792 26630
rect 24816 26628 24872 26630
rect 24576 25594 24632 25596
rect 24656 25594 24712 25596
rect 24736 25594 24792 25596
rect 24816 25594 24872 25596
rect 24576 25542 24622 25594
rect 24622 25542 24632 25594
rect 24656 25542 24686 25594
rect 24686 25542 24698 25594
rect 24698 25542 24712 25594
rect 24736 25542 24750 25594
rect 24750 25542 24762 25594
rect 24762 25542 24792 25594
rect 24816 25542 24826 25594
rect 24826 25542 24872 25594
rect 24576 25540 24632 25542
rect 24656 25540 24712 25542
rect 24736 25540 24792 25542
rect 24816 25540 24872 25542
rect 24576 24506 24632 24508
rect 24656 24506 24712 24508
rect 24736 24506 24792 24508
rect 24816 24506 24872 24508
rect 24576 24454 24622 24506
rect 24622 24454 24632 24506
rect 24656 24454 24686 24506
rect 24686 24454 24698 24506
rect 24698 24454 24712 24506
rect 24736 24454 24750 24506
rect 24750 24454 24762 24506
rect 24762 24454 24792 24506
rect 24816 24454 24826 24506
rect 24826 24454 24872 24506
rect 24576 24452 24632 24454
rect 24656 24452 24712 24454
rect 24736 24452 24792 24454
rect 24816 24452 24872 24454
rect 24576 23418 24632 23420
rect 24656 23418 24712 23420
rect 24736 23418 24792 23420
rect 24816 23418 24872 23420
rect 24576 23366 24622 23418
rect 24622 23366 24632 23418
rect 24656 23366 24686 23418
rect 24686 23366 24698 23418
rect 24698 23366 24712 23418
rect 24736 23366 24750 23418
rect 24750 23366 24762 23418
rect 24762 23366 24792 23418
rect 24816 23366 24826 23418
rect 24826 23366 24872 23418
rect 24576 23364 24632 23366
rect 24656 23364 24712 23366
rect 24736 23364 24792 23366
rect 24816 23364 24872 23366
rect 24576 22330 24632 22332
rect 24656 22330 24712 22332
rect 24736 22330 24792 22332
rect 24816 22330 24872 22332
rect 24576 22278 24622 22330
rect 24622 22278 24632 22330
rect 24656 22278 24686 22330
rect 24686 22278 24698 22330
rect 24698 22278 24712 22330
rect 24736 22278 24750 22330
rect 24750 22278 24762 22330
rect 24762 22278 24792 22330
rect 24816 22278 24826 22330
rect 24826 22278 24872 22330
rect 24576 22276 24632 22278
rect 24656 22276 24712 22278
rect 24736 22276 24792 22278
rect 24816 22276 24872 22278
rect 24576 21242 24632 21244
rect 24656 21242 24712 21244
rect 24736 21242 24792 21244
rect 24816 21242 24872 21244
rect 24576 21190 24622 21242
rect 24622 21190 24632 21242
rect 24656 21190 24686 21242
rect 24686 21190 24698 21242
rect 24698 21190 24712 21242
rect 24736 21190 24750 21242
rect 24750 21190 24762 21242
rect 24762 21190 24792 21242
rect 24816 21190 24826 21242
rect 24826 21190 24872 21242
rect 24576 21188 24632 21190
rect 24656 21188 24712 21190
rect 24736 21188 24792 21190
rect 24816 21188 24872 21190
rect 24576 20154 24632 20156
rect 24656 20154 24712 20156
rect 24736 20154 24792 20156
rect 24816 20154 24872 20156
rect 24576 20102 24622 20154
rect 24622 20102 24632 20154
rect 24656 20102 24686 20154
rect 24686 20102 24698 20154
rect 24698 20102 24712 20154
rect 24736 20102 24750 20154
rect 24750 20102 24762 20154
rect 24762 20102 24792 20154
rect 24816 20102 24826 20154
rect 24826 20102 24872 20154
rect 24576 20100 24632 20102
rect 24656 20100 24712 20102
rect 24736 20100 24792 20102
rect 24816 20100 24872 20102
rect 24576 19066 24632 19068
rect 24656 19066 24712 19068
rect 24736 19066 24792 19068
rect 24816 19066 24872 19068
rect 24576 19014 24622 19066
rect 24622 19014 24632 19066
rect 24656 19014 24686 19066
rect 24686 19014 24698 19066
rect 24698 19014 24712 19066
rect 24736 19014 24750 19066
rect 24750 19014 24762 19066
rect 24762 19014 24792 19066
rect 24816 19014 24826 19066
rect 24826 19014 24872 19066
rect 24576 19012 24632 19014
rect 24656 19012 24712 19014
rect 24736 19012 24792 19014
rect 24816 19012 24872 19014
rect 24576 17978 24632 17980
rect 24656 17978 24712 17980
rect 24736 17978 24792 17980
rect 24816 17978 24872 17980
rect 24576 17926 24622 17978
rect 24622 17926 24632 17978
rect 24656 17926 24686 17978
rect 24686 17926 24698 17978
rect 24698 17926 24712 17978
rect 24736 17926 24750 17978
rect 24750 17926 24762 17978
rect 24762 17926 24792 17978
rect 24816 17926 24826 17978
rect 24826 17926 24872 17978
rect 24576 17924 24632 17926
rect 24656 17924 24712 17926
rect 24736 17924 24792 17926
rect 24816 17924 24872 17926
rect 24576 16890 24632 16892
rect 24656 16890 24712 16892
rect 24736 16890 24792 16892
rect 24816 16890 24872 16892
rect 24576 16838 24622 16890
rect 24622 16838 24632 16890
rect 24656 16838 24686 16890
rect 24686 16838 24698 16890
rect 24698 16838 24712 16890
rect 24736 16838 24750 16890
rect 24750 16838 24762 16890
rect 24762 16838 24792 16890
rect 24816 16838 24826 16890
rect 24826 16838 24872 16890
rect 24576 16836 24632 16838
rect 24656 16836 24712 16838
rect 24736 16836 24792 16838
rect 24816 16836 24872 16838
rect 24576 15802 24632 15804
rect 24656 15802 24712 15804
rect 24736 15802 24792 15804
rect 24816 15802 24872 15804
rect 24576 15750 24622 15802
rect 24622 15750 24632 15802
rect 24656 15750 24686 15802
rect 24686 15750 24698 15802
rect 24698 15750 24712 15802
rect 24736 15750 24750 15802
rect 24750 15750 24762 15802
rect 24762 15750 24792 15802
rect 24816 15750 24826 15802
rect 24826 15750 24872 15802
rect 24576 15748 24632 15750
rect 24656 15748 24712 15750
rect 24736 15748 24792 15750
rect 24816 15748 24872 15750
rect 29300 31578 29356 31580
rect 29380 31578 29436 31580
rect 29460 31578 29516 31580
rect 29540 31578 29596 31580
rect 29300 31526 29346 31578
rect 29346 31526 29356 31578
rect 29380 31526 29410 31578
rect 29410 31526 29422 31578
rect 29422 31526 29436 31578
rect 29460 31526 29474 31578
rect 29474 31526 29486 31578
rect 29486 31526 29516 31578
rect 29540 31526 29550 31578
rect 29550 31526 29596 31578
rect 29300 31524 29356 31526
rect 29380 31524 29436 31526
rect 29460 31524 29516 31526
rect 29540 31524 29596 31526
rect 34024 31034 34080 31036
rect 34104 31034 34160 31036
rect 34184 31034 34240 31036
rect 34264 31034 34320 31036
rect 34024 30982 34070 31034
rect 34070 30982 34080 31034
rect 34104 30982 34134 31034
rect 34134 30982 34146 31034
rect 34146 30982 34160 31034
rect 34184 30982 34198 31034
rect 34198 30982 34210 31034
rect 34210 30982 34240 31034
rect 34264 30982 34274 31034
rect 34274 30982 34320 31034
rect 34024 30980 34080 30982
rect 34104 30980 34160 30982
rect 34184 30980 34240 30982
rect 34264 30980 34320 30982
rect 29300 30490 29356 30492
rect 29380 30490 29436 30492
rect 29460 30490 29516 30492
rect 29540 30490 29596 30492
rect 29300 30438 29346 30490
rect 29346 30438 29356 30490
rect 29380 30438 29410 30490
rect 29410 30438 29422 30490
rect 29422 30438 29436 30490
rect 29460 30438 29474 30490
rect 29474 30438 29486 30490
rect 29486 30438 29516 30490
rect 29540 30438 29550 30490
rect 29550 30438 29596 30490
rect 29300 30436 29356 30438
rect 29380 30436 29436 30438
rect 29460 30436 29516 30438
rect 29540 30436 29596 30438
rect 29300 29402 29356 29404
rect 29380 29402 29436 29404
rect 29460 29402 29516 29404
rect 29540 29402 29596 29404
rect 29300 29350 29346 29402
rect 29346 29350 29356 29402
rect 29380 29350 29410 29402
rect 29410 29350 29422 29402
rect 29422 29350 29436 29402
rect 29460 29350 29474 29402
rect 29474 29350 29486 29402
rect 29486 29350 29516 29402
rect 29540 29350 29550 29402
rect 29550 29350 29596 29402
rect 29300 29348 29356 29350
rect 29380 29348 29436 29350
rect 29460 29348 29516 29350
rect 29540 29348 29596 29350
rect 34024 29946 34080 29948
rect 34104 29946 34160 29948
rect 34184 29946 34240 29948
rect 34264 29946 34320 29948
rect 34024 29894 34070 29946
rect 34070 29894 34080 29946
rect 34104 29894 34134 29946
rect 34134 29894 34146 29946
rect 34146 29894 34160 29946
rect 34184 29894 34198 29946
rect 34198 29894 34210 29946
rect 34210 29894 34240 29946
rect 34264 29894 34274 29946
rect 34274 29894 34320 29946
rect 34024 29892 34080 29894
rect 34104 29892 34160 29894
rect 34184 29892 34240 29894
rect 34264 29892 34320 29894
rect 29300 28314 29356 28316
rect 29380 28314 29436 28316
rect 29460 28314 29516 28316
rect 29540 28314 29596 28316
rect 29300 28262 29346 28314
rect 29346 28262 29356 28314
rect 29380 28262 29410 28314
rect 29410 28262 29422 28314
rect 29422 28262 29436 28314
rect 29460 28262 29474 28314
rect 29474 28262 29486 28314
rect 29486 28262 29516 28314
rect 29540 28262 29550 28314
rect 29550 28262 29596 28314
rect 29300 28260 29356 28262
rect 29380 28260 29436 28262
rect 29460 28260 29516 28262
rect 29540 28260 29596 28262
rect 29300 27226 29356 27228
rect 29380 27226 29436 27228
rect 29460 27226 29516 27228
rect 29540 27226 29596 27228
rect 29300 27174 29346 27226
rect 29346 27174 29356 27226
rect 29380 27174 29410 27226
rect 29410 27174 29422 27226
rect 29422 27174 29436 27226
rect 29460 27174 29474 27226
rect 29474 27174 29486 27226
rect 29486 27174 29516 27226
rect 29540 27174 29550 27226
rect 29550 27174 29596 27226
rect 29300 27172 29356 27174
rect 29380 27172 29436 27174
rect 29460 27172 29516 27174
rect 29540 27172 29596 27174
rect 29300 26138 29356 26140
rect 29380 26138 29436 26140
rect 29460 26138 29516 26140
rect 29540 26138 29596 26140
rect 29300 26086 29346 26138
rect 29346 26086 29356 26138
rect 29380 26086 29410 26138
rect 29410 26086 29422 26138
rect 29422 26086 29436 26138
rect 29460 26086 29474 26138
rect 29474 26086 29486 26138
rect 29486 26086 29516 26138
rect 29540 26086 29550 26138
rect 29550 26086 29596 26138
rect 29300 26084 29356 26086
rect 29380 26084 29436 26086
rect 29460 26084 29516 26086
rect 29540 26084 29596 26086
rect 29300 25050 29356 25052
rect 29380 25050 29436 25052
rect 29460 25050 29516 25052
rect 29540 25050 29596 25052
rect 29300 24998 29346 25050
rect 29346 24998 29356 25050
rect 29380 24998 29410 25050
rect 29410 24998 29422 25050
rect 29422 24998 29436 25050
rect 29460 24998 29474 25050
rect 29474 24998 29486 25050
rect 29486 24998 29516 25050
rect 29540 24998 29550 25050
rect 29550 24998 29596 25050
rect 29300 24996 29356 24998
rect 29380 24996 29436 24998
rect 29460 24996 29516 24998
rect 29540 24996 29596 24998
rect 29300 23962 29356 23964
rect 29380 23962 29436 23964
rect 29460 23962 29516 23964
rect 29540 23962 29596 23964
rect 29300 23910 29346 23962
rect 29346 23910 29356 23962
rect 29380 23910 29410 23962
rect 29410 23910 29422 23962
rect 29422 23910 29436 23962
rect 29460 23910 29474 23962
rect 29474 23910 29486 23962
rect 29486 23910 29516 23962
rect 29540 23910 29550 23962
rect 29550 23910 29596 23962
rect 29300 23908 29356 23910
rect 29380 23908 29436 23910
rect 29460 23908 29516 23910
rect 29540 23908 29596 23910
rect 24576 14714 24632 14716
rect 24656 14714 24712 14716
rect 24736 14714 24792 14716
rect 24816 14714 24872 14716
rect 24576 14662 24622 14714
rect 24622 14662 24632 14714
rect 24656 14662 24686 14714
rect 24686 14662 24698 14714
rect 24698 14662 24712 14714
rect 24736 14662 24750 14714
rect 24750 14662 24762 14714
rect 24762 14662 24792 14714
rect 24816 14662 24826 14714
rect 24826 14662 24872 14714
rect 24576 14660 24632 14662
rect 24656 14660 24712 14662
rect 24736 14660 24792 14662
rect 24816 14660 24872 14662
rect 24576 13626 24632 13628
rect 24656 13626 24712 13628
rect 24736 13626 24792 13628
rect 24816 13626 24872 13628
rect 24576 13574 24622 13626
rect 24622 13574 24632 13626
rect 24656 13574 24686 13626
rect 24686 13574 24698 13626
rect 24698 13574 24712 13626
rect 24736 13574 24750 13626
rect 24750 13574 24762 13626
rect 24762 13574 24792 13626
rect 24816 13574 24826 13626
rect 24826 13574 24872 13626
rect 24576 13572 24632 13574
rect 24656 13572 24712 13574
rect 24736 13572 24792 13574
rect 24816 13572 24872 13574
rect 29300 22874 29356 22876
rect 29380 22874 29436 22876
rect 29460 22874 29516 22876
rect 29540 22874 29596 22876
rect 29300 22822 29346 22874
rect 29346 22822 29356 22874
rect 29380 22822 29410 22874
rect 29410 22822 29422 22874
rect 29422 22822 29436 22874
rect 29460 22822 29474 22874
rect 29474 22822 29486 22874
rect 29486 22822 29516 22874
rect 29540 22822 29550 22874
rect 29550 22822 29596 22874
rect 29300 22820 29356 22822
rect 29380 22820 29436 22822
rect 29460 22820 29516 22822
rect 29540 22820 29596 22822
rect 29300 21786 29356 21788
rect 29380 21786 29436 21788
rect 29460 21786 29516 21788
rect 29540 21786 29596 21788
rect 29300 21734 29346 21786
rect 29346 21734 29356 21786
rect 29380 21734 29410 21786
rect 29410 21734 29422 21786
rect 29422 21734 29436 21786
rect 29460 21734 29474 21786
rect 29474 21734 29486 21786
rect 29486 21734 29516 21786
rect 29540 21734 29550 21786
rect 29550 21734 29596 21786
rect 29300 21732 29356 21734
rect 29380 21732 29436 21734
rect 29460 21732 29516 21734
rect 29540 21732 29596 21734
rect 29300 20698 29356 20700
rect 29380 20698 29436 20700
rect 29460 20698 29516 20700
rect 29540 20698 29596 20700
rect 29300 20646 29346 20698
rect 29346 20646 29356 20698
rect 29380 20646 29410 20698
rect 29410 20646 29422 20698
rect 29422 20646 29436 20698
rect 29460 20646 29474 20698
rect 29474 20646 29486 20698
rect 29486 20646 29516 20698
rect 29540 20646 29550 20698
rect 29550 20646 29596 20698
rect 29300 20644 29356 20646
rect 29380 20644 29436 20646
rect 29460 20644 29516 20646
rect 29540 20644 29596 20646
rect 29300 19610 29356 19612
rect 29380 19610 29436 19612
rect 29460 19610 29516 19612
rect 29540 19610 29596 19612
rect 29300 19558 29346 19610
rect 29346 19558 29356 19610
rect 29380 19558 29410 19610
rect 29410 19558 29422 19610
rect 29422 19558 29436 19610
rect 29460 19558 29474 19610
rect 29474 19558 29486 19610
rect 29486 19558 29516 19610
rect 29540 19558 29550 19610
rect 29550 19558 29596 19610
rect 29300 19556 29356 19558
rect 29380 19556 29436 19558
rect 29460 19556 29516 19558
rect 29540 19556 29596 19558
rect 29300 18522 29356 18524
rect 29380 18522 29436 18524
rect 29460 18522 29516 18524
rect 29540 18522 29596 18524
rect 29300 18470 29346 18522
rect 29346 18470 29356 18522
rect 29380 18470 29410 18522
rect 29410 18470 29422 18522
rect 29422 18470 29436 18522
rect 29460 18470 29474 18522
rect 29474 18470 29486 18522
rect 29486 18470 29516 18522
rect 29540 18470 29550 18522
rect 29550 18470 29596 18522
rect 29300 18468 29356 18470
rect 29380 18468 29436 18470
rect 29460 18468 29516 18470
rect 29540 18468 29596 18470
rect 29300 17434 29356 17436
rect 29380 17434 29436 17436
rect 29460 17434 29516 17436
rect 29540 17434 29596 17436
rect 29300 17382 29346 17434
rect 29346 17382 29356 17434
rect 29380 17382 29410 17434
rect 29410 17382 29422 17434
rect 29422 17382 29436 17434
rect 29460 17382 29474 17434
rect 29474 17382 29486 17434
rect 29486 17382 29516 17434
rect 29540 17382 29550 17434
rect 29550 17382 29596 17434
rect 29300 17380 29356 17382
rect 29380 17380 29436 17382
rect 29460 17380 29516 17382
rect 29540 17380 29596 17382
rect 29300 16346 29356 16348
rect 29380 16346 29436 16348
rect 29460 16346 29516 16348
rect 29540 16346 29596 16348
rect 29300 16294 29346 16346
rect 29346 16294 29356 16346
rect 29380 16294 29410 16346
rect 29410 16294 29422 16346
rect 29422 16294 29436 16346
rect 29460 16294 29474 16346
rect 29474 16294 29486 16346
rect 29486 16294 29516 16346
rect 29540 16294 29550 16346
rect 29550 16294 29596 16346
rect 29300 16292 29356 16294
rect 29380 16292 29436 16294
rect 29460 16292 29516 16294
rect 29540 16292 29596 16294
rect 29300 15258 29356 15260
rect 29380 15258 29436 15260
rect 29460 15258 29516 15260
rect 29540 15258 29596 15260
rect 29300 15206 29346 15258
rect 29346 15206 29356 15258
rect 29380 15206 29410 15258
rect 29410 15206 29422 15258
rect 29422 15206 29436 15258
rect 29460 15206 29474 15258
rect 29474 15206 29486 15258
rect 29486 15206 29516 15258
rect 29540 15206 29550 15258
rect 29550 15206 29596 15258
rect 29300 15204 29356 15206
rect 29380 15204 29436 15206
rect 29460 15204 29516 15206
rect 29540 15204 29596 15206
rect 24576 12538 24632 12540
rect 24656 12538 24712 12540
rect 24736 12538 24792 12540
rect 24816 12538 24872 12540
rect 24576 12486 24622 12538
rect 24622 12486 24632 12538
rect 24656 12486 24686 12538
rect 24686 12486 24698 12538
rect 24698 12486 24712 12538
rect 24736 12486 24750 12538
rect 24750 12486 24762 12538
rect 24762 12486 24792 12538
rect 24816 12486 24826 12538
rect 24826 12486 24872 12538
rect 24576 12484 24632 12486
rect 24656 12484 24712 12486
rect 24736 12484 24792 12486
rect 24816 12484 24872 12486
rect 29300 14170 29356 14172
rect 29380 14170 29436 14172
rect 29460 14170 29516 14172
rect 29540 14170 29596 14172
rect 29300 14118 29346 14170
rect 29346 14118 29356 14170
rect 29380 14118 29410 14170
rect 29410 14118 29422 14170
rect 29422 14118 29436 14170
rect 29460 14118 29474 14170
rect 29474 14118 29486 14170
rect 29486 14118 29516 14170
rect 29540 14118 29550 14170
rect 29550 14118 29596 14170
rect 29300 14116 29356 14118
rect 29380 14116 29436 14118
rect 29460 14116 29516 14118
rect 29540 14116 29596 14118
rect 24576 11450 24632 11452
rect 24656 11450 24712 11452
rect 24736 11450 24792 11452
rect 24816 11450 24872 11452
rect 24576 11398 24622 11450
rect 24622 11398 24632 11450
rect 24656 11398 24686 11450
rect 24686 11398 24698 11450
rect 24698 11398 24712 11450
rect 24736 11398 24750 11450
rect 24750 11398 24762 11450
rect 24762 11398 24792 11450
rect 24816 11398 24826 11450
rect 24826 11398 24872 11450
rect 24576 11396 24632 11398
rect 24656 11396 24712 11398
rect 24736 11396 24792 11398
rect 24816 11396 24872 11398
rect 19852 9818 19908 9820
rect 19932 9818 19988 9820
rect 20012 9818 20068 9820
rect 20092 9818 20148 9820
rect 19852 9766 19898 9818
rect 19898 9766 19908 9818
rect 19932 9766 19962 9818
rect 19962 9766 19974 9818
rect 19974 9766 19988 9818
rect 20012 9766 20026 9818
rect 20026 9766 20038 9818
rect 20038 9766 20068 9818
rect 20092 9766 20102 9818
rect 20102 9766 20148 9818
rect 19852 9764 19908 9766
rect 19932 9764 19988 9766
rect 20012 9764 20068 9766
rect 20092 9764 20148 9766
rect 19852 8730 19908 8732
rect 19932 8730 19988 8732
rect 20012 8730 20068 8732
rect 20092 8730 20148 8732
rect 19852 8678 19898 8730
rect 19898 8678 19908 8730
rect 19932 8678 19962 8730
rect 19962 8678 19974 8730
rect 19974 8678 19988 8730
rect 20012 8678 20026 8730
rect 20026 8678 20038 8730
rect 20038 8678 20068 8730
rect 20092 8678 20102 8730
rect 20102 8678 20148 8730
rect 19852 8676 19908 8678
rect 19932 8676 19988 8678
rect 20012 8676 20068 8678
rect 20092 8676 20148 8678
rect 19852 7642 19908 7644
rect 19932 7642 19988 7644
rect 20012 7642 20068 7644
rect 20092 7642 20148 7644
rect 19852 7590 19898 7642
rect 19898 7590 19908 7642
rect 19932 7590 19962 7642
rect 19962 7590 19974 7642
rect 19974 7590 19988 7642
rect 20012 7590 20026 7642
rect 20026 7590 20038 7642
rect 20038 7590 20068 7642
rect 20092 7590 20102 7642
rect 20102 7590 20148 7642
rect 19852 7588 19908 7590
rect 19932 7588 19988 7590
rect 20012 7588 20068 7590
rect 20092 7588 20148 7590
rect 19852 6554 19908 6556
rect 19932 6554 19988 6556
rect 20012 6554 20068 6556
rect 20092 6554 20148 6556
rect 19852 6502 19898 6554
rect 19898 6502 19908 6554
rect 19932 6502 19962 6554
rect 19962 6502 19974 6554
rect 19974 6502 19988 6554
rect 20012 6502 20026 6554
rect 20026 6502 20038 6554
rect 20038 6502 20068 6554
rect 20092 6502 20102 6554
rect 20102 6502 20148 6554
rect 19852 6500 19908 6502
rect 19932 6500 19988 6502
rect 20012 6500 20068 6502
rect 20092 6500 20148 6502
rect 19852 5466 19908 5468
rect 19932 5466 19988 5468
rect 20012 5466 20068 5468
rect 20092 5466 20148 5468
rect 19852 5414 19898 5466
rect 19898 5414 19908 5466
rect 19932 5414 19962 5466
rect 19962 5414 19974 5466
rect 19974 5414 19988 5466
rect 20012 5414 20026 5466
rect 20026 5414 20038 5466
rect 20038 5414 20068 5466
rect 20092 5414 20102 5466
rect 20102 5414 20148 5466
rect 19852 5412 19908 5414
rect 19932 5412 19988 5414
rect 20012 5412 20068 5414
rect 20092 5412 20148 5414
rect 19852 4378 19908 4380
rect 19932 4378 19988 4380
rect 20012 4378 20068 4380
rect 20092 4378 20148 4380
rect 19852 4326 19898 4378
rect 19898 4326 19908 4378
rect 19932 4326 19962 4378
rect 19962 4326 19974 4378
rect 19974 4326 19988 4378
rect 20012 4326 20026 4378
rect 20026 4326 20038 4378
rect 20038 4326 20068 4378
rect 20092 4326 20102 4378
rect 20102 4326 20148 4378
rect 19852 4324 19908 4326
rect 19932 4324 19988 4326
rect 20012 4324 20068 4326
rect 20092 4324 20148 4326
rect 1490 1672 1546 1728
rect 10404 2202 10460 2204
rect 10484 2202 10540 2204
rect 10564 2202 10620 2204
rect 10644 2202 10700 2204
rect 10404 2150 10450 2202
rect 10450 2150 10460 2202
rect 10484 2150 10514 2202
rect 10514 2150 10526 2202
rect 10526 2150 10540 2202
rect 10564 2150 10578 2202
rect 10578 2150 10590 2202
rect 10590 2150 10620 2202
rect 10644 2150 10654 2202
rect 10654 2150 10700 2202
rect 10404 2148 10460 2150
rect 10484 2148 10540 2150
rect 10564 2148 10620 2150
rect 10644 2148 10700 2150
rect 19852 3290 19908 3292
rect 19932 3290 19988 3292
rect 20012 3290 20068 3292
rect 20092 3290 20148 3292
rect 19852 3238 19898 3290
rect 19898 3238 19908 3290
rect 19932 3238 19962 3290
rect 19962 3238 19974 3290
rect 19974 3238 19988 3290
rect 20012 3238 20026 3290
rect 20026 3238 20038 3290
rect 20038 3238 20068 3290
rect 20092 3238 20102 3290
rect 20102 3238 20148 3290
rect 19852 3236 19908 3238
rect 19932 3236 19988 3238
rect 20012 3236 20068 3238
rect 20092 3236 20148 3238
rect 24576 10362 24632 10364
rect 24656 10362 24712 10364
rect 24736 10362 24792 10364
rect 24816 10362 24872 10364
rect 24576 10310 24622 10362
rect 24622 10310 24632 10362
rect 24656 10310 24686 10362
rect 24686 10310 24698 10362
rect 24698 10310 24712 10362
rect 24736 10310 24750 10362
rect 24750 10310 24762 10362
rect 24762 10310 24792 10362
rect 24816 10310 24826 10362
rect 24826 10310 24872 10362
rect 24576 10308 24632 10310
rect 24656 10308 24712 10310
rect 24736 10308 24792 10310
rect 24816 10308 24872 10310
rect 29300 13082 29356 13084
rect 29380 13082 29436 13084
rect 29460 13082 29516 13084
rect 29540 13082 29596 13084
rect 29300 13030 29346 13082
rect 29346 13030 29356 13082
rect 29380 13030 29410 13082
rect 29410 13030 29422 13082
rect 29422 13030 29436 13082
rect 29460 13030 29474 13082
rect 29474 13030 29486 13082
rect 29486 13030 29516 13082
rect 29540 13030 29550 13082
rect 29550 13030 29596 13082
rect 29300 13028 29356 13030
rect 29380 13028 29436 13030
rect 29460 13028 29516 13030
rect 29540 13028 29596 13030
rect 34024 28858 34080 28860
rect 34104 28858 34160 28860
rect 34184 28858 34240 28860
rect 34264 28858 34320 28860
rect 34024 28806 34070 28858
rect 34070 28806 34080 28858
rect 34104 28806 34134 28858
rect 34134 28806 34146 28858
rect 34146 28806 34160 28858
rect 34184 28806 34198 28858
rect 34198 28806 34210 28858
rect 34210 28806 34240 28858
rect 34264 28806 34274 28858
rect 34274 28806 34320 28858
rect 34024 28804 34080 28806
rect 34104 28804 34160 28806
rect 34184 28804 34240 28806
rect 34264 28804 34320 28806
rect 34024 27770 34080 27772
rect 34104 27770 34160 27772
rect 34184 27770 34240 27772
rect 34264 27770 34320 27772
rect 34024 27718 34070 27770
rect 34070 27718 34080 27770
rect 34104 27718 34134 27770
rect 34134 27718 34146 27770
rect 34146 27718 34160 27770
rect 34184 27718 34198 27770
rect 34198 27718 34210 27770
rect 34210 27718 34240 27770
rect 34264 27718 34274 27770
rect 34274 27718 34320 27770
rect 34024 27716 34080 27718
rect 34104 27716 34160 27718
rect 34184 27716 34240 27718
rect 34264 27716 34320 27718
rect 29300 11994 29356 11996
rect 29380 11994 29436 11996
rect 29460 11994 29516 11996
rect 29540 11994 29596 11996
rect 29300 11942 29346 11994
rect 29346 11942 29356 11994
rect 29380 11942 29410 11994
rect 29410 11942 29422 11994
rect 29422 11942 29436 11994
rect 29460 11942 29474 11994
rect 29474 11942 29486 11994
rect 29486 11942 29516 11994
rect 29540 11942 29550 11994
rect 29550 11942 29596 11994
rect 29300 11940 29356 11942
rect 29380 11940 29436 11942
rect 29460 11940 29516 11942
rect 29540 11940 29596 11942
rect 29300 10906 29356 10908
rect 29380 10906 29436 10908
rect 29460 10906 29516 10908
rect 29540 10906 29596 10908
rect 29300 10854 29346 10906
rect 29346 10854 29356 10906
rect 29380 10854 29410 10906
rect 29410 10854 29422 10906
rect 29422 10854 29436 10906
rect 29460 10854 29474 10906
rect 29474 10854 29486 10906
rect 29486 10854 29516 10906
rect 29540 10854 29550 10906
rect 29550 10854 29596 10906
rect 29300 10852 29356 10854
rect 29380 10852 29436 10854
rect 29460 10852 29516 10854
rect 29540 10852 29596 10854
rect 24576 9274 24632 9276
rect 24656 9274 24712 9276
rect 24736 9274 24792 9276
rect 24816 9274 24872 9276
rect 24576 9222 24622 9274
rect 24622 9222 24632 9274
rect 24656 9222 24686 9274
rect 24686 9222 24698 9274
rect 24698 9222 24712 9274
rect 24736 9222 24750 9274
rect 24750 9222 24762 9274
rect 24762 9222 24792 9274
rect 24816 9222 24826 9274
rect 24826 9222 24872 9274
rect 24576 9220 24632 9222
rect 24656 9220 24712 9222
rect 24736 9220 24792 9222
rect 24816 9220 24872 9222
rect 29300 9818 29356 9820
rect 29380 9818 29436 9820
rect 29460 9818 29516 9820
rect 29540 9818 29596 9820
rect 29300 9766 29346 9818
rect 29346 9766 29356 9818
rect 29380 9766 29410 9818
rect 29410 9766 29422 9818
rect 29422 9766 29436 9818
rect 29460 9766 29474 9818
rect 29474 9766 29486 9818
rect 29486 9766 29516 9818
rect 29540 9766 29550 9818
rect 29550 9766 29596 9818
rect 29300 9764 29356 9766
rect 29380 9764 29436 9766
rect 29460 9764 29516 9766
rect 29540 9764 29596 9766
rect 29300 8730 29356 8732
rect 29380 8730 29436 8732
rect 29460 8730 29516 8732
rect 29540 8730 29596 8732
rect 29300 8678 29346 8730
rect 29346 8678 29356 8730
rect 29380 8678 29410 8730
rect 29410 8678 29422 8730
rect 29422 8678 29436 8730
rect 29460 8678 29474 8730
rect 29474 8678 29486 8730
rect 29486 8678 29516 8730
rect 29540 8678 29550 8730
rect 29550 8678 29596 8730
rect 29300 8676 29356 8678
rect 29380 8676 29436 8678
rect 29460 8676 29516 8678
rect 29540 8676 29596 8678
rect 24576 8186 24632 8188
rect 24656 8186 24712 8188
rect 24736 8186 24792 8188
rect 24816 8186 24872 8188
rect 24576 8134 24622 8186
rect 24622 8134 24632 8186
rect 24656 8134 24686 8186
rect 24686 8134 24698 8186
rect 24698 8134 24712 8186
rect 24736 8134 24750 8186
rect 24750 8134 24762 8186
rect 24762 8134 24792 8186
rect 24816 8134 24826 8186
rect 24826 8134 24872 8186
rect 24576 8132 24632 8134
rect 24656 8132 24712 8134
rect 24736 8132 24792 8134
rect 24816 8132 24872 8134
rect 29300 7642 29356 7644
rect 29380 7642 29436 7644
rect 29460 7642 29516 7644
rect 29540 7642 29596 7644
rect 29300 7590 29346 7642
rect 29346 7590 29356 7642
rect 29380 7590 29410 7642
rect 29410 7590 29422 7642
rect 29422 7590 29436 7642
rect 29460 7590 29474 7642
rect 29474 7590 29486 7642
rect 29486 7590 29516 7642
rect 29540 7590 29550 7642
rect 29550 7590 29596 7642
rect 29300 7588 29356 7590
rect 29380 7588 29436 7590
rect 29460 7588 29516 7590
rect 29540 7588 29596 7590
rect 24576 7098 24632 7100
rect 24656 7098 24712 7100
rect 24736 7098 24792 7100
rect 24816 7098 24872 7100
rect 24576 7046 24622 7098
rect 24622 7046 24632 7098
rect 24656 7046 24686 7098
rect 24686 7046 24698 7098
rect 24698 7046 24712 7098
rect 24736 7046 24750 7098
rect 24750 7046 24762 7098
rect 24762 7046 24792 7098
rect 24816 7046 24826 7098
rect 24826 7046 24872 7098
rect 24576 7044 24632 7046
rect 24656 7044 24712 7046
rect 24736 7044 24792 7046
rect 24816 7044 24872 7046
rect 24576 6010 24632 6012
rect 24656 6010 24712 6012
rect 24736 6010 24792 6012
rect 24816 6010 24872 6012
rect 24576 5958 24622 6010
rect 24622 5958 24632 6010
rect 24656 5958 24686 6010
rect 24686 5958 24698 6010
rect 24698 5958 24712 6010
rect 24736 5958 24750 6010
rect 24750 5958 24762 6010
rect 24762 5958 24792 6010
rect 24816 5958 24826 6010
rect 24826 5958 24872 6010
rect 24576 5956 24632 5958
rect 24656 5956 24712 5958
rect 24736 5956 24792 5958
rect 24816 5956 24872 5958
rect 29300 6554 29356 6556
rect 29380 6554 29436 6556
rect 29460 6554 29516 6556
rect 29540 6554 29596 6556
rect 29300 6502 29346 6554
rect 29346 6502 29356 6554
rect 29380 6502 29410 6554
rect 29410 6502 29422 6554
rect 29422 6502 29436 6554
rect 29460 6502 29474 6554
rect 29474 6502 29486 6554
rect 29486 6502 29516 6554
rect 29540 6502 29550 6554
rect 29550 6502 29596 6554
rect 29300 6500 29356 6502
rect 29380 6500 29436 6502
rect 29460 6500 29516 6502
rect 29540 6500 29596 6502
rect 34024 26682 34080 26684
rect 34104 26682 34160 26684
rect 34184 26682 34240 26684
rect 34264 26682 34320 26684
rect 34024 26630 34070 26682
rect 34070 26630 34080 26682
rect 34104 26630 34134 26682
rect 34134 26630 34146 26682
rect 34146 26630 34160 26682
rect 34184 26630 34198 26682
rect 34198 26630 34210 26682
rect 34210 26630 34240 26682
rect 34264 26630 34274 26682
rect 34274 26630 34320 26682
rect 34024 26628 34080 26630
rect 34104 26628 34160 26630
rect 34184 26628 34240 26630
rect 34264 26628 34320 26630
rect 34024 25594 34080 25596
rect 34104 25594 34160 25596
rect 34184 25594 34240 25596
rect 34264 25594 34320 25596
rect 34024 25542 34070 25594
rect 34070 25542 34080 25594
rect 34104 25542 34134 25594
rect 34134 25542 34146 25594
rect 34146 25542 34160 25594
rect 34184 25542 34198 25594
rect 34198 25542 34210 25594
rect 34210 25542 34240 25594
rect 34264 25542 34274 25594
rect 34274 25542 34320 25594
rect 34024 25540 34080 25542
rect 34104 25540 34160 25542
rect 34184 25540 34240 25542
rect 34264 25540 34320 25542
rect 34024 24506 34080 24508
rect 34104 24506 34160 24508
rect 34184 24506 34240 24508
rect 34264 24506 34320 24508
rect 34024 24454 34070 24506
rect 34070 24454 34080 24506
rect 34104 24454 34134 24506
rect 34134 24454 34146 24506
rect 34146 24454 34160 24506
rect 34184 24454 34198 24506
rect 34198 24454 34210 24506
rect 34210 24454 34240 24506
rect 34264 24454 34274 24506
rect 34274 24454 34320 24506
rect 34024 24452 34080 24454
rect 34104 24452 34160 24454
rect 34184 24452 34240 24454
rect 34264 24452 34320 24454
rect 34024 23418 34080 23420
rect 34104 23418 34160 23420
rect 34184 23418 34240 23420
rect 34264 23418 34320 23420
rect 34024 23366 34070 23418
rect 34070 23366 34080 23418
rect 34104 23366 34134 23418
rect 34134 23366 34146 23418
rect 34146 23366 34160 23418
rect 34184 23366 34198 23418
rect 34198 23366 34210 23418
rect 34210 23366 34240 23418
rect 34264 23366 34274 23418
rect 34274 23366 34320 23418
rect 34024 23364 34080 23366
rect 34104 23364 34160 23366
rect 34184 23364 34240 23366
rect 34264 23364 34320 23366
rect 34024 22330 34080 22332
rect 34104 22330 34160 22332
rect 34184 22330 34240 22332
rect 34264 22330 34320 22332
rect 34024 22278 34070 22330
rect 34070 22278 34080 22330
rect 34104 22278 34134 22330
rect 34134 22278 34146 22330
rect 34146 22278 34160 22330
rect 34184 22278 34198 22330
rect 34198 22278 34210 22330
rect 34210 22278 34240 22330
rect 34264 22278 34274 22330
rect 34274 22278 34320 22330
rect 34024 22276 34080 22278
rect 34104 22276 34160 22278
rect 34184 22276 34240 22278
rect 34264 22276 34320 22278
rect 34024 21242 34080 21244
rect 34104 21242 34160 21244
rect 34184 21242 34240 21244
rect 34264 21242 34320 21244
rect 34024 21190 34070 21242
rect 34070 21190 34080 21242
rect 34104 21190 34134 21242
rect 34134 21190 34146 21242
rect 34146 21190 34160 21242
rect 34184 21190 34198 21242
rect 34198 21190 34210 21242
rect 34210 21190 34240 21242
rect 34264 21190 34274 21242
rect 34274 21190 34320 21242
rect 34024 21188 34080 21190
rect 34104 21188 34160 21190
rect 34184 21188 34240 21190
rect 34264 21188 34320 21190
rect 34024 20154 34080 20156
rect 34104 20154 34160 20156
rect 34184 20154 34240 20156
rect 34264 20154 34320 20156
rect 34024 20102 34070 20154
rect 34070 20102 34080 20154
rect 34104 20102 34134 20154
rect 34134 20102 34146 20154
rect 34146 20102 34160 20154
rect 34184 20102 34198 20154
rect 34198 20102 34210 20154
rect 34210 20102 34240 20154
rect 34264 20102 34274 20154
rect 34274 20102 34320 20154
rect 34024 20100 34080 20102
rect 34104 20100 34160 20102
rect 34184 20100 34240 20102
rect 34264 20100 34320 20102
rect 34024 19066 34080 19068
rect 34104 19066 34160 19068
rect 34184 19066 34240 19068
rect 34264 19066 34320 19068
rect 34024 19014 34070 19066
rect 34070 19014 34080 19066
rect 34104 19014 34134 19066
rect 34134 19014 34146 19066
rect 34146 19014 34160 19066
rect 34184 19014 34198 19066
rect 34198 19014 34210 19066
rect 34210 19014 34240 19066
rect 34264 19014 34274 19066
rect 34274 19014 34320 19066
rect 34024 19012 34080 19014
rect 34104 19012 34160 19014
rect 34184 19012 34240 19014
rect 34264 19012 34320 19014
rect 34024 17978 34080 17980
rect 34104 17978 34160 17980
rect 34184 17978 34240 17980
rect 34264 17978 34320 17980
rect 34024 17926 34070 17978
rect 34070 17926 34080 17978
rect 34104 17926 34134 17978
rect 34134 17926 34146 17978
rect 34146 17926 34160 17978
rect 34184 17926 34198 17978
rect 34198 17926 34210 17978
rect 34210 17926 34240 17978
rect 34264 17926 34274 17978
rect 34274 17926 34320 17978
rect 34024 17924 34080 17926
rect 34104 17924 34160 17926
rect 34184 17924 34240 17926
rect 34264 17924 34320 17926
rect 34024 16890 34080 16892
rect 34104 16890 34160 16892
rect 34184 16890 34240 16892
rect 34264 16890 34320 16892
rect 34024 16838 34070 16890
rect 34070 16838 34080 16890
rect 34104 16838 34134 16890
rect 34134 16838 34146 16890
rect 34146 16838 34160 16890
rect 34184 16838 34198 16890
rect 34198 16838 34210 16890
rect 34210 16838 34240 16890
rect 34264 16838 34274 16890
rect 34274 16838 34320 16890
rect 34024 16836 34080 16838
rect 34104 16836 34160 16838
rect 34184 16836 34240 16838
rect 34264 16836 34320 16838
rect 34024 15802 34080 15804
rect 34104 15802 34160 15804
rect 34184 15802 34240 15804
rect 34264 15802 34320 15804
rect 34024 15750 34070 15802
rect 34070 15750 34080 15802
rect 34104 15750 34134 15802
rect 34134 15750 34146 15802
rect 34146 15750 34160 15802
rect 34184 15750 34198 15802
rect 34198 15750 34210 15802
rect 34210 15750 34240 15802
rect 34264 15750 34274 15802
rect 34274 15750 34320 15802
rect 34024 15748 34080 15750
rect 34104 15748 34160 15750
rect 34184 15748 34240 15750
rect 34264 15748 34320 15750
rect 34024 14714 34080 14716
rect 34104 14714 34160 14716
rect 34184 14714 34240 14716
rect 34264 14714 34320 14716
rect 34024 14662 34070 14714
rect 34070 14662 34080 14714
rect 34104 14662 34134 14714
rect 34134 14662 34146 14714
rect 34146 14662 34160 14714
rect 34184 14662 34198 14714
rect 34198 14662 34210 14714
rect 34210 14662 34240 14714
rect 34264 14662 34274 14714
rect 34274 14662 34320 14714
rect 34024 14660 34080 14662
rect 34104 14660 34160 14662
rect 34184 14660 34240 14662
rect 34264 14660 34320 14662
rect 34024 13626 34080 13628
rect 34104 13626 34160 13628
rect 34184 13626 34240 13628
rect 34264 13626 34320 13628
rect 34024 13574 34070 13626
rect 34070 13574 34080 13626
rect 34104 13574 34134 13626
rect 34134 13574 34146 13626
rect 34146 13574 34160 13626
rect 34184 13574 34198 13626
rect 34198 13574 34210 13626
rect 34210 13574 34240 13626
rect 34264 13574 34274 13626
rect 34274 13574 34320 13626
rect 34024 13572 34080 13574
rect 34104 13572 34160 13574
rect 34184 13572 34240 13574
rect 34264 13572 34320 13574
rect 34024 12538 34080 12540
rect 34104 12538 34160 12540
rect 34184 12538 34240 12540
rect 34264 12538 34320 12540
rect 34024 12486 34070 12538
rect 34070 12486 34080 12538
rect 34104 12486 34134 12538
rect 34134 12486 34146 12538
rect 34146 12486 34160 12538
rect 34184 12486 34198 12538
rect 34198 12486 34210 12538
rect 34210 12486 34240 12538
rect 34264 12486 34274 12538
rect 34274 12486 34320 12538
rect 34024 12484 34080 12486
rect 34104 12484 34160 12486
rect 34184 12484 34240 12486
rect 34264 12484 34320 12486
rect 34024 11450 34080 11452
rect 34104 11450 34160 11452
rect 34184 11450 34240 11452
rect 34264 11450 34320 11452
rect 34024 11398 34070 11450
rect 34070 11398 34080 11450
rect 34104 11398 34134 11450
rect 34134 11398 34146 11450
rect 34146 11398 34160 11450
rect 34184 11398 34198 11450
rect 34198 11398 34210 11450
rect 34210 11398 34240 11450
rect 34264 11398 34274 11450
rect 34274 11398 34320 11450
rect 34024 11396 34080 11398
rect 34104 11396 34160 11398
rect 34184 11396 34240 11398
rect 34264 11396 34320 11398
rect 34024 10362 34080 10364
rect 34104 10362 34160 10364
rect 34184 10362 34240 10364
rect 34264 10362 34320 10364
rect 34024 10310 34070 10362
rect 34070 10310 34080 10362
rect 34104 10310 34134 10362
rect 34134 10310 34146 10362
rect 34146 10310 34160 10362
rect 34184 10310 34198 10362
rect 34198 10310 34210 10362
rect 34210 10310 34240 10362
rect 34264 10310 34274 10362
rect 34274 10310 34320 10362
rect 34024 10308 34080 10310
rect 34104 10308 34160 10310
rect 34184 10308 34240 10310
rect 34264 10308 34320 10310
rect 34024 9274 34080 9276
rect 34104 9274 34160 9276
rect 34184 9274 34240 9276
rect 34264 9274 34320 9276
rect 34024 9222 34070 9274
rect 34070 9222 34080 9274
rect 34104 9222 34134 9274
rect 34134 9222 34146 9274
rect 34146 9222 34160 9274
rect 34184 9222 34198 9274
rect 34198 9222 34210 9274
rect 34210 9222 34240 9274
rect 34264 9222 34274 9274
rect 34274 9222 34320 9274
rect 34024 9220 34080 9222
rect 34104 9220 34160 9222
rect 34184 9220 34240 9222
rect 34264 9220 34320 9222
rect 34024 8186 34080 8188
rect 34104 8186 34160 8188
rect 34184 8186 34240 8188
rect 34264 8186 34320 8188
rect 34024 8134 34070 8186
rect 34070 8134 34080 8186
rect 34104 8134 34134 8186
rect 34134 8134 34146 8186
rect 34146 8134 34160 8186
rect 34184 8134 34198 8186
rect 34198 8134 34210 8186
rect 34210 8134 34240 8186
rect 34264 8134 34274 8186
rect 34274 8134 34320 8186
rect 34024 8132 34080 8134
rect 34104 8132 34160 8134
rect 34184 8132 34240 8134
rect 34264 8132 34320 8134
rect 34024 7098 34080 7100
rect 34104 7098 34160 7100
rect 34184 7098 34240 7100
rect 34264 7098 34320 7100
rect 34024 7046 34070 7098
rect 34070 7046 34080 7098
rect 34104 7046 34134 7098
rect 34134 7046 34146 7098
rect 34146 7046 34160 7098
rect 34184 7046 34198 7098
rect 34198 7046 34210 7098
rect 34210 7046 34240 7098
rect 34264 7046 34274 7098
rect 34274 7046 34320 7098
rect 34024 7044 34080 7046
rect 34104 7044 34160 7046
rect 34184 7044 34240 7046
rect 34264 7044 34320 7046
rect 24576 4922 24632 4924
rect 24656 4922 24712 4924
rect 24736 4922 24792 4924
rect 24816 4922 24872 4924
rect 24576 4870 24622 4922
rect 24622 4870 24632 4922
rect 24656 4870 24686 4922
rect 24686 4870 24698 4922
rect 24698 4870 24712 4922
rect 24736 4870 24750 4922
rect 24750 4870 24762 4922
rect 24762 4870 24792 4922
rect 24816 4870 24826 4922
rect 24826 4870 24872 4922
rect 24576 4868 24632 4870
rect 24656 4868 24712 4870
rect 24736 4868 24792 4870
rect 24816 4868 24872 4870
rect 24576 3834 24632 3836
rect 24656 3834 24712 3836
rect 24736 3834 24792 3836
rect 24816 3834 24872 3836
rect 24576 3782 24622 3834
rect 24622 3782 24632 3834
rect 24656 3782 24686 3834
rect 24686 3782 24698 3834
rect 24698 3782 24712 3834
rect 24736 3782 24750 3834
rect 24750 3782 24762 3834
rect 24762 3782 24792 3834
rect 24816 3782 24826 3834
rect 24826 3782 24872 3834
rect 24576 3780 24632 3782
rect 24656 3780 24712 3782
rect 24736 3780 24792 3782
rect 24816 3780 24872 3782
rect 29300 5466 29356 5468
rect 29380 5466 29436 5468
rect 29460 5466 29516 5468
rect 29540 5466 29596 5468
rect 29300 5414 29346 5466
rect 29346 5414 29356 5466
rect 29380 5414 29410 5466
rect 29410 5414 29422 5466
rect 29422 5414 29436 5466
rect 29460 5414 29474 5466
rect 29474 5414 29486 5466
rect 29486 5414 29516 5466
rect 29540 5414 29550 5466
rect 29550 5414 29596 5466
rect 29300 5412 29356 5414
rect 29380 5412 29436 5414
rect 29460 5412 29516 5414
rect 29540 5412 29596 5414
rect 29300 4378 29356 4380
rect 29380 4378 29436 4380
rect 29460 4378 29516 4380
rect 29540 4378 29596 4380
rect 29300 4326 29346 4378
rect 29346 4326 29356 4378
rect 29380 4326 29410 4378
rect 29410 4326 29422 4378
rect 29422 4326 29436 4378
rect 29460 4326 29474 4378
rect 29474 4326 29486 4378
rect 29486 4326 29516 4378
rect 29540 4326 29550 4378
rect 29550 4326 29596 4378
rect 29300 4324 29356 4326
rect 29380 4324 29436 4326
rect 29460 4324 29516 4326
rect 29540 4324 29596 4326
rect 34024 6010 34080 6012
rect 34104 6010 34160 6012
rect 34184 6010 34240 6012
rect 34264 6010 34320 6012
rect 34024 5958 34070 6010
rect 34070 5958 34080 6010
rect 34104 5958 34134 6010
rect 34134 5958 34146 6010
rect 34146 5958 34160 6010
rect 34184 5958 34198 6010
rect 34198 5958 34210 6010
rect 34210 5958 34240 6010
rect 34264 5958 34274 6010
rect 34274 5958 34320 6010
rect 34024 5956 34080 5958
rect 34104 5956 34160 5958
rect 34184 5956 34240 5958
rect 34264 5956 34320 5958
rect 34024 4922 34080 4924
rect 34104 4922 34160 4924
rect 34184 4922 34240 4924
rect 34264 4922 34320 4924
rect 34024 4870 34070 4922
rect 34070 4870 34080 4922
rect 34104 4870 34134 4922
rect 34134 4870 34146 4922
rect 34146 4870 34160 4922
rect 34184 4870 34198 4922
rect 34198 4870 34210 4922
rect 34210 4870 34240 4922
rect 34264 4870 34274 4922
rect 34274 4870 34320 4922
rect 34024 4868 34080 4870
rect 34104 4868 34160 4870
rect 34184 4868 34240 4870
rect 34264 4868 34320 4870
rect 24576 2746 24632 2748
rect 24656 2746 24712 2748
rect 24736 2746 24792 2748
rect 24816 2746 24872 2748
rect 24576 2694 24622 2746
rect 24622 2694 24632 2746
rect 24656 2694 24686 2746
rect 24686 2694 24698 2746
rect 24698 2694 24712 2746
rect 24736 2694 24750 2746
rect 24750 2694 24762 2746
rect 24762 2694 24792 2746
rect 24816 2694 24826 2746
rect 24826 2694 24872 2746
rect 24576 2692 24632 2694
rect 24656 2692 24712 2694
rect 24736 2692 24792 2694
rect 24816 2692 24872 2694
rect 29300 3290 29356 3292
rect 29380 3290 29436 3292
rect 29460 3290 29516 3292
rect 29540 3290 29596 3292
rect 29300 3238 29346 3290
rect 29346 3238 29356 3290
rect 29380 3238 29410 3290
rect 29410 3238 29422 3290
rect 29422 3238 29436 3290
rect 29460 3238 29474 3290
rect 29474 3238 29486 3290
rect 29486 3238 29516 3290
rect 29540 3238 29550 3290
rect 29550 3238 29596 3290
rect 29300 3236 29356 3238
rect 29380 3236 29436 3238
rect 29460 3236 29516 3238
rect 29540 3236 29596 3238
rect 34024 3834 34080 3836
rect 34104 3834 34160 3836
rect 34184 3834 34240 3836
rect 34264 3834 34320 3836
rect 34024 3782 34070 3834
rect 34070 3782 34080 3834
rect 34104 3782 34134 3834
rect 34134 3782 34146 3834
rect 34146 3782 34160 3834
rect 34184 3782 34198 3834
rect 34198 3782 34210 3834
rect 34210 3782 34240 3834
rect 34264 3782 34274 3834
rect 34274 3782 34320 3834
rect 34024 3780 34080 3782
rect 34104 3780 34160 3782
rect 34184 3780 34240 3782
rect 34264 3780 34320 3782
rect 34024 2746 34080 2748
rect 34104 2746 34160 2748
rect 34184 2746 34240 2748
rect 34264 2746 34320 2748
rect 34024 2694 34070 2746
rect 34070 2694 34080 2746
rect 34104 2694 34134 2746
rect 34134 2694 34146 2746
rect 34146 2694 34160 2746
rect 34184 2694 34198 2746
rect 34198 2694 34210 2746
rect 34210 2694 34240 2746
rect 34264 2694 34274 2746
rect 34274 2694 34320 2746
rect 34024 2692 34080 2694
rect 34104 2692 34160 2694
rect 34184 2692 34240 2694
rect 34264 2692 34320 2694
rect 19852 2202 19908 2204
rect 19932 2202 19988 2204
rect 20012 2202 20068 2204
rect 20092 2202 20148 2204
rect 19852 2150 19898 2202
rect 19898 2150 19908 2202
rect 19932 2150 19962 2202
rect 19962 2150 19974 2202
rect 19974 2150 19988 2202
rect 20012 2150 20026 2202
rect 20026 2150 20038 2202
rect 20038 2150 20068 2202
rect 20092 2150 20102 2202
rect 20102 2150 20148 2202
rect 19852 2148 19908 2150
rect 19932 2148 19988 2150
rect 20012 2148 20068 2150
rect 20092 2148 20148 2150
rect 29300 2202 29356 2204
rect 29380 2202 29436 2204
rect 29460 2202 29516 2204
rect 29540 2202 29596 2204
rect 29300 2150 29346 2202
rect 29346 2150 29356 2202
rect 29380 2150 29410 2202
rect 29410 2150 29422 2202
rect 29422 2150 29436 2202
rect 29460 2150 29474 2202
rect 29474 2150 29486 2202
rect 29486 2150 29516 2202
rect 29540 2150 29550 2202
rect 29550 2150 29596 2202
rect 29300 2148 29356 2150
rect 29380 2148 29436 2150
rect 29460 2148 29516 2150
rect 29540 2148 29596 2150
<< metal3 >>
rect 0 34370 800 34400
rect 1393 34370 1459 34373
rect 0 34368 1459 34370
rect 0 34312 1398 34368
rect 1454 34312 1459 34368
rect 0 34310 1459 34312
rect 0 34280 800 34310
rect 1393 34307 1459 34310
rect 10394 33760 10710 33761
rect 10394 33696 10400 33760
rect 10464 33696 10480 33760
rect 10544 33696 10560 33760
rect 10624 33696 10640 33760
rect 10704 33696 10710 33760
rect 10394 33695 10710 33696
rect 19842 33760 20158 33761
rect 19842 33696 19848 33760
rect 19912 33696 19928 33760
rect 19992 33696 20008 33760
rect 20072 33696 20088 33760
rect 20152 33696 20158 33760
rect 19842 33695 20158 33696
rect 29290 33760 29606 33761
rect 29290 33696 29296 33760
rect 29360 33696 29376 33760
rect 29440 33696 29456 33760
rect 29520 33696 29536 33760
rect 29600 33696 29606 33760
rect 29290 33695 29606 33696
rect 5670 33216 5986 33217
rect 5670 33152 5676 33216
rect 5740 33152 5756 33216
rect 5820 33152 5836 33216
rect 5900 33152 5916 33216
rect 5980 33152 5986 33216
rect 5670 33151 5986 33152
rect 15118 33216 15434 33217
rect 15118 33152 15124 33216
rect 15188 33152 15204 33216
rect 15268 33152 15284 33216
rect 15348 33152 15364 33216
rect 15428 33152 15434 33216
rect 15118 33151 15434 33152
rect 24566 33216 24882 33217
rect 24566 33152 24572 33216
rect 24636 33152 24652 33216
rect 24716 33152 24732 33216
rect 24796 33152 24812 33216
rect 24876 33152 24882 33216
rect 24566 33151 24882 33152
rect 34014 33216 34330 33217
rect 34014 33152 34020 33216
rect 34084 33152 34100 33216
rect 34164 33152 34180 33216
rect 34244 33152 34260 33216
rect 34324 33152 34330 33216
rect 34014 33151 34330 33152
rect 0 33010 800 33040
rect 1485 33010 1551 33013
rect 0 33008 1551 33010
rect 0 32952 1490 33008
rect 1546 32952 1551 33008
rect 0 32950 1551 32952
rect 0 32920 800 32950
rect 1485 32947 1551 32950
rect 10394 32672 10710 32673
rect 10394 32608 10400 32672
rect 10464 32608 10480 32672
rect 10544 32608 10560 32672
rect 10624 32608 10640 32672
rect 10704 32608 10710 32672
rect 10394 32607 10710 32608
rect 19842 32672 20158 32673
rect 19842 32608 19848 32672
rect 19912 32608 19928 32672
rect 19992 32608 20008 32672
rect 20072 32608 20088 32672
rect 20152 32608 20158 32672
rect 19842 32607 20158 32608
rect 29290 32672 29606 32673
rect 29290 32608 29296 32672
rect 29360 32608 29376 32672
rect 29440 32608 29456 32672
rect 29520 32608 29536 32672
rect 29600 32608 29606 32672
rect 29290 32607 29606 32608
rect 5670 32128 5986 32129
rect 5670 32064 5676 32128
rect 5740 32064 5756 32128
rect 5820 32064 5836 32128
rect 5900 32064 5916 32128
rect 5980 32064 5986 32128
rect 5670 32063 5986 32064
rect 15118 32128 15434 32129
rect 15118 32064 15124 32128
rect 15188 32064 15204 32128
rect 15268 32064 15284 32128
rect 15348 32064 15364 32128
rect 15428 32064 15434 32128
rect 15118 32063 15434 32064
rect 24566 32128 24882 32129
rect 24566 32064 24572 32128
rect 24636 32064 24652 32128
rect 24716 32064 24732 32128
rect 24796 32064 24812 32128
rect 24876 32064 24882 32128
rect 24566 32063 24882 32064
rect 34014 32128 34330 32129
rect 34014 32064 34020 32128
rect 34084 32064 34100 32128
rect 34164 32064 34180 32128
rect 34244 32064 34260 32128
rect 34324 32064 34330 32128
rect 34014 32063 34330 32064
rect 0 31650 800 31680
rect 1485 31650 1551 31653
rect 0 31648 1551 31650
rect 0 31592 1490 31648
rect 1546 31592 1551 31648
rect 0 31590 1551 31592
rect 0 31560 800 31590
rect 1485 31587 1551 31590
rect 10394 31584 10710 31585
rect 10394 31520 10400 31584
rect 10464 31520 10480 31584
rect 10544 31520 10560 31584
rect 10624 31520 10640 31584
rect 10704 31520 10710 31584
rect 10394 31519 10710 31520
rect 19842 31584 20158 31585
rect 19842 31520 19848 31584
rect 19912 31520 19928 31584
rect 19992 31520 20008 31584
rect 20072 31520 20088 31584
rect 20152 31520 20158 31584
rect 19842 31519 20158 31520
rect 29290 31584 29606 31585
rect 29290 31520 29296 31584
rect 29360 31520 29376 31584
rect 29440 31520 29456 31584
rect 29520 31520 29536 31584
rect 29600 31520 29606 31584
rect 29290 31519 29606 31520
rect 5670 31040 5986 31041
rect 5670 30976 5676 31040
rect 5740 30976 5756 31040
rect 5820 30976 5836 31040
rect 5900 30976 5916 31040
rect 5980 30976 5986 31040
rect 5670 30975 5986 30976
rect 15118 31040 15434 31041
rect 15118 30976 15124 31040
rect 15188 30976 15204 31040
rect 15268 30976 15284 31040
rect 15348 30976 15364 31040
rect 15428 30976 15434 31040
rect 15118 30975 15434 30976
rect 24566 31040 24882 31041
rect 24566 30976 24572 31040
rect 24636 30976 24652 31040
rect 24716 30976 24732 31040
rect 24796 30976 24812 31040
rect 24876 30976 24882 31040
rect 24566 30975 24882 30976
rect 34014 31040 34330 31041
rect 34014 30976 34020 31040
rect 34084 30976 34100 31040
rect 34164 30976 34180 31040
rect 34244 30976 34260 31040
rect 34324 30976 34330 31040
rect 34014 30975 34330 30976
rect 10394 30496 10710 30497
rect 10394 30432 10400 30496
rect 10464 30432 10480 30496
rect 10544 30432 10560 30496
rect 10624 30432 10640 30496
rect 10704 30432 10710 30496
rect 10394 30431 10710 30432
rect 19842 30496 20158 30497
rect 19842 30432 19848 30496
rect 19912 30432 19928 30496
rect 19992 30432 20008 30496
rect 20072 30432 20088 30496
rect 20152 30432 20158 30496
rect 19842 30431 20158 30432
rect 29290 30496 29606 30497
rect 29290 30432 29296 30496
rect 29360 30432 29376 30496
rect 29440 30432 29456 30496
rect 29520 30432 29536 30496
rect 29600 30432 29606 30496
rect 29290 30431 29606 30432
rect 0 30290 800 30320
rect 1485 30290 1551 30293
rect 0 30288 1551 30290
rect 0 30232 1490 30288
rect 1546 30232 1551 30288
rect 0 30230 1551 30232
rect 0 30200 800 30230
rect 1485 30227 1551 30230
rect 5670 29952 5986 29953
rect 5670 29888 5676 29952
rect 5740 29888 5756 29952
rect 5820 29888 5836 29952
rect 5900 29888 5916 29952
rect 5980 29888 5986 29952
rect 5670 29887 5986 29888
rect 15118 29952 15434 29953
rect 15118 29888 15124 29952
rect 15188 29888 15204 29952
rect 15268 29888 15284 29952
rect 15348 29888 15364 29952
rect 15428 29888 15434 29952
rect 15118 29887 15434 29888
rect 24566 29952 24882 29953
rect 24566 29888 24572 29952
rect 24636 29888 24652 29952
rect 24716 29888 24732 29952
rect 24796 29888 24812 29952
rect 24876 29888 24882 29952
rect 24566 29887 24882 29888
rect 34014 29952 34330 29953
rect 34014 29888 34020 29952
rect 34084 29888 34100 29952
rect 34164 29888 34180 29952
rect 34244 29888 34260 29952
rect 34324 29888 34330 29952
rect 34014 29887 34330 29888
rect 10394 29408 10710 29409
rect 10394 29344 10400 29408
rect 10464 29344 10480 29408
rect 10544 29344 10560 29408
rect 10624 29344 10640 29408
rect 10704 29344 10710 29408
rect 10394 29343 10710 29344
rect 19842 29408 20158 29409
rect 19842 29344 19848 29408
rect 19912 29344 19928 29408
rect 19992 29344 20008 29408
rect 20072 29344 20088 29408
rect 20152 29344 20158 29408
rect 19842 29343 20158 29344
rect 29290 29408 29606 29409
rect 29290 29344 29296 29408
rect 29360 29344 29376 29408
rect 29440 29344 29456 29408
rect 29520 29344 29536 29408
rect 29600 29344 29606 29408
rect 29290 29343 29606 29344
rect 0 28930 800 28960
rect 1485 28930 1551 28933
rect 0 28928 1551 28930
rect 0 28872 1490 28928
rect 1546 28872 1551 28928
rect 0 28870 1551 28872
rect 0 28840 800 28870
rect 1485 28867 1551 28870
rect 5670 28864 5986 28865
rect 5670 28800 5676 28864
rect 5740 28800 5756 28864
rect 5820 28800 5836 28864
rect 5900 28800 5916 28864
rect 5980 28800 5986 28864
rect 5670 28799 5986 28800
rect 15118 28864 15434 28865
rect 15118 28800 15124 28864
rect 15188 28800 15204 28864
rect 15268 28800 15284 28864
rect 15348 28800 15364 28864
rect 15428 28800 15434 28864
rect 15118 28799 15434 28800
rect 24566 28864 24882 28865
rect 24566 28800 24572 28864
rect 24636 28800 24652 28864
rect 24716 28800 24732 28864
rect 24796 28800 24812 28864
rect 24876 28800 24882 28864
rect 24566 28799 24882 28800
rect 34014 28864 34330 28865
rect 34014 28800 34020 28864
rect 34084 28800 34100 28864
rect 34164 28800 34180 28864
rect 34244 28800 34260 28864
rect 34324 28800 34330 28864
rect 34014 28799 34330 28800
rect 10394 28320 10710 28321
rect 10394 28256 10400 28320
rect 10464 28256 10480 28320
rect 10544 28256 10560 28320
rect 10624 28256 10640 28320
rect 10704 28256 10710 28320
rect 10394 28255 10710 28256
rect 19842 28320 20158 28321
rect 19842 28256 19848 28320
rect 19912 28256 19928 28320
rect 19992 28256 20008 28320
rect 20072 28256 20088 28320
rect 20152 28256 20158 28320
rect 19842 28255 20158 28256
rect 29290 28320 29606 28321
rect 29290 28256 29296 28320
rect 29360 28256 29376 28320
rect 29440 28256 29456 28320
rect 29520 28256 29536 28320
rect 29600 28256 29606 28320
rect 29290 28255 29606 28256
rect 5670 27776 5986 27777
rect 5670 27712 5676 27776
rect 5740 27712 5756 27776
rect 5820 27712 5836 27776
rect 5900 27712 5916 27776
rect 5980 27712 5986 27776
rect 5670 27711 5986 27712
rect 15118 27776 15434 27777
rect 15118 27712 15124 27776
rect 15188 27712 15204 27776
rect 15268 27712 15284 27776
rect 15348 27712 15364 27776
rect 15428 27712 15434 27776
rect 15118 27711 15434 27712
rect 24566 27776 24882 27777
rect 24566 27712 24572 27776
rect 24636 27712 24652 27776
rect 24716 27712 24732 27776
rect 24796 27712 24812 27776
rect 24876 27712 24882 27776
rect 24566 27711 24882 27712
rect 34014 27776 34330 27777
rect 34014 27712 34020 27776
rect 34084 27712 34100 27776
rect 34164 27712 34180 27776
rect 34244 27712 34260 27776
rect 34324 27712 34330 27776
rect 34014 27711 34330 27712
rect 0 27570 800 27600
rect 1485 27570 1551 27573
rect 0 27568 1551 27570
rect 0 27512 1490 27568
rect 1546 27512 1551 27568
rect 0 27510 1551 27512
rect 0 27480 800 27510
rect 1485 27507 1551 27510
rect 10394 27232 10710 27233
rect 10394 27168 10400 27232
rect 10464 27168 10480 27232
rect 10544 27168 10560 27232
rect 10624 27168 10640 27232
rect 10704 27168 10710 27232
rect 10394 27167 10710 27168
rect 19842 27232 20158 27233
rect 19842 27168 19848 27232
rect 19912 27168 19928 27232
rect 19992 27168 20008 27232
rect 20072 27168 20088 27232
rect 20152 27168 20158 27232
rect 19842 27167 20158 27168
rect 29290 27232 29606 27233
rect 29290 27168 29296 27232
rect 29360 27168 29376 27232
rect 29440 27168 29456 27232
rect 29520 27168 29536 27232
rect 29600 27168 29606 27232
rect 29290 27167 29606 27168
rect 5670 26688 5986 26689
rect 5670 26624 5676 26688
rect 5740 26624 5756 26688
rect 5820 26624 5836 26688
rect 5900 26624 5916 26688
rect 5980 26624 5986 26688
rect 5670 26623 5986 26624
rect 15118 26688 15434 26689
rect 15118 26624 15124 26688
rect 15188 26624 15204 26688
rect 15268 26624 15284 26688
rect 15348 26624 15364 26688
rect 15428 26624 15434 26688
rect 15118 26623 15434 26624
rect 24566 26688 24882 26689
rect 24566 26624 24572 26688
rect 24636 26624 24652 26688
rect 24716 26624 24732 26688
rect 24796 26624 24812 26688
rect 24876 26624 24882 26688
rect 24566 26623 24882 26624
rect 34014 26688 34330 26689
rect 34014 26624 34020 26688
rect 34084 26624 34100 26688
rect 34164 26624 34180 26688
rect 34244 26624 34260 26688
rect 34324 26624 34330 26688
rect 34014 26623 34330 26624
rect 0 26210 800 26240
rect 1485 26210 1551 26213
rect 0 26208 1551 26210
rect 0 26152 1490 26208
rect 1546 26152 1551 26208
rect 0 26150 1551 26152
rect 0 26120 800 26150
rect 1485 26147 1551 26150
rect 10394 26144 10710 26145
rect 10394 26080 10400 26144
rect 10464 26080 10480 26144
rect 10544 26080 10560 26144
rect 10624 26080 10640 26144
rect 10704 26080 10710 26144
rect 10394 26079 10710 26080
rect 19842 26144 20158 26145
rect 19842 26080 19848 26144
rect 19912 26080 19928 26144
rect 19992 26080 20008 26144
rect 20072 26080 20088 26144
rect 20152 26080 20158 26144
rect 19842 26079 20158 26080
rect 29290 26144 29606 26145
rect 29290 26080 29296 26144
rect 29360 26080 29376 26144
rect 29440 26080 29456 26144
rect 29520 26080 29536 26144
rect 29600 26080 29606 26144
rect 29290 26079 29606 26080
rect 5670 25600 5986 25601
rect 5670 25536 5676 25600
rect 5740 25536 5756 25600
rect 5820 25536 5836 25600
rect 5900 25536 5916 25600
rect 5980 25536 5986 25600
rect 5670 25535 5986 25536
rect 15118 25600 15434 25601
rect 15118 25536 15124 25600
rect 15188 25536 15204 25600
rect 15268 25536 15284 25600
rect 15348 25536 15364 25600
rect 15428 25536 15434 25600
rect 15118 25535 15434 25536
rect 24566 25600 24882 25601
rect 24566 25536 24572 25600
rect 24636 25536 24652 25600
rect 24716 25536 24732 25600
rect 24796 25536 24812 25600
rect 24876 25536 24882 25600
rect 24566 25535 24882 25536
rect 34014 25600 34330 25601
rect 34014 25536 34020 25600
rect 34084 25536 34100 25600
rect 34164 25536 34180 25600
rect 34244 25536 34260 25600
rect 34324 25536 34330 25600
rect 34014 25535 34330 25536
rect 10394 25056 10710 25057
rect 10394 24992 10400 25056
rect 10464 24992 10480 25056
rect 10544 24992 10560 25056
rect 10624 24992 10640 25056
rect 10704 24992 10710 25056
rect 10394 24991 10710 24992
rect 19842 25056 20158 25057
rect 19842 24992 19848 25056
rect 19912 24992 19928 25056
rect 19992 24992 20008 25056
rect 20072 24992 20088 25056
rect 20152 24992 20158 25056
rect 19842 24991 20158 24992
rect 29290 25056 29606 25057
rect 29290 24992 29296 25056
rect 29360 24992 29376 25056
rect 29440 24992 29456 25056
rect 29520 24992 29536 25056
rect 29600 24992 29606 25056
rect 29290 24991 29606 24992
rect 0 24850 800 24880
rect 1485 24850 1551 24853
rect 0 24848 1551 24850
rect 0 24792 1490 24848
rect 1546 24792 1551 24848
rect 0 24790 1551 24792
rect 0 24760 800 24790
rect 1485 24787 1551 24790
rect 5670 24512 5986 24513
rect 5670 24448 5676 24512
rect 5740 24448 5756 24512
rect 5820 24448 5836 24512
rect 5900 24448 5916 24512
rect 5980 24448 5986 24512
rect 5670 24447 5986 24448
rect 15118 24512 15434 24513
rect 15118 24448 15124 24512
rect 15188 24448 15204 24512
rect 15268 24448 15284 24512
rect 15348 24448 15364 24512
rect 15428 24448 15434 24512
rect 15118 24447 15434 24448
rect 24566 24512 24882 24513
rect 24566 24448 24572 24512
rect 24636 24448 24652 24512
rect 24716 24448 24732 24512
rect 24796 24448 24812 24512
rect 24876 24448 24882 24512
rect 24566 24447 24882 24448
rect 34014 24512 34330 24513
rect 34014 24448 34020 24512
rect 34084 24448 34100 24512
rect 34164 24448 34180 24512
rect 34244 24448 34260 24512
rect 34324 24448 34330 24512
rect 34014 24447 34330 24448
rect 10394 23968 10710 23969
rect 10394 23904 10400 23968
rect 10464 23904 10480 23968
rect 10544 23904 10560 23968
rect 10624 23904 10640 23968
rect 10704 23904 10710 23968
rect 10394 23903 10710 23904
rect 19842 23968 20158 23969
rect 19842 23904 19848 23968
rect 19912 23904 19928 23968
rect 19992 23904 20008 23968
rect 20072 23904 20088 23968
rect 20152 23904 20158 23968
rect 19842 23903 20158 23904
rect 29290 23968 29606 23969
rect 29290 23904 29296 23968
rect 29360 23904 29376 23968
rect 29440 23904 29456 23968
rect 29520 23904 29536 23968
rect 29600 23904 29606 23968
rect 29290 23903 29606 23904
rect 0 23490 800 23520
rect 1485 23490 1551 23493
rect 0 23488 1551 23490
rect 0 23432 1490 23488
rect 1546 23432 1551 23488
rect 0 23430 1551 23432
rect 0 23400 800 23430
rect 1485 23427 1551 23430
rect 5670 23424 5986 23425
rect 5670 23360 5676 23424
rect 5740 23360 5756 23424
rect 5820 23360 5836 23424
rect 5900 23360 5916 23424
rect 5980 23360 5986 23424
rect 5670 23359 5986 23360
rect 15118 23424 15434 23425
rect 15118 23360 15124 23424
rect 15188 23360 15204 23424
rect 15268 23360 15284 23424
rect 15348 23360 15364 23424
rect 15428 23360 15434 23424
rect 15118 23359 15434 23360
rect 24566 23424 24882 23425
rect 24566 23360 24572 23424
rect 24636 23360 24652 23424
rect 24716 23360 24732 23424
rect 24796 23360 24812 23424
rect 24876 23360 24882 23424
rect 24566 23359 24882 23360
rect 34014 23424 34330 23425
rect 34014 23360 34020 23424
rect 34084 23360 34100 23424
rect 34164 23360 34180 23424
rect 34244 23360 34260 23424
rect 34324 23360 34330 23424
rect 34014 23359 34330 23360
rect 10394 22880 10710 22881
rect 10394 22816 10400 22880
rect 10464 22816 10480 22880
rect 10544 22816 10560 22880
rect 10624 22816 10640 22880
rect 10704 22816 10710 22880
rect 10394 22815 10710 22816
rect 19842 22880 20158 22881
rect 19842 22816 19848 22880
rect 19912 22816 19928 22880
rect 19992 22816 20008 22880
rect 20072 22816 20088 22880
rect 20152 22816 20158 22880
rect 19842 22815 20158 22816
rect 29290 22880 29606 22881
rect 29290 22816 29296 22880
rect 29360 22816 29376 22880
rect 29440 22816 29456 22880
rect 29520 22816 29536 22880
rect 29600 22816 29606 22880
rect 29290 22815 29606 22816
rect 5670 22336 5986 22337
rect 5670 22272 5676 22336
rect 5740 22272 5756 22336
rect 5820 22272 5836 22336
rect 5900 22272 5916 22336
rect 5980 22272 5986 22336
rect 5670 22271 5986 22272
rect 15118 22336 15434 22337
rect 15118 22272 15124 22336
rect 15188 22272 15204 22336
rect 15268 22272 15284 22336
rect 15348 22272 15364 22336
rect 15428 22272 15434 22336
rect 15118 22271 15434 22272
rect 24566 22336 24882 22337
rect 24566 22272 24572 22336
rect 24636 22272 24652 22336
rect 24716 22272 24732 22336
rect 24796 22272 24812 22336
rect 24876 22272 24882 22336
rect 24566 22271 24882 22272
rect 34014 22336 34330 22337
rect 34014 22272 34020 22336
rect 34084 22272 34100 22336
rect 34164 22272 34180 22336
rect 34244 22272 34260 22336
rect 34324 22272 34330 22336
rect 34014 22271 34330 22272
rect 0 22130 800 22160
rect 1393 22130 1459 22133
rect 0 22128 1459 22130
rect 0 22072 1398 22128
rect 1454 22072 1459 22128
rect 0 22070 1459 22072
rect 0 22040 800 22070
rect 1393 22067 1459 22070
rect 10394 21792 10710 21793
rect 10394 21728 10400 21792
rect 10464 21728 10480 21792
rect 10544 21728 10560 21792
rect 10624 21728 10640 21792
rect 10704 21728 10710 21792
rect 10394 21727 10710 21728
rect 19842 21792 20158 21793
rect 19842 21728 19848 21792
rect 19912 21728 19928 21792
rect 19992 21728 20008 21792
rect 20072 21728 20088 21792
rect 20152 21728 20158 21792
rect 19842 21727 20158 21728
rect 29290 21792 29606 21793
rect 29290 21728 29296 21792
rect 29360 21728 29376 21792
rect 29440 21728 29456 21792
rect 29520 21728 29536 21792
rect 29600 21728 29606 21792
rect 29290 21727 29606 21728
rect 5670 21248 5986 21249
rect 5670 21184 5676 21248
rect 5740 21184 5756 21248
rect 5820 21184 5836 21248
rect 5900 21184 5916 21248
rect 5980 21184 5986 21248
rect 5670 21183 5986 21184
rect 15118 21248 15434 21249
rect 15118 21184 15124 21248
rect 15188 21184 15204 21248
rect 15268 21184 15284 21248
rect 15348 21184 15364 21248
rect 15428 21184 15434 21248
rect 15118 21183 15434 21184
rect 24566 21248 24882 21249
rect 24566 21184 24572 21248
rect 24636 21184 24652 21248
rect 24716 21184 24732 21248
rect 24796 21184 24812 21248
rect 24876 21184 24882 21248
rect 24566 21183 24882 21184
rect 34014 21248 34330 21249
rect 34014 21184 34020 21248
rect 34084 21184 34100 21248
rect 34164 21184 34180 21248
rect 34244 21184 34260 21248
rect 34324 21184 34330 21248
rect 34014 21183 34330 21184
rect 0 20770 800 20800
rect 1485 20770 1551 20773
rect 0 20768 1551 20770
rect 0 20712 1490 20768
rect 1546 20712 1551 20768
rect 0 20710 1551 20712
rect 0 20680 800 20710
rect 1485 20707 1551 20710
rect 10394 20704 10710 20705
rect 10394 20640 10400 20704
rect 10464 20640 10480 20704
rect 10544 20640 10560 20704
rect 10624 20640 10640 20704
rect 10704 20640 10710 20704
rect 10394 20639 10710 20640
rect 19842 20704 20158 20705
rect 19842 20640 19848 20704
rect 19912 20640 19928 20704
rect 19992 20640 20008 20704
rect 20072 20640 20088 20704
rect 20152 20640 20158 20704
rect 19842 20639 20158 20640
rect 29290 20704 29606 20705
rect 29290 20640 29296 20704
rect 29360 20640 29376 20704
rect 29440 20640 29456 20704
rect 29520 20640 29536 20704
rect 29600 20640 29606 20704
rect 29290 20639 29606 20640
rect 5670 20160 5986 20161
rect 5670 20096 5676 20160
rect 5740 20096 5756 20160
rect 5820 20096 5836 20160
rect 5900 20096 5916 20160
rect 5980 20096 5986 20160
rect 5670 20095 5986 20096
rect 15118 20160 15434 20161
rect 15118 20096 15124 20160
rect 15188 20096 15204 20160
rect 15268 20096 15284 20160
rect 15348 20096 15364 20160
rect 15428 20096 15434 20160
rect 15118 20095 15434 20096
rect 24566 20160 24882 20161
rect 24566 20096 24572 20160
rect 24636 20096 24652 20160
rect 24716 20096 24732 20160
rect 24796 20096 24812 20160
rect 24876 20096 24882 20160
rect 24566 20095 24882 20096
rect 34014 20160 34330 20161
rect 34014 20096 34020 20160
rect 34084 20096 34100 20160
rect 34164 20096 34180 20160
rect 34244 20096 34260 20160
rect 34324 20096 34330 20160
rect 34014 20095 34330 20096
rect 10394 19616 10710 19617
rect 10394 19552 10400 19616
rect 10464 19552 10480 19616
rect 10544 19552 10560 19616
rect 10624 19552 10640 19616
rect 10704 19552 10710 19616
rect 10394 19551 10710 19552
rect 19842 19616 20158 19617
rect 19842 19552 19848 19616
rect 19912 19552 19928 19616
rect 19992 19552 20008 19616
rect 20072 19552 20088 19616
rect 20152 19552 20158 19616
rect 19842 19551 20158 19552
rect 29290 19616 29606 19617
rect 29290 19552 29296 19616
rect 29360 19552 29376 19616
rect 29440 19552 29456 19616
rect 29520 19552 29536 19616
rect 29600 19552 29606 19616
rect 29290 19551 29606 19552
rect 0 19410 800 19440
rect 1485 19410 1551 19413
rect 0 19408 1551 19410
rect 0 19352 1490 19408
rect 1546 19352 1551 19408
rect 0 19350 1551 19352
rect 0 19320 800 19350
rect 1485 19347 1551 19350
rect 5670 19072 5986 19073
rect 5670 19008 5676 19072
rect 5740 19008 5756 19072
rect 5820 19008 5836 19072
rect 5900 19008 5916 19072
rect 5980 19008 5986 19072
rect 5670 19007 5986 19008
rect 15118 19072 15434 19073
rect 15118 19008 15124 19072
rect 15188 19008 15204 19072
rect 15268 19008 15284 19072
rect 15348 19008 15364 19072
rect 15428 19008 15434 19072
rect 15118 19007 15434 19008
rect 24566 19072 24882 19073
rect 24566 19008 24572 19072
rect 24636 19008 24652 19072
rect 24716 19008 24732 19072
rect 24796 19008 24812 19072
rect 24876 19008 24882 19072
rect 24566 19007 24882 19008
rect 34014 19072 34330 19073
rect 34014 19008 34020 19072
rect 34084 19008 34100 19072
rect 34164 19008 34180 19072
rect 34244 19008 34260 19072
rect 34324 19008 34330 19072
rect 34014 19007 34330 19008
rect 10394 18528 10710 18529
rect 10394 18464 10400 18528
rect 10464 18464 10480 18528
rect 10544 18464 10560 18528
rect 10624 18464 10640 18528
rect 10704 18464 10710 18528
rect 10394 18463 10710 18464
rect 19842 18528 20158 18529
rect 19842 18464 19848 18528
rect 19912 18464 19928 18528
rect 19992 18464 20008 18528
rect 20072 18464 20088 18528
rect 20152 18464 20158 18528
rect 19842 18463 20158 18464
rect 29290 18528 29606 18529
rect 29290 18464 29296 18528
rect 29360 18464 29376 18528
rect 29440 18464 29456 18528
rect 29520 18464 29536 18528
rect 29600 18464 29606 18528
rect 29290 18463 29606 18464
rect 0 18050 800 18080
rect 1485 18050 1551 18053
rect 0 18048 1551 18050
rect 0 17992 1490 18048
rect 1546 17992 1551 18048
rect 0 17990 1551 17992
rect 0 17960 800 17990
rect 1485 17987 1551 17990
rect 5670 17984 5986 17985
rect 5670 17920 5676 17984
rect 5740 17920 5756 17984
rect 5820 17920 5836 17984
rect 5900 17920 5916 17984
rect 5980 17920 5986 17984
rect 5670 17919 5986 17920
rect 15118 17984 15434 17985
rect 15118 17920 15124 17984
rect 15188 17920 15204 17984
rect 15268 17920 15284 17984
rect 15348 17920 15364 17984
rect 15428 17920 15434 17984
rect 15118 17919 15434 17920
rect 24566 17984 24882 17985
rect 24566 17920 24572 17984
rect 24636 17920 24652 17984
rect 24716 17920 24732 17984
rect 24796 17920 24812 17984
rect 24876 17920 24882 17984
rect 24566 17919 24882 17920
rect 34014 17984 34330 17985
rect 34014 17920 34020 17984
rect 34084 17920 34100 17984
rect 34164 17920 34180 17984
rect 34244 17920 34260 17984
rect 34324 17920 34330 17984
rect 34014 17919 34330 17920
rect 10394 17440 10710 17441
rect 10394 17376 10400 17440
rect 10464 17376 10480 17440
rect 10544 17376 10560 17440
rect 10624 17376 10640 17440
rect 10704 17376 10710 17440
rect 10394 17375 10710 17376
rect 19842 17440 20158 17441
rect 19842 17376 19848 17440
rect 19912 17376 19928 17440
rect 19992 17376 20008 17440
rect 20072 17376 20088 17440
rect 20152 17376 20158 17440
rect 19842 17375 20158 17376
rect 29290 17440 29606 17441
rect 29290 17376 29296 17440
rect 29360 17376 29376 17440
rect 29440 17376 29456 17440
rect 29520 17376 29536 17440
rect 29600 17376 29606 17440
rect 29290 17375 29606 17376
rect 5670 16896 5986 16897
rect 5670 16832 5676 16896
rect 5740 16832 5756 16896
rect 5820 16832 5836 16896
rect 5900 16832 5916 16896
rect 5980 16832 5986 16896
rect 5670 16831 5986 16832
rect 15118 16896 15434 16897
rect 15118 16832 15124 16896
rect 15188 16832 15204 16896
rect 15268 16832 15284 16896
rect 15348 16832 15364 16896
rect 15428 16832 15434 16896
rect 15118 16831 15434 16832
rect 24566 16896 24882 16897
rect 24566 16832 24572 16896
rect 24636 16832 24652 16896
rect 24716 16832 24732 16896
rect 24796 16832 24812 16896
rect 24876 16832 24882 16896
rect 24566 16831 24882 16832
rect 34014 16896 34330 16897
rect 34014 16832 34020 16896
rect 34084 16832 34100 16896
rect 34164 16832 34180 16896
rect 34244 16832 34260 16896
rect 34324 16832 34330 16896
rect 34014 16831 34330 16832
rect 0 16690 800 16720
rect 1485 16690 1551 16693
rect 0 16688 1551 16690
rect 0 16632 1490 16688
rect 1546 16632 1551 16688
rect 0 16630 1551 16632
rect 0 16600 800 16630
rect 1485 16627 1551 16630
rect 10394 16352 10710 16353
rect 10394 16288 10400 16352
rect 10464 16288 10480 16352
rect 10544 16288 10560 16352
rect 10624 16288 10640 16352
rect 10704 16288 10710 16352
rect 10394 16287 10710 16288
rect 19842 16352 20158 16353
rect 19842 16288 19848 16352
rect 19912 16288 19928 16352
rect 19992 16288 20008 16352
rect 20072 16288 20088 16352
rect 20152 16288 20158 16352
rect 19842 16287 20158 16288
rect 29290 16352 29606 16353
rect 29290 16288 29296 16352
rect 29360 16288 29376 16352
rect 29440 16288 29456 16352
rect 29520 16288 29536 16352
rect 29600 16288 29606 16352
rect 29290 16287 29606 16288
rect 5670 15808 5986 15809
rect 5670 15744 5676 15808
rect 5740 15744 5756 15808
rect 5820 15744 5836 15808
rect 5900 15744 5916 15808
rect 5980 15744 5986 15808
rect 5670 15743 5986 15744
rect 15118 15808 15434 15809
rect 15118 15744 15124 15808
rect 15188 15744 15204 15808
rect 15268 15744 15284 15808
rect 15348 15744 15364 15808
rect 15428 15744 15434 15808
rect 15118 15743 15434 15744
rect 24566 15808 24882 15809
rect 24566 15744 24572 15808
rect 24636 15744 24652 15808
rect 24716 15744 24732 15808
rect 24796 15744 24812 15808
rect 24876 15744 24882 15808
rect 24566 15743 24882 15744
rect 34014 15808 34330 15809
rect 34014 15744 34020 15808
rect 34084 15744 34100 15808
rect 34164 15744 34180 15808
rect 34244 15744 34260 15808
rect 34324 15744 34330 15808
rect 34014 15743 34330 15744
rect 0 15330 800 15360
rect 1485 15330 1551 15333
rect 0 15328 1551 15330
rect 0 15272 1490 15328
rect 1546 15272 1551 15328
rect 0 15270 1551 15272
rect 0 15240 800 15270
rect 1485 15267 1551 15270
rect 10394 15264 10710 15265
rect 10394 15200 10400 15264
rect 10464 15200 10480 15264
rect 10544 15200 10560 15264
rect 10624 15200 10640 15264
rect 10704 15200 10710 15264
rect 10394 15199 10710 15200
rect 19842 15264 20158 15265
rect 19842 15200 19848 15264
rect 19912 15200 19928 15264
rect 19992 15200 20008 15264
rect 20072 15200 20088 15264
rect 20152 15200 20158 15264
rect 19842 15199 20158 15200
rect 29290 15264 29606 15265
rect 29290 15200 29296 15264
rect 29360 15200 29376 15264
rect 29440 15200 29456 15264
rect 29520 15200 29536 15264
rect 29600 15200 29606 15264
rect 29290 15199 29606 15200
rect 5670 14720 5986 14721
rect 5670 14656 5676 14720
rect 5740 14656 5756 14720
rect 5820 14656 5836 14720
rect 5900 14656 5916 14720
rect 5980 14656 5986 14720
rect 5670 14655 5986 14656
rect 15118 14720 15434 14721
rect 15118 14656 15124 14720
rect 15188 14656 15204 14720
rect 15268 14656 15284 14720
rect 15348 14656 15364 14720
rect 15428 14656 15434 14720
rect 15118 14655 15434 14656
rect 24566 14720 24882 14721
rect 24566 14656 24572 14720
rect 24636 14656 24652 14720
rect 24716 14656 24732 14720
rect 24796 14656 24812 14720
rect 24876 14656 24882 14720
rect 24566 14655 24882 14656
rect 34014 14720 34330 14721
rect 34014 14656 34020 14720
rect 34084 14656 34100 14720
rect 34164 14656 34180 14720
rect 34244 14656 34260 14720
rect 34324 14656 34330 14720
rect 34014 14655 34330 14656
rect 10394 14176 10710 14177
rect 10394 14112 10400 14176
rect 10464 14112 10480 14176
rect 10544 14112 10560 14176
rect 10624 14112 10640 14176
rect 10704 14112 10710 14176
rect 10394 14111 10710 14112
rect 19842 14176 20158 14177
rect 19842 14112 19848 14176
rect 19912 14112 19928 14176
rect 19992 14112 20008 14176
rect 20072 14112 20088 14176
rect 20152 14112 20158 14176
rect 19842 14111 20158 14112
rect 29290 14176 29606 14177
rect 29290 14112 29296 14176
rect 29360 14112 29376 14176
rect 29440 14112 29456 14176
rect 29520 14112 29536 14176
rect 29600 14112 29606 14176
rect 29290 14111 29606 14112
rect 0 13970 800 14000
rect 1485 13970 1551 13973
rect 0 13968 1551 13970
rect 0 13912 1490 13968
rect 1546 13912 1551 13968
rect 0 13910 1551 13912
rect 0 13880 800 13910
rect 1485 13907 1551 13910
rect 5670 13632 5986 13633
rect 5670 13568 5676 13632
rect 5740 13568 5756 13632
rect 5820 13568 5836 13632
rect 5900 13568 5916 13632
rect 5980 13568 5986 13632
rect 5670 13567 5986 13568
rect 15118 13632 15434 13633
rect 15118 13568 15124 13632
rect 15188 13568 15204 13632
rect 15268 13568 15284 13632
rect 15348 13568 15364 13632
rect 15428 13568 15434 13632
rect 15118 13567 15434 13568
rect 24566 13632 24882 13633
rect 24566 13568 24572 13632
rect 24636 13568 24652 13632
rect 24716 13568 24732 13632
rect 24796 13568 24812 13632
rect 24876 13568 24882 13632
rect 24566 13567 24882 13568
rect 34014 13632 34330 13633
rect 34014 13568 34020 13632
rect 34084 13568 34100 13632
rect 34164 13568 34180 13632
rect 34244 13568 34260 13632
rect 34324 13568 34330 13632
rect 34014 13567 34330 13568
rect 10394 13088 10710 13089
rect 10394 13024 10400 13088
rect 10464 13024 10480 13088
rect 10544 13024 10560 13088
rect 10624 13024 10640 13088
rect 10704 13024 10710 13088
rect 10394 13023 10710 13024
rect 19842 13088 20158 13089
rect 19842 13024 19848 13088
rect 19912 13024 19928 13088
rect 19992 13024 20008 13088
rect 20072 13024 20088 13088
rect 20152 13024 20158 13088
rect 19842 13023 20158 13024
rect 29290 13088 29606 13089
rect 29290 13024 29296 13088
rect 29360 13024 29376 13088
rect 29440 13024 29456 13088
rect 29520 13024 29536 13088
rect 29600 13024 29606 13088
rect 29290 13023 29606 13024
rect 0 12610 800 12640
rect 1485 12610 1551 12613
rect 0 12608 1551 12610
rect 0 12552 1490 12608
rect 1546 12552 1551 12608
rect 0 12550 1551 12552
rect 0 12520 800 12550
rect 1485 12547 1551 12550
rect 5670 12544 5986 12545
rect 5670 12480 5676 12544
rect 5740 12480 5756 12544
rect 5820 12480 5836 12544
rect 5900 12480 5916 12544
rect 5980 12480 5986 12544
rect 5670 12479 5986 12480
rect 15118 12544 15434 12545
rect 15118 12480 15124 12544
rect 15188 12480 15204 12544
rect 15268 12480 15284 12544
rect 15348 12480 15364 12544
rect 15428 12480 15434 12544
rect 15118 12479 15434 12480
rect 24566 12544 24882 12545
rect 24566 12480 24572 12544
rect 24636 12480 24652 12544
rect 24716 12480 24732 12544
rect 24796 12480 24812 12544
rect 24876 12480 24882 12544
rect 24566 12479 24882 12480
rect 34014 12544 34330 12545
rect 34014 12480 34020 12544
rect 34084 12480 34100 12544
rect 34164 12480 34180 12544
rect 34244 12480 34260 12544
rect 34324 12480 34330 12544
rect 34014 12479 34330 12480
rect 10394 12000 10710 12001
rect 10394 11936 10400 12000
rect 10464 11936 10480 12000
rect 10544 11936 10560 12000
rect 10624 11936 10640 12000
rect 10704 11936 10710 12000
rect 10394 11935 10710 11936
rect 19842 12000 20158 12001
rect 19842 11936 19848 12000
rect 19912 11936 19928 12000
rect 19992 11936 20008 12000
rect 20072 11936 20088 12000
rect 20152 11936 20158 12000
rect 19842 11935 20158 11936
rect 29290 12000 29606 12001
rect 29290 11936 29296 12000
rect 29360 11936 29376 12000
rect 29440 11936 29456 12000
rect 29520 11936 29536 12000
rect 29600 11936 29606 12000
rect 29290 11935 29606 11936
rect 5670 11456 5986 11457
rect 5670 11392 5676 11456
rect 5740 11392 5756 11456
rect 5820 11392 5836 11456
rect 5900 11392 5916 11456
rect 5980 11392 5986 11456
rect 5670 11391 5986 11392
rect 15118 11456 15434 11457
rect 15118 11392 15124 11456
rect 15188 11392 15204 11456
rect 15268 11392 15284 11456
rect 15348 11392 15364 11456
rect 15428 11392 15434 11456
rect 15118 11391 15434 11392
rect 24566 11456 24882 11457
rect 24566 11392 24572 11456
rect 24636 11392 24652 11456
rect 24716 11392 24732 11456
rect 24796 11392 24812 11456
rect 24876 11392 24882 11456
rect 24566 11391 24882 11392
rect 34014 11456 34330 11457
rect 34014 11392 34020 11456
rect 34084 11392 34100 11456
rect 34164 11392 34180 11456
rect 34244 11392 34260 11456
rect 34324 11392 34330 11456
rect 34014 11391 34330 11392
rect 0 11250 800 11280
rect 1485 11250 1551 11253
rect 0 11248 1551 11250
rect 0 11192 1490 11248
rect 1546 11192 1551 11248
rect 0 11190 1551 11192
rect 0 11160 800 11190
rect 1485 11187 1551 11190
rect 10394 10912 10710 10913
rect 10394 10848 10400 10912
rect 10464 10848 10480 10912
rect 10544 10848 10560 10912
rect 10624 10848 10640 10912
rect 10704 10848 10710 10912
rect 10394 10847 10710 10848
rect 19842 10912 20158 10913
rect 19842 10848 19848 10912
rect 19912 10848 19928 10912
rect 19992 10848 20008 10912
rect 20072 10848 20088 10912
rect 20152 10848 20158 10912
rect 19842 10847 20158 10848
rect 29290 10912 29606 10913
rect 29290 10848 29296 10912
rect 29360 10848 29376 10912
rect 29440 10848 29456 10912
rect 29520 10848 29536 10912
rect 29600 10848 29606 10912
rect 29290 10847 29606 10848
rect 5670 10368 5986 10369
rect 5670 10304 5676 10368
rect 5740 10304 5756 10368
rect 5820 10304 5836 10368
rect 5900 10304 5916 10368
rect 5980 10304 5986 10368
rect 5670 10303 5986 10304
rect 15118 10368 15434 10369
rect 15118 10304 15124 10368
rect 15188 10304 15204 10368
rect 15268 10304 15284 10368
rect 15348 10304 15364 10368
rect 15428 10304 15434 10368
rect 15118 10303 15434 10304
rect 24566 10368 24882 10369
rect 24566 10304 24572 10368
rect 24636 10304 24652 10368
rect 24716 10304 24732 10368
rect 24796 10304 24812 10368
rect 24876 10304 24882 10368
rect 24566 10303 24882 10304
rect 34014 10368 34330 10369
rect 34014 10304 34020 10368
rect 34084 10304 34100 10368
rect 34164 10304 34180 10368
rect 34244 10304 34260 10368
rect 34324 10304 34330 10368
rect 34014 10303 34330 10304
rect 0 9890 800 9920
rect 1485 9890 1551 9893
rect 0 9888 1551 9890
rect 0 9832 1490 9888
rect 1546 9832 1551 9888
rect 0 9830 1551 9832
rect 0 9800 800 9830
rect 1485 9827 1551 9830
rect 10394 9824 10710 9825
rect 10394 9760 10400 9824
rect 10464 9760 10480 9824
rect 10544 9760 10560 9824
rect 10624 9760 10640 9824
rect 10704 9760 10710 9824
rect 10394 9759 10710 9760
rect 19842 9824 20158 9825
rect 19842 9760 19848 9824
rect 19912 9760 19928 9824
rect 19992 9760 20008 9824
rect 20072 9760 20088 9824
rect 20152 9760 20158 9824
rect 19842 9759 20158 9760
rect 29290 9824 29606 9825
rect 29290 9760 29296 9824
rect 29360 9760 29376 9824
rect 29440 9760 29456 9824
rect 29520 9760 29536 9824
rect 29600 9760 29606 9824
rect 29290 9759 29606 9760
rect 5670 9280 5986 9281
rect 5670 9216 5676 9280
rect 5740 9216 5756 9280
rect 5820 9216 5836 9280
rect 5900 9216 5916 9280
rect 5980 9216 5986 9280
rect 5670 9215 5986 9216
rect 15118 9280 15434 9281
rect 15118 9216 15124 9280
rect 15188 9216 15204 9280
rect 15268 9216 15284 9280
rect 15348 9216 15364 9280
rect 15428 9216 15434 9280
rect 15118 9215 15434 9216
rect 24566 9280 24882 9281
rect 24566 9216 24572 9280
rect 24636 9216 24652 9280
rect 24716 9216 24732 9280
rect 24796 9216 24812 9280
rect 24876 9216 24882 9280
rect 24566 9215 24882 9216
rect 34014 9280 34330 9281
rect 34014 9216 34020 9280
rect 34084 9216 34100 9280
rect 34164 9216 34180 9280
rect 34244 9216 34260 9280
rect 34324 9216 34330 9280
rect 34014 9215 34330 9216
rect 10394 8736 10710 8737
rect 10394 8672 10400 8736
rect 10464 8672 10480 8736
rect 10544 8672 10560 8736
rect 10624 8672 10640 8736
rect 10704 8672 10710 8736
rect 10394 8671 10710 8672
rect 19842 8736 20158 8737
rect 19842 8672 19848 8736
rect 19912 8672 19928 8736
rect 19992 8672 20008 8736
rect 20072 8672 20088 8736
rect 20152 8672 20158 8736
rect 19842 8671 20158 8672
rect 29290 8736 29606 8737
rect 29290 8672 29296 8736
rect 29360 8672 29376 8736
rect 29440 8672 29456 8736
rect 29520 8672 29536 8736
rect 29600 8672 29606 8736
rect 29290 8671 29606 8672
rect 0 8530 800 8560
rect 1485 8530 1551 8533
rect 0 8528 1551 8530
rect 0 8472 1490 8528
rect 1546 8472 1551 8528
rect 0 8470 1551 8472
rect 0 8440 800 8470
rect 1485 8467 1551 8470
rect 5670 8192 5986 8193
rect 5670 8128 5676 8192
rect 5740 8128 5756 8192
rect 5820 8128 5836 8192
rect 5900 8128 5916 8192
rect 5980 8128 5986 8192
rect 5670 8127 5986 8128
rect 15118 8192 15434 8193
rect 15118 8128 15124 8192
rect 15188 8128 15204 8192
rect 15268 8128 15284 8192
rect 15348 8128 15364 8192
rect 15428 8128 15434 8192
rect 15118 8127 15434 8128
rect 24566 8192 24882 8193
rect 24566 8128 24572 8192
rect 24636 8128 24652 8192
rect 24716 8128 24732 8192
rect 24796 8128 24812 8192
rect 24876 8128 24882 8192
rect 24566 8127 24882 8128
rect 34014 8192 34330 8193
rect 34014 8128 34020 8192
rect 34084 8128 34100 8192
rect 34164 8128 34180 8192
rect 34244 8128 34260 8192
rect 34324 8128 34330 8192
rect 34014 8127 34330 8128
rect 10394 7648 10710 7649
rect 10394 7584 10400 7648
rect 10464 7584 10480 7648
rect 10544 7584 10560 7648
rect 10624 7584 10640 7648
rect 10704 7584 10710 7648
rect 10394 7583 10710 7584
rect 19842 7648 20158 7649
rect 19842 7584 19848 7648
rect 19912 7584 19928 7648
rect 19992 7584 20008 7648
rect 20072 7584 20088 7648
rect 20152 7584 20158 7648
rect 19842 7583 20158 7584
rect 29290 7648 29606 7649
rect 29290 7584 29296 7648
rect 29360 7584 29376 7648
rect 29440 7584 29456 7648
rect 29520 7584 29536 7648
rect 29600 7584 29606 7648
rect 29290 7583 29606 7584
rect 0 7170 800 7200
rect 1485 7170 1551 7173
rect 0 7168 1551 7170
rect 0 7112 1490 7168
rect 1546 7112 1551 7168
rect 0 7110 1551 7112
rect 0 7080 800 7110
rect 1485 7107 1551 7110
rect 5670 7104 5986 7105
rect 5670 7040 5676 7104
rect 5740 7040 5756 7104
rect 5820 7040 5836 7104
rect 5900 7040 5916 7104
rect 5980 7040 5986 7104
rect 5670 7039 5986 7040
rect 15118 7104 15434 7105
rect 15118 7040 15124 7104
rect 15188 7040 15204 7104
rect 15268 7040 15284 7104
rect 15348 7040 15364 7104
rect 15428 7040 15434 7104
rect 15118 7039 15434 7040
rect 24566 7104 24882 7105
rect 24566 7040 24572 7104
rect 24636 7040 24652 7104
rect 24716 7040 24732 7104
rect 24796 7040 24812 7104
rect 24876 7040 24882 7104
rect 24566 7039 24882 7040
rect 34014 7104 34330 7105
rect 34014 7040 34020 7104
rect 34084 7040 34100 7104
rect 34164 7040 34180 7104
rect 34244 7040 34260 7104
rect 34324 7040 34330 7104
rect 34014 7039 34330 7040
rect 10394 6560 10710 6561
rect 10394 6496 10400 6560
rect 10464 6496 10480 6560
rect 10544 6496 10560 6560
rect 10624 6496 10640 6560
rect 10704 6496 10710 6560
rect 10394 6495 10710 6496
rect 19842 6560 20158 6561
rect 19842 6496 19848 6560
rect 19912 6496 19928 6560
rect 19992 6496 20008 6560
rect 20072 6496 20088 6560
rect 20152 6496 20158 6560
rect 19842 6495 20158 6496
rect 29290 6560 29606 6561
rect 29290 6496 29296 6560
rect 29360 6496 29376 6560
rect 29440 6496 29456 6560
rect 29520 6496 29536 6560
rect 29600 6496 29606 6560
rect 29290 6495 29606 6496
rect 5670 6016 5986 6017
rect 5670 5952 5676 6016
rect 5740 5952 5756 6016
rect 5820 5952 5836 6016
rect 5900 5952 5916 6016
rect 5980 5952 5986 6016
rect 5670 5951 5986 5952
rect 15118 6016 15434 6017
rect 15118 5952 15124 6016
rect 15188 5952 15204 6016
rect 15268 5952 15284 6016
rect 15348 5952 15364 6016
rect 15428 5952 15434 6016
rect 15118 5951 15434 5952
rect 24566 6016 24882 6017
rect 24566 5952 24572 6016
rect 24636 5952 24652 6016
rect 24716 5952 24732 6016
rect 24796 5952 24812 6016
rect 24876 5952 24882 6016
rect 24566 5951 24882 5952
rect 34014 6016 34330 6017
rect 34014 5952 34020 6016
rect 34084 5952 34100 6016
rect 34164 5952 34180 6016
rect 34244 5952 34260 6016
rect 34324 5952 34330 6016
rect 34014 5951 34330 5952
rect 0 5810 800 5840
rect 1485 5810 1551 5813
rect 0 5808 1551 5810
rect 0 5752 1490 5808
rect 1546 5752 1551 5808
rect 0 5750 1551 5752
rect 0 5720 800 5750
rect 1485 5747 1551 5750
rect 10394 5472 10710 5473
rect 10394 5408 10400 5472
rect 10464 5408 10480 5472
rect 10544 5408 10560 5472
rect 10624 5408 10640 5472
rect 10704 5408 10710 5472
rect 10394 5407 10710 5408
rect 19842 5472 20158 5473
rect 19842 5408 19848 5472
rect 19912 5408 19928 5472
rect 19992 5408 20008 5472
rect 20072 5408 20088 5472
rect 20152 5408 20158 5472
rect 19842 5407 20158 5408
rect 29290 5472 29606 5473
rect 29290 5408 29296 5472
rect 29360 5408 29376 5472
rect 29440 5408 29456 5472
rect 29520 5408 29536 5472
rect 29600 5408 29606 5472
rect 29290 5407 29606 5408
rect 5670 4928 5986 4929
rect 5670 4864 5676 4928
rect 5740 4864 5756 4928
rect 5820 4864 5836 4928
rect 5900 4864 5916 4928
rect 5980 4864 5986 4928
rect 5670 4863 5986 4864
rect 15118 4928 15434 4929
rect 15118 4864 15124 4928
rect 15188 4864 15204 4928
rect 15268 4864 15284 4928
rect 15348 4864 15364 4928
rect 15428 4864 15434 4928
rect 15118 4863 15434 4864
rect 24566 4928 24882 4929
rect 24566 4864 24572 4928
rect 24636 4864 24652 4928
rect 24716 4864 24732 4928
rect 24796 4864 24812 4928
rect 24876 4864 24882 4928
rect 24566 4863 24882 4864
rect 34014 4928 34330 4929
rect 34014 4864 34020 4928
rect 34084 4864 34100 4928
rect 34164 4864 34180 4928
rect 34244 4864 34260 4928
rect 34324 4864 34330 4928
rect 34014 4863 34330 4864
rect 0 4450 800 4480
rect 1485 4450 1551 4453
rect 0 4448 1551 4450
rect 0 4392 1490 4448
rect 1546 4392 1551 4448
rect 0 4390 1551 4392
rect 0 4360 800 4390
rect 1485 4387 1551 4390
rect 10394 4384 10710 4385
rect 10394 4320 10400 4384
rect 10464 4320 10480 4384
rect 10544 4320 10560 4384
rect 10624 4320 10640 4384
rect 10704 4320 10710 4384
rect 10394 4319 10710 4320
rect 19842 4384 20158 4385
rect 19842 4320 19848 4384
rect 19912 4320 19928 4384
rect 19992 4320 20008 4384
rect 20072 4320 20088 4384
rect 20152 4320 20158 4384
rect 19842 4319 20158 4320
rect 29290 4384 29606 4385
rect 29290 4320 29296 4384
rect 29360 4320 29376 4384
rect 29440 4320 29456 4384
rect 29520 4320 29536 4384
rect 29600 4320 29606 4384
rect 29290 4319 29606 4320
rect 5670 3840 5986 3841
rect 5670 3776 5676 3840
rect 5740 3776 5756 3840
rect 5820 3776 5836 3840
rect 5900 3776 5916 3840
rect 5980 3776 5986 3840
rect 5670 3775 5986 3776
rect 15118 3840 15434 3841
rect 15118 3776 15124 3840
rect 15188 3776 15204 3840
rect 15268 3776 15284 3840
rect 15348 3776 15364 3840
rect 15428 3776 15434 3840
rect 15118 3775 15434 3776
rect 24566 3840 24882 3841
rect 24566 3776 24572 3840
rect 24636 3776 24652 3840
rect 24716 3776 24732 3840
rect 24796 3776 24812 3840
rect 24876 3776 24882 3840
rect 24566 3775 24882 3776
rect 34014 3840 34330 3841
rect 34014 3776 34020 3840
rect 34084 3776 34100 3840
rect 34164 3776 34180 3840
rect 34244 3776 34260 3840
rect 34324 3776 34330 3840
rect 34014 3775 34330 3776
rect 10394 3296 10710 3297
rect 10394 3232 10400 3296
rect 10464 3232 10480 3296
rect 10544 3232 10560 3296
rect 10624 3232 10640 3296
rect 10704 3232 10710 3296
rect 10394 3231 10710 3232
rect 19842 3296 20158 3297
rect 19842 3232 19848 3296
rect 19912 3232 19928 3296
rect 19992 3232 20008 3296
rect 20072 3232 20088 3296
rect 20152 3232 20158 3296
rect 19842 3231 20158 3232
rect 29290 3296 29606 3297
rect 29290 3232 29296 3296
rect 29360 3232 29376 3296
rect 29440 3232 29456 3296
rect 29520 3232 29536 3296
rect 29600 3232 29606 3296
rect 29290 3231 29606 3232
rect 0 3090 800 3120
rect 1485 3090 1551 3093
rect 0 3088 1551 3090
rect 0 3032 1490 3088
rect 1546 3032 1551 3088
rect 0 3030 1551 3032
rect 0 3000 800 3030
rect 1485 3027 1551 3030
rect 5670 2752 5986 2753
rect 5670 2688 5676 2752
rect 5740 2688 5756 2752
rect 5820 2688 5836 2752
rect 5900 2688 5916 2752
rect 5980 2688 5986 2752
rect 5670 2687 5986 2688
rect 15118 2752 15434 2753
rect 15118 2688 15124 2752
rect 15188 2688 15204 2752
rect 15268 2688 15284 2752
rect 15348 2688 15364 2752
rect 15428 2688 15434 2752
rect 15118 2687 15434 2688
rect 24566 2752 24882 2753
rect 24566 2688 24572 2752
rect 24636 2688 24652 2752
rect 24716 2688 24732 2752
rect 24796 2688 24812 2752
rect 24876 2688 24882 2752
rect 24566 2687 24882 2688
rect 34014 2752 34330 2753
rect 34014 2688 34020 2752
rect 34084 2688 34100 2752
rect 34164 2688 34180 2752
rect 34244 2688 34260 2752
rect 34324 2688 34330 2752
rect 34014 2687 34330 2688
rect 10394 2208 10710 2209
rect 10394 2144 10400 2208
rect 10464 2144 10480 2208
rect 10544 2144 10560 2208
rect 10624 2144 10640 2208
rect 10704 2144 10710 2208
rect 10394 2143 10710 2144
rect 19842 2208 20158 2209
rect 19842 2144 19848 2208
rect 19912 2144 19928 2208
rect 19992 2144 20008 2208
rect 20072 2144 20088 2208
rect 20152 2144 20158 2208
rect 19842 2143 20158 2144
rect 29290 2208 29606 2209
rect 29290 2144 29296 2208
rect 29360 2144 29376 2208
rect 29440 2144 29456 2208
rect 29520 2144 29536 2208
rect 29600 2144 29606 2208
rect 29290 2143 29606 2144
rect 0 1730 800 1760
rect 1485 1730 1551 1733
rect 0 1728 1551 1730
rect 0 1672 1490 1728
rect 1546 1672 1551 1728
rect 0 1670 1551 1672
rect 0 1640 800 1670
rect 1485 1667 1551 1670
<< via3 >>
rect 10400 33756 10464 33760
rect 10400 33700 10404 33756
rect 10404 33700 10460 33756
rect 10460 33700 10464 33756
rect 10400 33696 10464 33700
rect 10480 33756 10544 33760
rect 10480 33700 10484 33756
rect 10484 33700 10540 33756
rect 10540 33700 10544 33756
rect 10480 33696 10544 33700
rect 10560 33756 10624 33760
rect 10560 33700 10564 33756
rect 10564 33700 10620 33756
rect 10620 33700 10624 33756
rect 10560 33696 10624 33700
rect 10640 33756 10704 33760
rect 10640 33700 10644 33756
rect 10644 33700 10700 33756
rect 10700 33700 10704 33756
rect 10640 33696 10704 33700
rect 19848 33756 19912 33760
rect 19848 33700 19852 33756
rect 19852 33700 19908 33756
rect 19908 33700 19912 33756
rect 19848 33696 19912 33700
rect 19928 33756 19992 33760
rect 19928 33700 19932 33756
rect 19932 33700 19988 33756
rect 19988 33700 19992 33756
rect 19928 33696 19992 33700
rect 20008 33756 20072 33760
rect 20008 33700 20012 33756
rect 20012 33700 20068 33756
rect 20068 33700 20072 33756
rect 20008 33696 20072 33700
rect 20088 33756 20152 33760
rect 20088 33700 20092 33756
rect 20092 33700 20148 33756
rect 20148 33700 20152 33756
rect 20088 33696 20152 33700
rect 29296 33756 29360 33760
rect 29296 33700 29300 33756
rect 29300 33700 29356 33756
rect 29356 33700 29360 33756
rect 29296 33696 29360 33700
rect 29376 33756 29440 33760
rect 29376 33700 29380 33756
rect 29380 33700 29436 33756
rect 29436 33700 29440 33756
rect 29376 33696 29440 33700
rect 29456 33756 29520 33760
rect 29456 33700 29460 33756
rect 29460 33700 29516 33756
rect 29516 33700 29520 33756
rect 29456 33696 29520 33700
rect 29536 33756 29600 33760
rect 29536 33700 29540 33756
rect 29540 33700 29596 33756
rect 29596 33700 29600 33756
rect 29536 33696 29600 33700
rect 5676 33212 5740 33216
rect 5676 33156 5680 33212
rect 5680 33156 5736 33212
rect 5736 33156 5740 33212
rect 5676 33152 5740 33156
rect 5756 33212 5820 33216
rect 5756 33156 5760 33212
rect 5760 33156 5816 33212
rect 5816 33156 5820 33212
rect 5756 33152 5820 33156
rect 5836 33212 5900 33216
rect 5836 33156 5840 33212
rect 5840 33156 5896 33212
rect 5896 33156 5900 33212
rect 5836 33152 5900 33156
rect 5916 33212 5980 33216
rect 5916 33156 5920 33212
rect 5920 33156 5976 33212
rect 5976 33156 5980 33212
rect 5916 33152 5980 33156
rect 15124 33212 15188 33216
rect 15124 33156 15128 33212
rect 15128 33156 15184 33212
rect 15184 33156 15188 33212
rect 15124 33152 15188 33156
rect 15204 33212 15268 33216
rect 15204 33156 15208 33212
rect 15208 33156 15264 33212
rect 15264 33156 15268 33212
rect 15204 33152 15268 33156
rect 15284 33212 15348 33216
rect 15284 33156 15288 33212
rect 15288 33156 15344 33212
rect 15344 33156 15348 33212
rect 15284 33152 15348 33156
rect 15364 33212 15428 33216
rect 15364 33156 15368 33212
rect 15368 33156 15424 33212
rect 15424 33156 15428 33212
rect 15364 33152 15428 33156
rect 24572 33212 24636 33216
rect 24572 33156 24576 33212
rect 24576 33156 24632 33212
rect 24632 33156 24636 33212
rect 24572 33152 24636 33156
rect 24652 33212 24716 33216
rect 24652 33156 24656 33212
rect 24656 33156 24712 33212
rect 24712 33156 24716 33212
rect 24652 33152 24716 33156
rect 24732 33212 24796 33216
rect 24732 33156 24736 33212
rect 24736 33156 24792 33212
rect 24792 33156 24796 33212
rect 24732 33152 24796 33156
rect 24812 33212 24876 33216
rect 24812 33156 24816 33212
rect 24816 33156 24872 33212
rect 24872 33156 24876 33212
rect 24812 33152 24876 33156
rect 34020 33212 34084 33216
rect 34020 33156 34024 33212
rect 34024 33156 34080 33212
rect 34080 33156 34084 33212
rect 34020 33152 34084 33156
rect 34100 33212 34164 33216
rect 34100 33156 34104 33212
rect 34104 33156 34160 33212
rect 34160 33156 34164 33212
rect 34100 33152 34164 33156
rect 34180 33212 34244 33216
rect 34180 33156 34184 33212
rect 34184 33156 34240 33212
rect 34240 33156 34244 33212
rect 34180 33152 34244 33156
rect 34260 33212 34324 33216
rect 34260 33156 34264 33212
rect 34264 33156 34320 33212
rect 34320 33156 34324 33212
rect 34260 33152 34324 33156
rect 10400 32668 10464 32672
rect 10400 32612 10404 32668
rect 10404 32612 10460 32668
rect 10460 32612 10464 32668
rect 10400 32608 10464 32612
rect 10480 32668 10544 32672
rect 10480 32612 10484 32668
rect 10484 32612 10540 32668
rect 10540 32612 10544 32668
rect 10480 32608 10544 32612
rect 10560 32668 10624 32672
rect 10560 32612 10564 32668
rect 10564 32612 10620 32668
rect 10620 32612 10624 32668
rect 10560 32608 10624 32612
rect 10640 32668 10704 32672
rect 10640 32612 10644 32668
rect 10644 32612 10700 32668
rect 10700 32612 10704 32668
rect 10640 32608 10704 32612
rect 19848 32668 19912 32672
rect 19848 32612 19852 32668
rect 19852 32612 19908 32668
rect 19908 32612 19912 32668
rect 19848 32608 19912 32612
rect 19928 32668 19992 32672
rect 19928 32612 19932 32668
rect 19932 32612 19988 32668
rect 19988 32612 19992 32668
rect 19928 32608 19992 32612
rect 20008 32668 20072 32672
rect 20008 32612 20012 32668
rect 20012 32612 20068 32668
rect 20068 32612 20072 32668
rect 20008 32608 20072 32612
rect 20088 32668 20152 32672
rect 20088 32612 20092 32668
rect 20092 32612 20148 32668
rect 20148 32612 20152 32668
rect 20088 32608 20152 32612
rect 29296 32668 29360 32672
rect 29296 32612 29300 32668
rect 29300 32612 29356 32668
rect 29356 32612 29360 32668
rect 29296 32608 29360 32612
rect 29376 32668 29440 32672
rect 29376 32612 29380 32668
rect 29380 32612 29436 32668
rect 29436 32612 29440 32668
rect 29376 32608 29440 32612
rect 29456 32668 29520 32672
rect 29456 32612 29460 32668
rect 29460 32612 29516 32668
rect 29516 32612 29520 32668
rect 29456 32608 29520 32612
rect 29536 32668 29600 32672
rect 29536 32612 29540 32668
rect 29540 32612 29596 32668
rect 29596 32612 29600 32668
rect 29536 32608 29600 32612
rect 5676 32124 5740 32128
rect 5676 32068 5680 32124
rect 5680 32068 5736 32124
rect 5736 32068 5740 32124
rect 5676 32064 5740 32068
rect 5756 32124 5820 32128
rect 5756 32068 5760 32124
rect 5760 32068 5816 32124
rect 5816 32068 5820 32124
rect 5756 32064 5820 32068
rect 5836 32124 5900 32128
rect 5836 32068 5840 32124
rect 5840 32068 5896 32124
rect 5896 32068 5900 32124
rect 5836 32064 5900 32068
rect 5916 32124 5980 32128
rect 5916 32068 5920 32124
rect 5920 32068 5976 32124
rect 5976 32068 5980 32124
rect 5916 32064 5980 32068
rect 15124 32124 15188 32128
rect 15124 32068 15128 32124
rect 15128 32068 15184 32124
rect 15184 32068 15188 32124
rect 15124 32064 15188 32068
rect 15204 32124 15268 32128
rect 15204 32068 15208 32124
rect 15208 32068 15264 32124
rect 15264 32068 15268 32124
rect 15204 32064 15268 32068
rect 15284 32124 15348 32128
rect 15284 32068 15288 32124
rect 15288 32068 15344 32124
rect 15344 32068 15348 32124
rect 15284 32064 15348 32068
rect 15364 32124 15428 32128
rect 15364 32068 15368 32124
rect 15368 32068 15424 32124
rect 15424 32068 15428 32124
rect 15364 32064 15428 32068
rect 24572 32124 24636 32128
rect 24572 32068 24576 32124
rect 24576 32068 24632 32124
rect 24632 32068 24636 32124
rect 24572 32064 24636 32068
rect 24652 32124 24716 32128
rect 24652 32068 24656 32124
rect 24656 32068 24712 32124
rect 24712 32068 24716 32124
rect 24652 32064 24716 32068
rect 24732 32124 24796 32128
rect 24732 32068 24736 32124
rect 24736 32068 24792 32124
rect 24792 32068 24796 32124
rect 24732 32064 24796 32068
rect 24812 32124 24876 32128
rect 24812 32068 24816 32124
rect 24816 32068 24872 32124
rect 24872 32068 24876 32124
rect 24812 32064 24876 32068
rect 34020 32124 34084 32128
rect 34020 32068 34024 32124
rect 34024 32068 34080 32124
rect 34080 32068 34084 32124
rect 34020 32064 34084 32068
rect 34100 32124 34164 32128
rect 34100 32068 34104 32124
rect 34104 32068 34160 32124
rect 34160 32068 34164 32124
rect 34100 32064 34164 32068
rect 34180 32124 34244 32128
rect 34180 32068 34184 32124
rect 34184 32068 34240 32124
rect 34240 32068 34244 32124
rect 34180 32064 34244 32068
rect 34260 32124 34324 32128
rect 34260 32068 34264 32124
rect 34264 32068 34320 32124
rect 34320 32068 34324 32124
rect 34260 32064 34324 32068
rect 10400 31580 10464 31584
rect 10400 31524 10404 31580
rect 10404 31524 10460 31580
rect 10460 31524 10464 31580
rect 10400 31520 10464 31524
rect 10480 31580 10544 31584
rect 10480 31524 10484 31580
rect 10484 31524 10540 31580
rect 10540 31524 10544 31580
rect 10480 31520 10544 31524
rect 10560 31580 10624 31584
rect 10560 31524 10564 31580
rect 10564 31524 10620 31580
rect 10620 31524 10624 31580
rect 10560 31520 10624 31524
rect 10640 31580 10704 31584
rect 10640 31524 10644 31580
rect 10644 31524 10700 31580
rect 10700 31524 10704 31580
rect 10640 31520 10704 31524
rect 19848 31580 19912 31584
rect 19848 31524 19852 31580
rect 19852 31524 19908 31580
rect 19908 31524 19912 31580
rect 19848 31520 19912 31524
rect 19928 31580 19992 31584
rect 19928 31524 19932 31580
rect 19932 31524 19988 31580
rect 19988 31524 19992 31580
rect 19928 31520 19992 31524
rect 20008 31580 20072 31584
rect 20008 31524 20012 31580
rect 20012 31524 20068 31580
rect 20068 31524 20072 31580
rect 20008 31520 20072 31524
rect 20088 31580 20152 31584
rect 20088 31524 20092 31580
rect 20092 31524 20148 31580
rect 20148 31524 20152 31580
rect 20088 31520 20152 31524
rect 29296 31580 29360 31584
rect 29296 31524 29300 31580
rect 29300 31524 29356 31580
rect 29356 31524 29360 31580
rect 29296 31520 29360 31524
rect 29376 31580 29440 31584
rect 29376 31524 29380 31580
rect 29380 31524 29436 31580
rect 29436 31524 29440 31580
rect 29376 31520 29440 31524
rect 29456 31580 29520 31584
rect 29456 31524 29460 31580
rect 29460 31524 29516 31580
rect 29516 31524 29520 31580
rect 29456 31520 29520 31524
rect 29536 31580 29600 31584
rect 29536 31524 29540 31580
rect 29540 31524 29596 31580
rect 29596 31524 29600 31580
rect 29536 31520 29600 31524
rect 5676 31036 5740 31040
rect 5676 30980 5680 31036
rect 5680 30980 5736 31036
rect 5736 30980 5740 31036
rect 5676 30976 5740 30980
rect 5756 31036 5820 31040
rect 5756 30980 5760 31036
rect 5760 30980 5816 31036
rect 5816 30980 5820 31036
rect 5756 30976 5820 30980
rect 5836 31036 5900 31040
rect 5836 30980 5840 31036
rect 5840 30980 5896 31036
rect 5896 30980 5900 31036
rect 5836 30976 5900 30980
rect 5916 31036 5980 31040
rect 5916 30980 5920 31036
rect 5920 30980 5976 31036
rect 5976 30980 5980 31036
rect 5916 30976 5980 30980
rect 15124 31036 15188 31040
rect 15124 30980 15128 31036
rect 15128 30980 15184 31036
rect 15184 30980 15188 31036
rect 15124 30976 15188 30980
rect 15204 31036 15268 31040
rect 15204 30980 15208 31036
rect 15208 30980 15264 31036
rect 15264 30980 15268 31036
rect 15204 30976 15268 30980
rect 15284 31036 15348 31040
rect 15284 30980 15288 31036
rect 15288 30980 15344 31036
rect 15344 30980 15348 31036
rect 15284 30976 15348 30980
rect 15364 31036 15428 31040
rect 15364 30980 15368 31036
rect 15368 30980 15424 31036
rect 15424 30980 15428 31036
rect 15364 30976 15428 30980
rect 24572 31036 24636 31040
rect 24572 30980 24576 31036
rect 24576 30980 24632 31036
rect 24632 30980 24636 31036
rect 24572 30976 24636 30980
rect 24652 31036 24716 31040
rect 24652 30980 24656 31036
rect 24656 30980 24712 31036
rect 24712 30980 24716 31036
rect 24652 30976 24716 30980
rect 24732 31036 24796 31040
rect 24732 30980 24736 31036
rect 24736 30980 24792 31036
rect 24792 30980 24796 31036
rect 24732 30976 24796 30980
rect 24812 31036 24876 31040
rect 24812 30980 24816 31036
rect 24816 30980 24872 31036
rect 24872 30980 24876 31036
rect 24812 30976 24876 30980
rect 34020 31036 34084 31040
rect 34020 30980 34024 31036
rect 34024 30980 34080 31036
rect 34080 30980 34084 31036
rect 34020 30976 34084 30980
rect 34100 31036 34164 31040
rect 34100 30980 34104 31036
rect 34104 30980 34160 31036
rect 34160 30980 34164 31036
rect 34100 30976 34164 30980
rect 34180 31036 34244 31040
rect 34180 30980 34184 31036
rect 34184 30980 34240 31036
rect 34240 30980 34244 31036
rect 34180 30976 34244 30980
rect 34260 31036 34324 31040
rect 34260 30980 34264 31036
rect 34264 30980 34320 31036
rect 34320 30980 34324 31036
rect 34260 30976 34324 30980
rect 10400 30492 10464 30496
rect 10400 30436 10404 30492
rect 10404 30436 10460 30492
rect 10460 30436 10464 30492
rect 10400 30432 10464 30436
rect 10480 30492 10544 30496
rect 10480 30436 10484 30492
rect 10484 30436 10540 30492
rect 10540 30436 10544 30492
rect 10480 30432 10544 30436
rect 10560 30492 10624 30496
rect 10560 30436 10564 30492
rect 10564 30436 10620 30492
rect 10620 30436 10624 30492
rect 10560 30432 10624 30436
rect 10640 30492 10704 30496
rect 10640 30436 10644 30492
rect 10644 30436 10700 30492
rect 10700 30436 10704 30492
rect 10640 30432 10704 30436
rect 19848 30492 19912 30496
rect 19848 30436 19852 30492
rect 19852 30436 19908 30492
rect 19908 30436 19912 30492
rect 19848 30432 19912 30436
rect 19928 30492 19992 30496
rect 19928 30436 19932 30492
rect 19932 30436 19988 30492
rect 19988 30436 19992 30492
rect 19928 30432 19992 30436
rect 20008 30492 20072 30496
rect 20008 30436 20012 30492
rect 20012 30436 20068 30492
rect 20068 30436 20072 30492
rect 20008 30432 20072 30436
rect 20088 30492 20152 30496
rect 20088 30436 20092 30492
rect 20092 30436 20148 30492
rect 20148 30436 20152 30492
rect 20088 30432 20152 30436
rect 29296 30492 29360 30496
rect 29296 30436 29300 30492
rect 29300 30436 29356 30492
rect 29356 30436 29360 30492
rect 29296 30432 29360 30436
rect 29376 30492 29440 30496
rect 29376 30436 29380 30492
rect 29380 30436 29436 30492
rect 29436 30436 29440 30492
rect 29376 30432 29440 30436
rect 29456 30492 29520 30496
rect 29456 30436 29460 30492
rect 29460 30436 29516 30492
rect 29516 30436 29520 30492
rect 29456 30432 29520 30436
rect 29536 30492 29600 30496
rect 29536 30436 29540 30492
rect 29540 30436 29596 30492
rect 29596 30436 29600 30492
rect 29536 30432 29600 30436
rect 5676 29948 5740 29952
rect 5676 29892 5680 29948
rect 5680 29892 5736 29948
rect 5736 29892 5740 29948
rect 5676 29888 5740 29892
rect 5756 29948 5820 29952
rect 5756 29892 5760 29948
rect 5760 29892 5816 29948
rect 5816 29892 5820 29948
rect 5756 29888 5820 29892
rect 5836 29948 5900 29952
rect 5836 29892 5840 29948
rect 5840 29892 5896 29948
rect 5896 29892 5900 29948
rect 5836 29888 5900 29892
rect 5916 29948 5980 29952
rect 5916 29892 5920 29948
rect 5920 29892 5976 29948
rect 5976 29892 5980 29948
rect 5916 29888 5980 29892
rect 15124 29948 15188 29952
rect 15124 29892 15128 29948
rect 15128 29892 15184 29948
rect 15184 29892 15188 29948
rect 15124 29888 15188 29892
rect 15204 29948 15268 29952
rect 15204 29892 15208 29948
rect 15208 29892 15264 29948
rect 15264 29892 15268 29948
rect 15204 29888 15268 29892
rect 15284 29948 15348 29952
rect 15284 29892 15288 29948
rect 15288 29892 15344 29948
rect 15344 29892 15348 29948
rect 15284 29888 15348 29892
rect 15364 29948 15428 29952
rect 15364 29892 15368 29948
rect 15368 29892 15424 29948
rect 15424 29892 15428 29948
rect 15364 29888 15428 29892
rect 24572 29948 24636 29952
rect 24572 29892 24576 29948
rect 24576 29892 24632 29948
rect 24632 29892 24636 29948
rect 24572 29888 24636 29892
rect 24652 29948 24716 29952
rect 24652 29892 24656 29948
rect 24656 29892 24712 29948
rect 24712 29892 24716 29948
rect 24652 29888 24716 29892
rect 24732 29948 24796 29952
rect 24732 29892 24736 29948
rect 24736 29892 24792 29948
rect 24792 29892 24796 29948
rect 24732 29888 24796 29892
rect 24812 29948 24876 29952
rect 24812 29892 24816 29948
rect 24816 29892 24872 29948
rect 24872 29892 24876 29948
rect 24812 29888 24876 29892
rect 34020 29948 34084 29952
rect 34020 29892 34024 29948
rect 34024 29892 34080 29948
rect 34080 29892 34084 29948
rect 34020 29888 34084 29892
rect 34100 29948 34164 29952
rect 34100 29892 34104 29948
rect 34104 29892 34160 29948
rect 34160 29892 34164 29948
rect 34100 29888 34164 29892
rect 34180 29948 34244 29952
rect 34180 29892 34184 29948
rect 34184 29892 34240 29948
rect 34240 29892 34244 29948
rect 34180 29888 34244 29892
rect 34260 29948 34324 29952
rect 34260 29892 34264 29948
rect 34264 29892 34320 29948
rect 34320 29892 34324 29948
rect 34260 29888 34324 29892
rect 10400 29404 10464 29408
rect 10400 29348 10404 29404
rect 10404 29348 10460 29404
rect 10460 29348 10464 29404
rect 10400 29344 10464 29348
rect 10480 29404 10544 29408
rect 10480 29348 10484 29404
rect 10484 29348 10540 29404
rect 10540 29348 10544 29404
rect 10480 29344 10544 29348
rect 10560 29404 10624 29408
rect 10560 29348 10564 29404
rect 10564 29348 10620 29404
rect 10620 29348 10624 29404
rect 10560 29344 10624 29348
rect 10640 29404 10704 29408
rect 10640 29348 10644 29404
rect 10644 29348 10700 29404
rect 10700 29348 10704 29404
rect 10640 29344 10704 29348
rect 19848 29404 19912 29408
rect 19848 29348 19852 29404
rect 19852 29348 19908 29404
rect 19908 29348 19912 29404
rect 19848 29344 19912 29348
rect 19928 29404 19992 29408
rect 19928 29348 19932 29404
rect 19932 29348 19988 29404
rect 19988 29348 19992 29404
rect 19928 29344 19992 29348
rect 20008 29404 20072 29408
rect 20008 29348 20012 29404
rect 20012 29348 20068 29404
rect 20068 29348 20072 29404
rect 20008 29344 20072 29348
rect 20088 29404 20152 29408
rect 20088 29348 20092 29404
rect 20092 29348 20148 29404
rect 20148 29348 20152 29404
rect 20088 29344 20152 29348
rect 29296 29404 29360 29408
rect 29296 29348 29300 29404
rect 29300 29348 29356 29404
rect 29356 29348 29360 29404
rect 29296 29344 29360 29348
rect 29376 29404 29440 29408
rect 29376 29348 29380 29404
rect 29380 29348 29436 29404
rect 29436 29348 29440 29404
rect 29376 29344 29440 29348
rect 29456 29404 29520 29408
rect 29456 29348 29460 29404
rect 29460 29348 29516 29404
rect 29516 29348 29520 29404
rect 29456 29344 29520 29348
rect 29536 29404 29600 29408
rect 29536 29348 29540 29404
rect 29540 29348 29596 29404
rect 29596 29348 29600 29404
rect 29536 29344 29600 29348
rect 5676 28860 5740 28864
rect 5676 28804 5680 28860
rect 5680 28804 5736 28860
rect 5736 28804 5740 28860
rect 5676 28800 5740 28804
rect 5756 28860 5820 28864
rect 5756 28804 5760 28860
rect 5760 28804 5816 28860
rect 5816 28804 5820 28860
rect 5756 28800 5820 28804
rect 5836 28860 5900 28864
rect 5836 28804 5840 28860
rect 5840 28804 5896 28860
rect 5896 28804 5900 28860
rect 5836 28800 5900 28804
rect 5916 28860 5980 28864
rect 5916 28804 5920 28860
rect 5920 28804 5976 28860
rect 5976 28804 5980 28860
rect 5916 28800 5980 28804
rect 15124 28860 15188 28864
rect 15124 28804 15128 28860
rect 15128 28804 15184 28860
rect 15184 28804 15188 28860
rect 15124 28800 15188 28804
rect 15204 28860 15268 28864
rect 15204 28804 15208 28860
rect 15208 28804 15264 28860
rect 15264 28804 15268 28860
rect 15204 28800 15268 28804
rect 15284 28860 15348 28864
rect 15284 28804 15288 28860
rect 15288 28804 15344 28860
rect 15344 28804 15348 28860
rect 15284 28800 15348 28804
rect 15364 28860 15428 28864
rect 15364 28804 15368 28860
rect 15368 28804 15424 28860
rect 15424 28804 15428 28860
rect 15364 28800 15428 28804
rect 24572 28860 24636 28864
rect 24572 28804 24576 28860
rect 24576 28804 24632 28860
rect 24632 28804 24636 28860
rect 24572 28800 24636 28804
rect 24652 28860 24716 28864
rect 24652 28804 24656 28860
rect 24656 28804 24712 28860
rect 24712 28804 24716 28860
rect 24652 28800 24716 28804
rect 24732 28860 24796 28864
rect 24732 28804 24736 28860
rect 24736 28804 24792 28860
rect 24792 28804 24796 28860
rect 24732 28800 24796 28804
rect 24812 28860 24876 28864
rect 24812 28804 24816 28860
rect 24816 28804 24872 28860
rect 24872 28804 24876 28860
rect 24812 28800 24876 28804
rect 34020 28860 34084 28864
rect 34020 28804 34024 28860
rect 34024 28804 34080 28860
rect 34080 28804 34084 28860
rect 34020 28800 34084 28804
rect 34100 28860 34164 28864
rect 34100 28804 34104 28860
rect 34104 28804 34160 28860
rect 34160 28804 34164 28860
rect 34100 28800 34164 28804
rect 34180 28860 34244 28864
rect 34180 28804 34184 28860
rect 34184 28804 34240 28860
rect 34240 28804 34244 28860
rect 34180 28800 34244 28804
rect 34260 28860 34324 28864
rect 34260 28804 34264 28860
rect 34264 28804 34320 28860
rect 34320 28804 34324 28860
rect 34260 28800 34324 28804
rect 10400 28316 10464 28320
rect 10400 28260 10404 28316
rect 10404 28260 10460 28316
rect 10460 28260 10464 28316
rect 10400 28256 10464 28260
rect 10480 28316 10544 28320
rect 10480 28260 10484 28316
rect 10484 28260 10540 28316
rect 10540 28260 10544 28316
rect 10480 28256 10544 28260
rect 10560 28316 10624 28320
rect 10560 28260 10564 28316
rect 10564 28260 10620 28316
rect 10620 28260 10624 28316
rect 10560 28256 10624 28260
rect 10640 28316 10704 28320
rect 10640 28260 10644 28316
rect 10644 28260 10700 28316
rect 10700 28260 10704 28316
rect 10640 28256 10704 28260
rect 19848 28316 19912 28320
rect 19848 28260 19852 28316
rect 19852 28260 19908 28316
rect 19908 28260 19912 28316
rect 19848 28256 19912 28260
rect 19928 28316 19992 28320
rect 19928 28260 19932 28316
rect 19932 28260 19988 28316
rect 19988 28260 19992 28316
rect 19928 28256 19992 28260
rect 20008 28316 20072 28320
rect 20008 28260 20012 28316
rect 20012 28260 20068 28316
rect 20068 28260 20072 28316
rect 20008 28256 20072 28260
rect 20088 28316 20152 28320
rect 20088 28260 20092 28316
rect 20092 28260 20148 28316
rect 20148 28260 20152 28316
rect 20088 28256 20152 28260
rect 29296 28316 29360 28320
rect 29296 28260 29300 28316
rect 29300 28260 29356 28316
rect 29356 28260 29360 28316
rect 29296 28256 29360 28260
rect 29376 28316 29440 28320
rect 29376 28260 29380 28316
rect 29380 28260 29436 28316
rect 29436 28260 29440 28316
rect 29376 28256 29440 28260
rect 29456 28316 29520 28320
rect 29456 28260 29460 28316
rect 29460 28260 29516 28316
rect 29516 28260 29520 28316
rect 29456 28256 29520 28260
rect 29536 28316 29600 28320
rect 29536 28260 29540 28316
rect 29540 28260 29596 28316
rect 29596 28260 29600 28316
rect 29536 28256 29600 28260
rect 5676 27772 5740 27776
rect 5676 27716 5680 27772
rect 5680 27716 5736 27772
rect 5736 27716 5740 27772
rect 5676 27712 5740 27716
rect 5756 27772 5820 27776
rect 5756 27716 5760 27772
rect 5760 27716 5816 27772
rect 5816 27716 5820 27772
rect 5756 27712 5820 27716
rect 5836 27772 5900 27776
rect 5836 27716 5840 27772
rect 5840 27716 5896 27772
rect 5896 27716 5900 27772
rect 5836 27712 5900 27716
rect 5916 27772 5980 27776
rect 5916 27716 5920 27772
rect 5920 27716 5976 27772
rect 5976 27716 5980 27772
rect 5916 27712 5980 27716
rect 15124 27772 15188 27776
rect 15124 27716 15128 27772
rect 15128 27716 15184 27772
rect 15184 27716 15188 27772
rect 15124 27712 15188 27716
rect 15204 27772 15268 27776
rect 15204 27716 15208 27772
rect 15208 27716 15264 27772
rect 15264 27716 15268 27772
rect 15204 27712 15268 27716
rect 15284 27772 15348 27776
rect 15284 27716 15288 27772
rect 15288 27716 15344 27772
rect 15344 27716 15348 27772
rect 15284 27712 15348 27716
rect 15364 27772 15428 27776
rect 15364 27716 15368 27772
rect 15368 27716 15424 27772
rect 15424 27716 15428 27772
rect 15364 27712 15428 27716
rect 24572 27772 24636 27776
rect 24572 27716 24576 27772
rect 24576 27716 24632 27772
rect 24632 27716 24636 27772
rect 24572 27712 24636 27716
rect 24652 27772 24716 27776
rect 24652 27716 24656 27772
rect 24656 27716 24712 27772
rect 24712 27716 24716 27772
rect 24652 27712 24716 27716
rect 24732 27772 24796 27776
rect 24732 27716 24736 27772
rect 24736 27716 24792 27772
rect 24792 27716 24796 27772
rect 24732 27712 24796 27716
rect 24812 27772 24876 27776
rect 24812 27716 24816 27772
rect 24816 27716 24872 27772
rect 24872 27716 24876 27772
rect 24812 27712 24876 27716
rect 34020 27772 34084 27776
rect 34020 27716 34024 27772
rect 34024 27716 34080 27772
rect 34080 27716 34084 27772
rect 34020 27712 34084 27716
rect 34100 27772 34164 27776
rect 34100 27716 34104 27772
rect 34104 27716 34160 27772
rect 34160 27716 34164 27772
rect 34100 27712 34164 27716
rect 34180 27772 34244 27776
rect 34180 27716 34184 27772
rect 34184 27716 34240 27772
rect 34240 27716 34244 27772
rect 34180 27712 34244 27716
rect 34260 27772 34324 27776
rect 34260 27716 34264 27772
rect 34264 27716 34320 27772
rect 34320 27716 34324 27772
rect 34260 27712 34324 27716
rect 10400 27228 10464 27232
rect 10400 27172 10404 27228
rect 10404 27172 10460 27228
rect 10460 27172 10464 27228
rect 10400 27168 10464 27172
rect 10480 27228 10544 27232
rect 10480 27172 10484 27228
rect 10484 27172 10540 27228
rect 10540 27172 10544 27228
rect 10480 27168 10544 27172
rect 10560 27228 10624 27232
rect 10560 27172 10564 27228
rect 10564 27172 10620 27228
rect 10620 27172 10624 27228
rect 10560 27168 10624 27172
rect 10640 27228 10704 27232
rect 10640 27172 10644 27228
rect 10644 27172 10700 27228
rect 10700 27172 10704 27228
rect 10640 27168 10704 27172
rect 19848 27228 19912 27232
rect 19848 27172 19852 27228
rect 19852 27172 19908 27228
rect 19908 27172 19912 27228
rect 19848 27168 19912 27172
rect 19928 27228 19992 27232
rect 19928 27172 19932 27228
rect 19932 27172 19988 27228
rect 19988 27172 19992 27228
rect 19928 27168 19992 27172
rect 20008 27228 20072 27232
rect 20008 27172 20012 27228
rect 20012 27172 20068 27228
rect 20068 27172 20072 27228
rect 20008 27168 20072 27172
rect 20088 27228 20152 27232
rect 20088 27172 20092 27228
rect 20092 27172 20148 27228
rect 20148 27172 20152 27228
rect 20088 27168 20152 27172
rect 29296 27228 29360 27232
rect 29296 27172 29300 27228
rect 29300 27172 29356 27228
rect 29356 27172 29360 27228
rect 29296 27168 29360 27172
rect 29376 27228 29440 27232
rect 29376 27172 29380 27228
rect 29380 27172 29436 27228
rect 29436 27172 29440 27228
rect 29376 27168 29440 27172
rect 29456 27228 29520 27232
rect 29456 27172 29460 27228
rect 29460 27172 29516 27228
rect 29516 27172 29520 27228
rect 29456 27168 29520 27172
rect 29536 27228 29600 27232
rect 29536 27172 29540 27228
rect 29540 27172 29596 27228
rect 29596 27172 29600 27228
rect 29536 27168 29600 27172
rect 5676 26684 5740 26688
rect 5676 26628 5680 26684
rect 5680 26628 5736 26684
rect 5736 26628 5740 26684
rect 5676 26624 5740 26628
rect 5756 26684 5820 26688
rect 5756 26628 5760 26684
rect 5760 26628 5816 26684
rect 5816 26628 5820 26684
rect 5756 26624 5820 26628
rect 5836 26684 5900 26688
rect 5836 26628 5840 26684
rect 5840 26628 5896 26684
rect 5896 26628 5900 26684
rect 5836 26624 5900 26628
rect 5916 26684 5980 26688
rect 5916 26628 5920 26684
rect 5920 26628 5976 26684
rect 5976 26628 5980 26684
rect 5916 26624 5980 26628
rect 15124 26684 15188 26688
rect 15124 26628 15128 26684
rect 15128 26628 15184 26684
rect 15184 26628 15188 26684
rect 15124 26624 15188 26628
rect 15204 26684 15268 26688
rect 15204 26628 15208 26684
rect 15208 26628 15264 26684
rect 15264 26628 15268 26684
rect 15204 26624 15268 26628
rect 15284 26684 15348 26688
rect 15284 26628 15288 26684
rect 15288 26628 15344 26684
rect 15344 26628 15348 26684
rect 15284 26624 15348 26628
rect 15364 26684 15428 26688
rect 15364 26628 15368 26684
rect 15368 26628 15424 26684
rect 15424 26628 15428 26684
rect 15364 26624 15428 26628
rect 24572 26684 24636 26688
rect 24572 26628 24576 26684
rect 24576 26628 24632 26684
rect 24632 26628 24636 26684
rect 24572 26624 24636 26628
rect 24652 26684 24716 26688
rect 24652 26628 24656 26684
rect 24656 26628 24712 26684
rect 24712 26628 24716 26684
rect 24652 26624 24716 26628
rect 24732 26684 24796 26688
rect 24732 26628 24736 26684
rect 24736 26628 24792 26684
rect 24792 26628 24796 26684
rect 24732 26624 24796 26628
rect 24812 26684 24876 26688
rect 24812 26628 24816 26684
rect 24816 26628 24872 26684
rect 24872 26628 24876 26684
rect 24812 26624 24876 26628
rect 34020 26684 34084 26688
rect 34020 26628 34024 26684
rect 34024 26628 34080 26684
rect 34080 26628 34084 26684
rect 34020 26624 34084 26628
rect 34100 26684 34164 26688
rect 34100 26628 34104 26684
rect 34104 26628 34160 26684
rect 34160 26628 34164 26684
rect 34100 26624 34164 26628
rect 34180 26684 34244 26688
rect 34180 26628 34184 26684
rect 34184 26628 34240 26684
rect 34240 26628 34244 26684
rect 34180 26624 34244 26628
rect 34260 26684 34324 26688
rect 34260 26628 34264 26684
rect 34264 26628 34320 26684
rect 34320 26628 34324 26684
rect 34260 26624 34324 26628
rect 10400 26140 10464 26144
rect 10400 26084 10404 26140
rect 10404 26084 10460 26140
rect 10460 26084 10464 26140
rect 10400 26080 10464 26084
rect 10480 26140 10544 26144
rect 10480 26084 10484 26140
rect 10484 26084 10540 26140
rect 10540 26084 10544 26140
rect 10480 26080 10544 26084
rect 10560 26140 10624 26144
rect 10560 26084 10564 26140
rect 10564 26084 10620 26140
rect 10620 26084 10624 26140
rect 10560 26080 10624 26084
rect 10640 26140 10704 26144
rect 10640 26084 10644 26140
rect 10644 26084 10700 26140
rect 10700 26084 10704 26140
rect 10640 26080 10704 26084
rect 19848 26140 19912 26144
rect 19848 26084 19852 26140
rect 19852 26084 19908 26140
rect 19908 26084 19912 26140
rect 19848 26080 19912 26084
rect 19928 26140 19992 26144
rect 19928 26084 19932 26140
rect 19932 26084 19988 26140
rect 19988 26084 19992 26140
rect 19928 26080 19992 26084
rect 20008 26140 20072 26144
rect 20008 26084 20012 26140
rect 20012 26084 20068 26140
rect 20068 26084 20072 26140
rect 20008 26080 20072 26084
rect 20088 26140 20152 26144
rect 20088 26084 20092 26140
rect 20092 26084 20148 26140
rect 20148 26084 20152 26140
rect 20088 26080 20152 26084
rect 29296 26140 29360 26144
rect 29296 26084 29300 26140
rect 29300 26084 29356 26140
rect 29356 26084 29360 26140
rect 29296 26080 29360 26084
rect 29376 26140 29440 26144
rect 29376 26084 29380 26140
rect 29380 26084 29436 26140
rect 29436 26084 29440 26140
rect 29376 26080 29440 26084
rect 29456 26140 29520 26144
rect 29456 26084 29460 26140
rect 29460 26084 29516 26140
rect 29516 26084 29520 26140
rect 29456 26080 29520 26084
rect 29536 26140 29600 26144
rect 29536 26084 29540 26140
rect 29540 26084 29596 26140
rect 29596 26084 29600 26140
rect 29536 26080 29600 26084
rect 5676 25596 5740 25600
rect 5676 25540 5680 25596
rect 5680 25540 5736 25596
rect 5736 25540 5740 25596
rect 5676 25536 5740 25540
rect 5756 25596 5820 25600
rect 5756 25540 5760 25596
rect 5760 25540 5816 25596
rect 5816 25540 5820 25596
rect 5756 25536 5820 25540
rect 5836 25596 5900 25600
rect 5836 25540 5840 25596
rect 5840 25540 5896 25596
rect 5896 25540 5900 25596
rect 5836 25536 5900 25540
rect 5916 25596 5980 25600
rect 5916 25540 5920 25596
rect 5920 25540 5976 25596
rect 5976 25540 5980 25596
rect 5916 25536 5980 25540
rect 15124 25596 15188 25600
rect 15124 25540 15128 25596
rect 15128 25540 15184 25596
rect 15184 25540 15188 25596
rect 15124 25536 15188 25540
rect 15204 25596 15268 25600
rect 15204 25540 15208 25596
rect 15208 25540 15264 25596
rect 15264 25540 15268 25596
rect 15204 25536 15268 25540
rect 15284 25596 15348 25600
rect 15284 25540 15288 25596
rect 15288 25540 15344 25596
rect 15344 25540 15348 25596
rect 15284 25536 15348 25540
rect 15364 25596 15428 25600
rect 15364 25540 15368 25596
rect 15368 25540 15424 25596
rect 15424 25540 15428 25596
rect 15364 25536 15428 25540
rect 24572 25596 24636 25600
rect 24572 25540 24576 25596
rect 24576 25540 24632 25596
rect 24632 25540 24636 25596
rect 24572 25536 24636 25540
rect 24652 25596 24716 25600
rect 24652 25540 24656 25596
rect 24656 25540 24712 25596
rect 24712 25540 24716 25596
rect 24652 25536 24716 25540
rect 24732 25596 24796 25600
rect 24732 25540 24736 25596
rect 24736 25540 24792 25596
rect 24792 25540 24796 25596
rect 24732 25536 24796 25540
rect 24812 25596 24876 25600
rect 24812 25540 24816 25596
rect 24816 25540 24872 25596
rect 24872 25540 24876 25596
rect 24812 25536 24876 25540
rect 34020 25596 34084 25600
rect 34020 25540 34024 25596
rect 34024 25540 34080 25596
rect 34080 25540 34084 25596
rect 34020 25536 34084 25540
rect 34100 25596 34164 25600
rect 34100 25540 34104 25596
rect 34104 25540 34160 25596
rect 34160 25540 34164 25596
rect 34100 25536 34164 25540
rect 34180 25596 34244 25600
rect 34180 25540 34184 25596
rect 34184 25540 34240 25596
rect 34240 25540 34244 25596
rect 34180 25536 34244 25540
rect 34260 25596 34324 25600
rect 34260 25540 34264 25596
rect 34264 25540 34320 25596
rect 34320 25540 34324 25596
rect 34260 25536 34324 25540
rect 10400 25052 10464 25056
rect 10400 24996 10404 25052
rect 10404 24996 10460 25052
rect 10460 24996 10464 25052
rect 10400 24992 10464 24996
rect 10480 25052 10544 25056
rect 10480 24996 10484 25052
rect 10484 24996 10540 25052
rect 10540 24996 10544 25052
rect 10480 24992 10544 24996
rect 10560 25052 10624 25056
rect 10560 24996 10564 25052
rect 10564 24996 10620 25052
rect 10620 24996 10624 25052
rect 10560 24992 10624 24996
rect 10640 25052 10704 25056
rect 10640 24996 10644 25052
rect 10644 24996 10700 25052
rect 10700 24996 10704 25052
rect 10640 24992 10704 24996
rect 19848 25052 19912 25056
rect 19848 24996 19852 25052
rect 19852 24996 19908 25052
rect 19908 24996 19912 25052
rect 19848 24992 19912 24996
rect 19928 25052 19992 25056
rect 19928 24996 19932 25052
rect 19932 24996 19988 25052
rect 19988 24996 19992 25052
rect 19928 24992 19992 24996
rect 20008 25052 20072 25056
rect 20008 24996 20012 25052
rect 20012 24996 20068 25052
rect 20068 24996 20072 25052
rect 20008 24992 20072 24996
rect 20088 25052 20152 25056
rect 20088 24996 20092 25052
rect 20092 24996 20148 25052
rect 20148 24996 20152 25052
rect 20088 24992 20152 24996
rect 29296 25052 29360 25056
rect 29296 24996 29300 25052
rect 29300 24996 29356 25052
rect 29356 24996 29360 25052
rect 29296 24992 29360 24996
rect 29376 25052 29440 25056
rect 29376 24996 29380 25052
rect 29380 24996 29436 25052
rect 29436 24996 29440 25052
rect 29376 24992 29440 24996
rect 29456 25052 29520 25056
rect 29456 24996 29460 25052
rect 29460 24996 29516 25052
rect 29516 24996 29520 25052
rect 29456 24992 29520 24996
rect 29536 25052 29600 25056
rect 29536 24996 29540 25052
rect 29540 24996 29596 25052
rect 29596 24996 29600 25052
rect 29536 24992 29600 24996
rect 5676 24508 5740 24512
rect 5676 24452 5680 24508
rect 5680 24452 5736 24508
rect 5736 24452 5740 24508
rect 5676 24448 5740 24452
rect 5756 24508 5820 24512
rect 5756 24452 5760 24508
rect 5760 24452 5816 24508
rect 5816 24452 5820 24508
rect 5756 24448 5820 24452
rect 5836 24508 5900 24512
rect 5836 24452 5840 24508
rect 5840 24452 5896 24508
rect 5896 24452 5900 24508
rect 5836 24448 5900 24452
rect 5916 24508 5980 24512
rect 5916 24452 5920 24508
rect 5920 24452 5976 24508
rect 5976 24452 5980 24508
rect 5916 24448 5980 24452
rect 15124 24508 15188 24512
rect 15124 24452 15128 24508
rect 15128 24452 15184 24508
rect 15184 24452 15188 24508
rect 15124 24448 15188 24452
rect 15204 24508 15268 24512
rect 15204 24452 15208 24508
rect 15208 24452 15264 24508
rect 15264 24452 15268 24508
rect 15204 24448 15268 24452
rect 15284 24508 15348 24512
rect 15284 24452 15288 24508
rect 15288 24452 15344 24508
rect 15344 24452 15348 24508
rect 15284 24448 15348 24452
rect 15364 24508 15428 24512
rect 15364 24452 15368 24508
rect 15368 24452 15424 24508
rect 15424 24452 15428 24508
rect 15364 24448 15428 24452
rect 24572 24508 24636 24512
rect 24572 24452 24576 24508
rect 24576 24452 24632 24508
rect 24632 24452 24636 24508
rect 24572 24448 24636 24452
rect 24652 24508 24716 24512
rect 24652 24452 24656 24508
rect 24656 24452 24712 24508
rect 24712 24452 24716 24508
rect 24652 24448 24716 24452
rect 24732 24508 24796 24512
rect 24732 24452 24736 24508
rect 24736 24452 24792 24508
rect 24792 24452 24796 24508
rect 24732 24448 24796 24452
rect 24812 24508 24876 24512
rect 24812 24452 24816 24508
rect 24816 24452 24872 24508
rect 24872 24452 24876 24508
rect 24812 24448 24876 24452
rect 34020 24508 34084 24512
rect 34020 24452 34024 24508
rect 34024 24452 34080 24508
rect 34080 24452 34084 24508
rect 34020 24448 34084 24452
rect 34100 24508 34164 24512
rect 34100 24452 34104 24508
rect 34104 24452 34160 24508
rect 34160 24452 34164 24508
rect 34100 24448 34164 24452
rect 34180 24508 34244 24512
rect 34180 24452 34184 24508
rect 34184 24452 34240 24508
rect 34240 24452 34244 24508
rect 34180 24448 34244 24452
rect 34260 24508 34324 24512
rect 34260 24452 34264 24508
rect 34264 24452 34320 24508
rect 34320 24452 34324 24508
rect 34260 24448 34324 24452
rect 10400 23964 10464 23968
rect 10400 23908 10404 23964
rect 10404 23908 10460 23964
rect 10460 23908 10464 23964
rect 10400 23904 10464 23908
rect 10480 23964 10544 23968
rect 10480 23908 10484 23964
rect 10484 23908 10540 23964
rect 10540 23908 10544 23964
rect 10480 23904 10544 23908
rect 10560 23964 10624 23968
rect 10560 23908 10564 23964
rect 10564 23908 10620 23964
rect 10620 23908 10624 23964
rect 10560 23904 10624 23908
rect 10640 23964 10704 23968
rect 10640 23908 10644 23964
rect 10644 23908 10700 23964
rect 10700 23908 10704 23964
rect 10640 23904 10704 23908
rect 19848 23964 19912 23968
rect 19848 23908 19852 23964
rect 19852 23908 19908 23964
rect 19908 23908 19912 23964
rect 19848 23904 19912 23908
rect 19928 23964 19992 23968
rect 19928 23908 19932 23964
rect 19932 23908 19988 23964
rect 19988 23908 19992 23964
rect 19928 23904 19992 23908
rect 20008 23964 20072 23968
rect 20008 23908 20012 23964
rect 20012 23908 20068 23964
rect 20068 23908 20072 23964
rect 20008 23904 20072 23908
rect 20088 23964 20152 23968
rect 20088 23908 20092 23964
rect 20092 23908 20148 23964
rect 20148 23908 20152 23964
rect 20088 23904 20152 23908
rect 29296 23964 29360 23968
rect 29296 23908 29300 23964
rect 29300 23908 29356 23964
rect 29356 23908 29360 23964
rect 29296 23904 29360 23908
rect 29376 23964 29440 23968
rect 29376 23908 29380 23964
rect 29380 23908 29436 23964
rect 29436 23908 29440 23964
rect 29376 23904 29440 23908
rect 29456 23964 29520 23968
rect 29456 23908 29460 23964
rect 29460 23908 29516 23964
rect 29516 23908 29520 23964
rect 29456 23904 29520 23908
rect 29536 23964 29600 23968
rect 29536 23908 29540 23964
rect 29540 23908 29596 23964
rect 29596 23908 29600 23964
rect 29536 23904 29600 23908
rect 5676 23420 5740 23424
rect 5676 23364 5680 23420
rect 5680 23364 5736 23420
rect 5736 23364 5740 23420
rect 5676 23360 5740 23364
rect 5756 23420 5820 23424
rect 5756 23364 5760 23420
rect 5760 23364 5816 23420
rect 5816 23364 5820 23420
rect 5756 23360 5820 23364
rect 5836 23420 5900 23424
rect 5836 23364 5840 23420
rect 5840 23364 5896 23420
rect 5896 23364 5900 23420
rect 5836 23360 5900 23364
rect 5916 23420 5980 23424
rect 5916 23364 5920 23420
rect 5920 23364 5976 23420
rect 5976 23364 5980 23420
rect 5916 23360 5980 23364
rect 15124 23420 15188 23424
rect 15124 23364 15128 23420
rect 15128 23364 15184 23420
rect 15184 23364 15188 23420
rect 15124 23360 15188 23364
rect 15204 23420 15268 23424
rect 15204 23364 15208 23420
rect 15208 23364 15264 23420
rect 15264 23364 15268 23420
rect 15204 23360 15268 23364
rect 15284 23420 15348 23424
rect 15284 23364 15288 23420
rect 15288 23364 15344 23420
rect 15344 23364 15348 23420
rect 15284 23360 15348 23364
rect 15364 23420 15428 23424
rect 15364 23364 15368 23420
rect 15368 23364 15424 23420
rect 15424 23364 15428 23420
rect 15364 23360 15428 23364
rect 24572 23420 24636 23424
rect 24572 23364 24576 23420
rect 24576 23364 24632 23420
rect 24632 23364 24636 23420
rect 24572 23360 24636 23364
rect 24652 23420 24716 23424
rect 24652 23364 24656 23420
rect 24656 23364 24712 23420
rect 24712 23364 24716 23420
rect 24652 23360 24716 23364
rect 24732 23420 24796 23424
rect 24732 23364 24736 23420
rect 24736 23364 24792 23420
rect 24792 23364 24796 23420
rect 24732 23360 24796 23364
rect 24812 23420 24876 23424
rect 24812 23364 24816 23420
rect 24816 23364 24872 23420
rect 24872 23364 24876 23420
rect 24812 23360 24876 23364
rect 34020 23420 34084 23424
rect 34020 23364 34024 23420
rect 34024 23364 34080 23420
rect 34080 23364 34084 23420
rect 34020 23360 34084 23364
rect 34100 23420 34164 23424
rect 34100 23364 34104 23420
rect 34104 23364 34160 23420
rect 34160 23364 34164 23420
rect 34100 23360 34164 23364
rect 34180 23420 34244 23424
rect 34180 23364 34184 23420
rect 34184 23364 34240 23420
rect 34240 23364 34244 23420
rect 34180 23360 34244 23364
rect 34260 23420 34324 23424
rect 34260 23364 34264 23420
rect 34264 23364 34320 23420
rect 34320 23364 34324 23420
rect 34260 23360 34324 23364
rect 10400 22876 10464 22880
rect 10400 22820 10404 22876
rect 10404 22820 10460 22876
rect 10460 22820 10464 22876
rect 10400 22816 10464 22820
rect 10480 22876 10544 22880
rect 10480 22820 10484 22876
rect 10484 22820 10540 22876
rect 10540 22820 10544 22876
rect 10480 22816 10544 22820
rect 10560 22876 10624 22880
rect 10560 22820 10564 22876
rect 10564 22820 10620 22876
rect 10620 22820 10624 22876
rect 10560 22816 10624 22820
rect 10640 22876 10704 22880
rect 10640 22820 10644 22876
rect 10644 22820 10700 22876
rect 10700 22820 10704 22876
rect 10640 22816 10704 22820
rect 19848 22876 19912 22880
rect 19848 22820 19852 22876
rect 19852 22820 19908 22876
rect 19908 22820 19912 22876
rect 19848 22816 19912 22820
rect 19928 22876 19992 22880
rect 19928 22820 19932 22876
rect 19932 22820 19988 22876
rect 19988 22820 19992 22876
rect 19928 22816 19992 22820
rect 20008 22876 20072 22880
rect 20008 22820 20012 22876
rect 20012 22820 20068 22876
rect 20068 22820 20072 22876
rect 20008 22816 20072 22820
rect 20088 22876 20152 22880
rect 20088 22820 20092 22876
rect 20092 22820 20148 22876
rect 20148 22820 20152 22876
rect 20088 22816 20152 22820
rect 29296 22876 29360 22880
rect 29296 22820 29300 22876
rect 29300 22820 29356 22876
rect 29356 22820 29360 22876
rect 29296 22816 29360 22820
rect 29376 22876 29440 22880
rect 29376 22820 29380 22876
rect 29380 22820 29436 22876
rect 29436 22820 29440 22876
rect 29376 22816 29440 22820
rect 29456 22876 29520 22880
rect 29456 22820 29460 22876
rect 29460 22820 29516 22876
rect 29516 22820 29520 22876
rect 29456 22816 29520 22820
rect 29536 22876 29600 22880
rect 29536 22820 29540 22876
rect 29540 22820 29596 22876
rect 29596 22820 29600 22876
rect 29536 22816 29600 22820
rect 5676 22332 5740 22336
rect 5676 22276 5680 22332
rect 5680 22276 5736 22332
rect 5736 22276 5740 22332
rect 5676 22272 5740 22276
rect 5756 22332 5820 22336
rect 5756 22276 5760 22332
rect 5760 22276 5816 22332
rect 5816 22276 5820 22332
rect 5756 22272 5820 22276
rect 5836 22332 5900 22336
rect 5836 22276 5840 22332
rect 5840 22276 5896 22332
rect 5896 22276 5900 22332
rect 5836 22272 5900 22276
rect 5916 22332 5980 22336
rect 5916 22276 5920 22332
rect 5920 22276 5976 22332
rect 5976 22276 5980 22332
rect 5916 22272 5980 22276
rect 15124 22332 15188 22336
rect 15124 22276 15128 22332
rect 15128 22276 15184 22332
rect 15184 22276 15188 22332
rect 15124 22272 15188 22276
rect 15204 22332 15268 22336
rect 15204 22276 15208 22332
rect 15208 22276 15264 22332
rect 15264 22276 15268 22332
rect 15204 22272 15268 22276
rect 15284 22332 15348 22336
rect 15284 22276 15288 22332
rect 15288 22276 15344 22332
rect 15344 22276 15348 22332
rect 15284 22272 15348 22276
rect 15364 22332 15428 22336
rect 15364 22276 15368 22332
rect 15368 22276 15424 22332
rect 15424 22276 15428 22332
rect 15364 22272 15428 22276
rect 24572 22332 24636 22336
rect 24572 22276 24576 22332
rect 24576 22276 24632 22332
rect 24632 22276 24636 22332
rect 24572 22272 24636 22276
rect 24652 22332 24716 22336
rect 24652 22276 24656 22332
rect 24656 22276 24712 22332
rect 24712 22276 24716 22332
rect 24652 22272 24716 22276
rect 24732 22332 24796 22336
rect 24732 22276 24736 22332
rect 24736 22276 24792 22332
rect 24792 22276 24796 22332
rect 24732 22272 24796 22276
rect 24812 22332 24876 22336
rect 24812 22276 24816 22332
rect 24816 22276 24872 22332
rect 24872 22276 24876 22332
rect 24812 22272 24876 22276
rect 34020 22332 34084 22336
rect 34020 22276 34024 22332
rect 34024 22276 34080 22332
rect 34080 22276 34084 22332
rect 34020 22272 34084 22276
rect 34100 22332 34164 22336
rect 34100 22276 34104 22332
rect 34104 22276 34160 22332
rect 34160 22276 34164 22332
rect 34100 22272 34164 22276
rect 34180 22332 34244 22336
rect 34180 22276 34184 22332
rect 34184 22276 34240 22332
rect 34240 22276 34244 22332
rect 34180 22272 34244 22276
rect 34260 22332 34324 22336
rect 34260 22276 34264 22332
rect 34264 22276 34320 22332
rect 34320 22276 34324 22332
rect 34260 22272 34324 22276
rect 10400 21788 10464 21792
rect 10400 21732 10404 21788
rect 10404 21732 10460 21788
rect 10460 21732 10464 21788
rect 10400 21728 10464 21732
rect 10480 21788 10544 21792
rect 10480 21732 10484 21788
rect 10484 21732 10540 21788
rect 10540 21732 10544 21788
rect 10480 21728 10544 21732
rect 10560 21788 10624 21792
rect 10560 21732 10564 21788
rect 10564 21732 10620 21788
rect 10620 21732 10624 21788
rect 10560 21728 10624 21732
rect 10640 21788 10704 21792
rect 10640 21732 10644 21788
rect 10644 21732 10700 21788
rect 10700 21732 10704 21788
rect 10640 21728 10704 21732
rect 19848 21788 19912 21792
rect 19848 21732 19852 21788
rect 19852 21732 19908 21788
rect 19908 21732 19912 21788
rect 19848 21728 19912 21732
rect 19928 21788 19992 21792
rect 19928 21732 19932 21788
rect 19932 21732 19988 21788
rect 19988 21732 19992 21788
rect 19928 21728 19992 21732
rect 20008 21788 20072 21792
rect 20008 21732 20012 21788
rect 20012 21732 20068 21788
rect 20068 21732 20072 21788
rect 20008 21728 20072 21732
rect 20088 21788 20152 21792
rect 20088 21732 20092 21788
rect 20092 21732 20148 21788
rect 20148 21732 20152 21788
rect 20088 21728 20152 21732
rect 29296 21788 29360 21792
rect 29296 21732 29300 21788
rect 29300 21732 29356 21788
rect 29356 21732 29360 21788
rect 29296 21728 29360 21732
rect 29376 21788 29440 21792
rect 29376 21732 29380 21788
rect 29380 21732 29436 21788
rect 29436 21732 29440 21788
rect 29376 21728 29440 21732
rect 29456 21788 29520 21792
rect 29456 21732 29460 21788
rect 29460 21732 29516 21788
rect 29516 21732 29520 21788
rect 29456 21728 29520 21732
rect 29536 21788 29600 21792
rect 29536 21732 29540 21788
rect 29540 21732 29596 21788
rect 29596 21732 29600 21788
rect 29536 21728 29600 21732
rect 5676 21244 5740 21248
rect 5676 21188 5680 21244
rect 5680 21188 5736 21244
rect 5736 21188 5740 21244
rect 5676 21184 5740 21188
rect 5756 21244 5820 21248
rect 5756 21188 5760 21244
rect 5760 21188 5816 21244
rect 5816 21188 5820 21244
rect 5756 21184 5820 21188
rect 5836 21244 5900 21248
rect 5836 21188 5840 21244
rect 5840 21188 5896 21244
rect 5896 21188 5900 21244
rect 5836 21184 5900 21188
rect 5916 21244 5980 21248
rect 5916 21188 5920 21244
rect 5920 21188 5976 21244
rect 5976 21188 5980 21244
rect 5916 21184 5980 21188
rect 15124 21244 15188 21248
rect 15124 21188 15128 21244
rect 15128 21188 15184 21244
rect 15184 21188 15188 21244
rect 15124 21184 15188 21188
rect 15204 21244 15268 21248
rect 15204 21188 15208 21244
rect 15208 21188 15264 21244
rect 15264 21188 15268 21244
rect 15204 21184 15268 21188
rect 15284 21244 15348 21248
rect 15284 21188 15288 21244
rect 15288 21188 15344 21244
rect 15344 21188 15348 21244
rect 15284 21184 15348 21188
rect 15364 21244 15428 21248
rect 15364 21188 15368 21244
rect 15368 21188 15424 21244
rect 15424 21188 15428 21244
rect 15364 21184 15428 21188
rect 24572 21244 24636 21248
rect 24572 21188 24576 21244
rect 24576 21188 24632 21244
rect 24632 21188 24636 21244
rect 24572 21184 24636 21188
rect 24652 21244 24716 21248
rect 24652 21188 24656 21244
rect 24656 21188 24712 21244
rect 24712 21188 24716 21244
rect 24652 21184 24716 21188
rect 24732 21244 24796 21248
rect 24732 21188 24736 21244
rect 24736 21188 24792 21244
rect 24792 21188 24796 21244
rect 24732 21184 24796 21188
rect 24812 21244 24876 21248
rect 24812 21188 24816 21244
rect 24816 21188 24872 21244
rect 24872 21188 24876 21244
rect 24812 21184 24876 21188
rect 34020 21244 34084 21248
rect 34020 21188 34024 21244
rect 34024 21188 34080 21244
rect 34080 21188 34084 21244
rect 34020 21184 34084 21188
rect 34100 21244 34164 21248
rect 34100 21188 34104 21244
rect 34104 21188 34160 21244
rect 34160 21188 34164 21244
rect 34100 21184 34164 21188
rect 34180 21244 34244 21248
rect 34180 21188 34184 21244
rect 34184 21188 34240 21244
rect 34240 21188 34244 21244
rect 34180 21184 34244 21188
rect 34260 21244 34324 21248
rect 34260 21188 34264 21244
rect 34264 21188 34320 21244
rect 34320 21188 34324 21244
rect 34260 21184 34324 21188
rect 10400 20700 10464 20704
rect 10400 20644 10404 20700
rect 10404 20644 10460 20700
rect 10460 20644 10464 20700
rect 10400 20640 10464 20644
rect 10480 20700 10544 20704
rect 10480 20644 10484 20700
rect 10484 20644 10540 20700
rect 10540 20644 10544 20700
rect 10480 20640 10544 20644
rect 10560 20700 10624 20704
rect 10560 20644 10564 20700
rect 10564 20644 10620 20700
rect 10620 20644 10624 20700
rect 10560 20640 10624 20644
rect 10640 20700 10704 20704
rect 10640 20644 10644 20700
rect 10644 20644 10700 20700
rect 10700 20644 10704 20700
rect 10640 20640 10704 20644
rect 19848 20700 19912 20704
rect 19848 20644 19852 20700
rect 19852 20644 19908 20700
rect 19908 20644 19912 20700
rect 19848 20640 19912 20644
rect 19928 20700 19992 20704
rect 19928 20644 19932 20700
rect 19932 20644 19988 20700
rect 19988 20644 19992 20700
rect 19928 20640 19992 20644
rect 20008 20700 20072 20704
rect 20008 20644 20012 20700
rect 20012 20644 20068 20700
rect 20068 20644 20072 20700
rect 20008 20640 20072 20644
rect 20088 20700 20152 20704
rect 20088 20644 20092 20700
rect 20092 20644 20148 20700
rect 20148 20644 20152 20700
rect 20088 20640 20152 20644
rect 29296 20700 29360 20704
rect 29296 20644 29300 20700
rect 29300 20644 29356 20700
rect 29356 20644 29360 20700
rect 29296 20640 29360 20644
rect 29376 20700 29440 20704
rect 29376 20644 29380 20700
rect 29380 20644 29436 20700
rect 29436 20644 29440 20700
rect 29376 20640 29440 20644
rect 29456 20700 29520 20704
rect 29456 20644 29460 20700
rect 29460 20644 29516 20700
rect 29516 20644 29520 20700
rect 29456 20640 29520 20644
rect 29536 20700 29600 20704
rect 29536 20644 29540 20700
rect 29540 20644 29596 20700
rect 29596 20644 29600 20700
rect 29536 20640 29600 20644
rect 5676 20156 5740 20160
rect 5676 20100 5680 20156
rect 5680 20100 5736 20156
rect 5736 20100 5740 20156
rect 5676 20096 5740 20100
rect 5756 20156 5820 20160
rect 5756 20100 5760 20156
rect 5760 20100 5816 20156
rect 5816 20100 5820 20156
rect 5756 20096 5820 20100
rect 5836 20156 5900 20160
rect 5836 20100 5840 20156
rect 5840 20100 5896 20156
rect 5896 20100 5900 20156
rect 5836 20096 5900 20100
rect 5916 20156 5980 20160
rect 5916 20100 5920 20156
rect 5920 20100 5976 20156
rect 5976 20100 5980 20156
rect 5916 20096 5980 20100
rect 15124 20156 15188 20160
rect 15124 20100 15128 20156
rect 15128 20100 15184 20156
rect 15184 20100 15188 20156
rect 15124 20096 15188 20100
rect 15204 20156 15268 20160
rect 15204 20100 15208 20156
rect 15208 20100 15264 20156
rect 15264 20100 15268 20156
rect 15204 20096 15268 20100
rect 15284 20156 15348 20160
rect 15284 20100 15288 20156
rect 15288 20100 15344 20156
rect 15344 20100 15348 20156
rect 15284 20096 15348 20100
rect 15364 20156 15428 20160
rect 15364 20100 15368 20156
rect 15368 20100 15424 20156
rect 15424 20100 15428 20156
rect 15364 20096 15428 20100
rect 24572 20156 24636 20160
rect 24572 20100 24576 20156
rect 24576 20100 24632 20156
rect 24632 20100 24636 20156
rect 24572 20096 24636 20100
rect 24652 20156 24716 20160
rect 24652 20100 24656 20156
rect 24656 20100 24712 20156
rect 24712 20100 24716 20156
rect 24652 20096 24716 20100
rect 24732 20156 24796 20160
rect 24732 20100 24736 20156
rect 24736 20100 24792 20156
rect 24792 20100 24796 20156
rect 24732 20096 24796 20100
rect 24812 20156 24876 20160
rect 24812 20100 24816 20156
rect 24816 20100 24872 20156
rect 24872 20100 24876 20156
rect 24812 20096 24876 20100
rect 34020 20156 34084 20160
rect 34020 20100 34024 20156
rect 34024 20100 34080 20156
rect 34080 20100 34084 20156
rect 34020 20096 34084 20100
rect 34100 20156 34164 20160
rect 34100 20100 34104 20156
rect 34104 20100 34160 20156
rect 34160 20100 34164 20156
rect 34100 20096 34164 20100
rect 34180 20156 34244 20160
rect 34180 20100 34184 20156
rect 34184 20100 34240 20156
rect 34240 20100 34244 20156
rect 34180 20096 34244 20100
rect 34260 20156 34324 20160
rect 34260 20100 34264 20156
rect 34264 20100 34320 20156
rect 34320 20100 34324 20156
rect 34260 20096 34324 20100
rect 10400 19612 10464 19616
rect 10400 19556 10404 19612
rect 10404 19556 10460 19612
rect 10460 19556 10464 19612
rect 10400 19552 10464 19556
rect 10480 19612 10544 19616
rect 10480 19556 10484 19612
rect 10484 19556 10540 19612
rect 10540 19556 10544 19612
rect 10480 19552 10544 19556
rect 10560 19612 10624 19616
rect 10560 19556 10564 19612
rect 10564 19556 10620 19612
rect 10620 19556 10624 19612
rect 10560 19552 10624 19556
rect 10640 19612 10704 19616
rect 10640 19556 10644 19612
rect 10644 19556 10700 19612
rect 10700 19556 10704 19612
rect 10640 19552 10704 19556
rect 19848 19612 19912 19616
rect 19848 19556 19852 19612
rect 19852 19556 19908 19612
rect 19908 19556 19912 19612
rect 19848 19552 19912 19556
rect 19928 19612 19992 19616
rect 19928 19556 19932 19612
rect 19932 19556 19988 19612
rect 19988 19556 19992 19612
rect 19928 19552 19992 19556
rect 20008 19612 20072 19616
rect 20008 19556 20012 19612
rect 20012 19556 20068 19612
rect 20068 19556 20072 19612
rect 20008 19552 20072 19556
rect 20088 19612 20152 19616
rect 20088 19556 20092 19612
rect 20092 19556 20148 19612
rect 20148 19556 20152 19612
rect 20088 19552 20152 19556
rect 29296 19612 29360 19616
rect 29296 19556 29300 19612
rect 29300 19556 29356 19612
rect 29356 19556 29360 19612
rect 29296 19552 29360 19556
rect 29376 19612 29440 19616
rect 29376 19556 29380 19612
rect 29380 19556 29436 19612
rect 29436 19556 29440 19612
rect 29376 19552 29440 19556
rect 29456 19612 29520 19616
rect 29456 19556 29460 19612
rect 29460 19556 29516 19612
rect 29516 19556 29520 19612
rect 29456 19552 29520 19556
rect 29536 19612 29600 19616
rect 29536 19556 29540 19612
rect 29540 19556 29596 19612
rect 29596 19556 29600 19612
rect 29536 19552 29600 19556
rect 5676 19068 5740 19072
rect 5676 19012 5680 19068
rect 5680 19012 5736 19068
rect 5736 19012 5740 19068
rect 5676 19008 5740 19012
rect 5756 19068 5820 19072
rect 5756 19012 5760 19068
rect 5760 19012 5816 19068
rect 5816 19012 5820 19068
rect 5756 19008 5820 19012
rect 5836 19068 5900 19072
rect 5836 19012 5840 19068
rect 5840 19012 5896 19068
rect 5896 19012 5900 19068
rect 5836 19008 5900 19012
rect 5916 19068 5980 19072
rect 5916 19012 5920 19068
rect 5920 19012 5976 19068
rect 5976 19012 5980 19068
rect 5916 19008 5980 19012
rect 15124 19068 15188 19072
rect 15124 19012 15128 19068
rect 15128 19012 15184 19068
rect 15184 19012 15188 19068
rect 15124 19008 15188 19012
rect 15204 19068 15268 19072
rect 15204 19012 15208 19068
rect 15208 19012 15264 19068
rect 15264 19012 15268 19068
rect 15204 19008 15268 19012
rect 15284 19068 15348 19072
rect 15284 19012 15288 19068
rect 15288 19012 15344 19068
rect 15344 19012 15348 19068
rect 15284 19008 15348 19012
rect 15364 19068 15428 19072
rect 15364 19012 15368 19068
rect 15368 19012 15424 19068
rect 15424 19012 15428 19068
rect 15364 19008 15428 19012
rect 24572 19068 24636 19072
rect 24572 19012 24576 19068
rect 24576 19012 24632 19068
rect 24632 19012 24636 19068
rect 24572 19008 24636 19012
rect 24652 19068 24716 19072
rect 24652 19012 24656 19068
rect 24656 19012 24712 19068
rect 24712 19012 24716 19068
rect 24652 19008 24716 19012
rect 24732 19068 24796 19072
rect 24732 19012 24736 19068
rect 24736 19012 24792 19068
rect 24792 19012 24796 19068
rect 24732 19008 24796 19012
rect 24812 19068 24876 19072
rect 24812 19012 24816 19068
rect 24816 19012 24872 19068
rect 24872 19012 24876 19068
rect 24812 19008 24876 19012
rect 34020 19068 34084 19072
rect 34020 19012 34024 19068
rect 34024 19012 34080 19068
rect 34080 19012 34084 19068
rect 34020 19008 34084 19012
rect 34100 19068 34164 19072
rect 34100 19012 34104 19068
rect 34104 19012 34160 19068
rect 34160 19012 34164 19068
rect 34100 19008 34164 19012
rect 34180 19068 34244 19072
rect 34180 19012 34184 19068
rect 34184 19012 34240 19068
rect 34240 19012 34244 19068
rect 34180 19008 34244 19012
rect 34260 19068 34324 19072
rect 34260 19012 34264 19068
rect 34264 19012 34320 19068
rect 34320 19012 34324 19068
rect 34260 19008 34324 19012
rect 10400 18524 10464 18528
rect 10400 18468 10404 18524
rect 10404 18468 10460 18524
rect 10460 18468 10464 18524
rect 10400 18464 10464 18468
rect 10480 18524 10544 18528
rect 10480 18468 10484 18524
rect 10484 18468 10540 18524
rect 10540 18468 10544 18524
rect 10480 18464 10544 18468
rect 10560 18524 10624 18528
rect 10560 18468 10564 18524
rect 10564 18468 10620 18524
rect 10620 18468 10624 18524
rect 10560 18464 10624 18468
rect 10640 18524 10704 18528
rect 10640 18468 10644 18524
rect 10644 18468 10700 18524
rect 10700 18468 10704 18524
rect 10640 18464 10704 18468
rect 19848 18524 19912 18528
rect 19848 18468 19852 18524
rect 19852 18468 19908 18524
rect 19908 18468 19912 18524
rect 19848 18464 19912 18468
rect 19928 18524 19992 18528
rect 19928 18468 19932 18524
rect 19932 18468 19988 18524
rect 19988 18468 19992 18524
rect 19928 18464 19992 18468
rect 20008 18524 20072 18528
rect 20008 18468 20012 18524
rect 20012 18468 20068 18524
rect 20068 18468 20072 18524
rect 20008 18464 20072 18468
rect 20088 18524 20152 18528
rect 20088 18468 20092 18524
rect 20092 18468 20148 18524
rect 20148 18468 20152 18524
rect 20088 18464 20152 18468
rect 29296 18524 29360 18528
rect 29296 18468 29300 18524
rect 29300 18468 29356 18524
rect 29356 18468 29360 18524
rect 29296 18464 29360 18468
rect 29376 18524 29440 18528
rect 29376 18468 29380 18524
rect 29380 18468 29436 18524
rect 29436 18468 29440 18524
rect 29376 18464 29440 18468
rect 29456 18524 29520 18528
rect 29456 18468 29460 18524
rect 29460 18468 29516 18524
rect 29516 18468 29520 18524
rect 29456 18464 29520 18468
rect 29536 18524 29600 18528
rect 29536 18468 29540 18524
rect 29540 18468 29596 18524
rect 29596 18468 29600 18524
rect 29536 18464 29600 18468
rect 5676 17980 5740 17984
rect 5676 17924 5680 17980
rect 5680 17924 5736 17980
rect 5736 17924 5740 17980
rect 5676 17920 5740 17924
rect 5756 17980 5820 17984
rect 5756 17924 5760 17980
rect 5760 17924 5816 17980
rect 5816 17924 5820 17980
rect 5756 17920 5820 17924
rect 5836 17980 5900 17984
rect 5836 17924 5840 17980
rect 5840 17924 5896 17980
rect 5896 17924 5900 17980
rect 5836 17920 5900 17924
rect 5916 17980 5980 17984
rect 5916 17924 5920 17980
rect 5920 17924 5976 17980
rect 5976 17924 5980 17980
rect 5916 17920 5980 17924
rect 15124 17980 15188 17984
rect 15124 17924 15128 17980
rect 15128 17924 15184 17980
rect 15184 17924 15188 17980
rect 15124 17920 15188 17924
rect 15204 17980 15268 17984
rect 15204 17924 15208 17980
rect 15208 17924 15264 17980
rect 15264 17924 15268 17980
rect 15204 17920 15268 17924
rect 15284 17980 15348 17984
rect 15284 17924 15288 17980
rect 15288 17924 15344 17980
rect 15344 17924 15348 17980
rect 15284 17920 15348 17924
rect 15364 17980 15428 17984
rect 15364 17924 15368 17980
rect 15368 17924 15424 17980
rect 15424 17924 15428 17980
rect 15364 17920 15428 17924
rect 24572 17980 24636 17984
rect 24572 17924 24576 17980
rect 24576 17924 24632 17980
rect 24632 17924 24636 17980
rect 24572 17920 24636 17924
rect 24652 17980 24716 17984
rect 24652 17924 24656 17980
rect 24656 17924 24712 17980
rect 24712 17924 24716 17980
rect 24652 17920 24716 17924
rect 24732 17980 24796 17984
rect 24732 17924 24736 17980
rect 24736 17924 24792 17980
rect 24792 17924 24796 17980
rect 24732 17920 24796 17924
rect 24812 17980 24876 17984
rect 24812 17924 24816 17980
rect 24816 17924 24872 17980
rect 24872 17924 24876 17980
rect 24812 17920 24876 17924
rect 34020 17980 34084 17984
rect 34020 17924 34024 17980
rect 34024 17924 34080 17980
rect 34080 17924 34084 17980
rect 34020 17920 34084 17924
rect 34100 17980 34164 17984
rect 34100 17924 34104 17980
rect 34104 17924 34160 17980
rect 34160 17924 34164 17980
rect 34100 17920 34164 17924
rect 34180 17980 34244 17984
rect 34180 17924 34184 17980
rect 34184 17924 34240 17980
rect 34240 17924 34244 17980
rect 34180 17920 34244 17924
rect 34260 17980 34324 17984
rect 34260 17924 34264 17980
rect 34264 17924 34320 17980
rect 34320 17924 34324 17980
rect 34260 17920 34324 17924
rect 10400 17436 10464 17440
rect 10400 17380 10404 17436
rect 10404 17380 10460 17436
rect 10460 17380 10464 17436
rect 10400 17376 10464 17380
rect 10480 17436 10544 17440
rect 10480 17380 10484 17436
rect 10484 17380 10540 17436
rect 10540 17380 10544 17436
rect 10480 17376 10544 17380
rect 10560 17436 10624 17440
rect 10560 17380 10564 17436
rect 10564 17380 10620 17436
rect 10620 17380 10624 17436
rect 10560 17376 10624 17380
rect 10640 17436 10704 17440
rect 10640 17380 10644 17436
rect 10644 17380 10700 17436
rect 10700 17380 10704 17436
rect 10640 17376 10704 17380
rect 19848 17436 19912 17440
rect 19848 17380 19852 17436
rect 19852 17380 19908 17436
rect 19908 17380 19912 17436
rect 19848 17376 19912 17380
rect 19928 17436 19992 17440
rect 19928 17380 19932 17436
rect 19932 17380 19988 17436
rect 19988 17380 19992 17436
rect 19928 17376 19992 17380
rect 20008 17436 20072 17440
rect 20008 17380 20012 17436
rect 20012 17380 20068 17436
rect 20068 17380 20072 17436
rect 20008 17376 20072 17380
rect 20088 17436 20152 17440
rect 20088 17380 20092 17436
rect 20092 17380 20148 17436
rect 20148 17380 20152 17436
rect 20088 17376 20152 17380
rect 29296 17436 29360 17440
rect 29296 17380 29300 17436
rect 29300 17380 29356 17436
rect 29356 17380 29360 17436
rect 29296 17376 29360 17380
rect 29376 17436 29440 17440
rect 29376 17380 29380 17436
rect 29380 17380 29436 17436
rect 29436 17380 29440 17436
rect 29376 17376 29440 17380
rect 29456 17436 29520 17440
rect 29456 17380 29460 17436
rect 29460 17380 29516 17436
rect 29516 17380 29520 17436
rect 29456 17376 29520 17380
rect 29536 17436 29600 17440
rect 29536 17380 29540 17436
rect 29540 17380 29596 17436
rect 29596 17380 29600 17436
rect 29536 17376 29600 17380
rect 5676 16892 5740 16896
rect 5676 16836 5680 16892
rect 5680 16836 5736 16892
rect 5736 16836 5740 16892
rect 5676 16832 5740 16836
rect 5756 16892 5820 16896
rect 5756 16836 5760 16892
rect 5760 16836 5816 16892
rect 5816 16836 5820 16892
rect 5756 16832 5820 16836
rect 5836 16892 5900 16896
rect 5836 16836 5840 16892
rect 5840 16836 5896 16892
rect 5896 16836 5900 16892
rect 5836 16832 5900 16836
rect 5916 16892 5980 16896
rect 5916 16836 5920 16892
rect 5920 16836 5976 16892
rect 5976 16836 5980 16892
rect 5916 16832 5980 16836
rect 15124 16892 15188 16896
rect 15124 16836 15128 16892
rect 15128 16836 15184 16892
rect 15184 16836 15188 16892
rect 15124 16832 15188 16836
rect 15204 16892 15268 16896
rect 15204 16836 15208 16892
rect 15208 16836 15264 16892
rect 15264 16836 15268 16892
rect 15204 16832 15268 16836
rect 15284 16892 15348 16896
rect 15284 16836 15288 16892
rect 15288 16836 15344 16892
rect 15344 16836 15348 16892
rect 15284 16832 15348 16836
rect 15364 16892 15428 16896
rect 15364 16836 15368 16892
rect 15368 16836 15424 16892
rect 15424 16836 15428 16892
rect 15364 16832 15428 16836
rect 24572 16892 24636 16896
rect 24572 16836 24576 16892
rect 24576 16836 24632 16892
rect 24632 16836 24636 16892
rect 24572 16832 24636 16836
rect 24652 16892 24716 16896
rect 24652 16836 24656 16892
rect 24656 16836 24712 16892
rect 24712 16836 24716 16892
rect 24652 16832 24716 16836
rect 24732 16892 24796 16896
rect 24732 16836 24736 16892
rect 24736 16836 24792 16892
rect 24792 16836 24796 16892
rect 24732 16832 24796 16836
rect 24812 16892 24876 16896
rect 24812 16836 24816 16892
rect 24816 16836 24872 16892
rect 24872 16836 24876 16892
rect 24812 16832 24876 16836
rect 34020 16892 34084 16896
rect 34020 16836 34024 16892
rect 34024 16836 34080 16892
rect 34080 16836 34084 16892
rect 34020 16832 34084 16836
rect 34100 16892 34164 16896
rect 34100 16836 34104 16892
rect 34104 16836 34160 16892
rect 34160 16836 34164 16892
rect 34100 16832 34164 16836
rect 34180 16892 34244 16896
rect 34180 16836 34184 16892
rect 34184 16836 34240 16892
rect 34240 16836 34244 16892
rect 34180 16832 34244 16836
rect 34260 16892 34324 16896
rect 34260 16836 34264 16892
rect 34264 16836 34320 16892
rect 34320 16836 34324 16892
rect 34260 16832 34324 16836
rect 10400 16348 10464 16352
rect 10400 16292 10404 16348
rect 10404 16292 10460 16348
rect 10460 16292 10464 16348
rect 10400 16288 10464 16292
rect 10480 16348 10544 16352
rect 10480 16292 10484 16348
rect 10484 16292 10540 16348
rect 10540 16292 10544 16348
rect 10480 16288 10544 16292
rect 10560 16348 10624 16352
rect 10560 16292 10564 16348
rect 10564 16292 10620 16348
rect 10620 16292 10624 16348
rect 10560 16288 10624 16292
rect 10640 16348 10704 16352
rect 10640 16292 10644 16348
rect 10644 16292 10700 16348
rect 10700 16292 10704 16348
rect 10640 16288 10704 16292
rect 19848 16348 19912 16352
rect 19848 16292 19852 16348
rect 19852 16292 19908 16348
rect 19908 16292 19912 16348
rect 19848 16288 19912 16292
rect 19928 16348 19992 16352
rect 19928 16292 19932 16348
rect 19932 16292 19988 16348
rect 19988 16292 19992 16348
rect 19928 16288 19992 16292
rect 20008 16348 20072 16352
rect 20008 16292 20012 16348
rect 20012 16292 20068 16348
rect 20068 16292 20072 16348
rect 20008 16288 20072 16292
rect 20088 16348 20152 16352
rect 20088 16292 20092 16348
rect 20092 16292 20148 16348
rect 20148 16292 20152 16348
rect 20088 16288 20152 16292
rect 29296 16348 29360 16352
rect 29296 16292 29300 16348
rect 29300 16292 29356 16348
rect 29356 16292 29360 16348
rect 29296 16288 29360 16292
rect 29376 16348 29440 16352
rect 29376 16292 29380 16348
rect 29380 16292 29436 16348
rect 29436 16292 29440 16348
rect 29376 16288 29440 16292
rect 29456 16348 29520 16352
rect 29456 16292 29460 16348
rect 29460 16292 29516 16348
rect 29516 16292 29520 16348
rect 29456 16288 29520 16292
rect 29536 16348 29600 16352
rect 29536 16292 29540 16348
rect 29540 16292 29596 16348
rect 29596 16292 29600 16348
rect 29536 16288 29600 16292
rect 5676 15804 5740 15808
rect 5676 15748 5680 15804
rect 5680 15748 5736 15804
rect 5736 15748 5740 15804
rect 5676 15744 5740 15748
rect 5756 15804 5820 15808
rect 5756 15748 5760 15804
rect 5760 15748 5816 15804
rect 5816 15748 5820 15804
rect 5756 15744 5820 15748
rect 5836 15804 5900 15808
rect 5836 15748 5840 15804
rect 5840 15748 5896 15804
rect 5896 15748 5900 15804
rect 5836 15744 5900 15748
rect 5916 15804 5980 15808
rect 5916 15748 5920 15804
rect 5920 15748 5976 15804
rect 5976 15748 5980 15804
rect 5916 15744 5980 15748
rect 15124 15804 15188 15808
rect 15124 15748 15128 15804
rect 15128 15748 15184 15804
rect 15184 15748 15188 15804
rect 15124 15744 15188 15748
rect 15204 15804 15268 15808
rect 15204 15748 15208 15804
rect 15208 15748 15264 15804
rect 15264 15748 15268 15804
rect 15204 15744 15268 15748
rect 15284 15804 15348 15808
rect 15284 15748 15288 15804
rect 15288 15748 15344 15804
rect 15344 15748 15348 15804
rect 15284 15744 15348 15748
rect 15364 15804 15428 15808
rect 15364 15748 15368 15804
rect 15368 15748 15424 15804
rect 15424 15748 15428 15804
rect 15364 15744 15428 15748
rect 24572 15804 24636 15808
rect 24572 15748 24576 15804
rect 24576 15748 24632 15804
rect 24632 15748 24636 15804
rect 24572 15744 24636 15748
rect 24652 15804 24716 15808
rect 24652 15748 24656 15804
rect 24656 15748 24712 15804
rect 24712 15748 24716 15804
rect 24652 15744 24716 15748
rect 24732 15804 24796 15808
rect 24732 15748 24736 15804
rect 24736 15748 24792 15804
rect 24792 15748 24796 15804
rect 24732 15744 24796 15748
rect 24812 15804 24876 15808
rect 24812 15748 24816 15804
rect 24816 15748 24872 15804
rect 24872 15748 24876 15804
rect 24812 15744 24876 15748
rect 34020 15804 34084 15808
rect 34020 15748 34024 15804
rect 34024 15748 34080 15804
rect 34080 15748 34084 15804
rect 34020 15744 34084 15748
rect 34100 15804 34164 15808
rect 34100 15748 34104 15804
rect 34104 15748 34160 15804
rect 34160 15748 34164 15804
rect 34100 15744 34164 15748
rect 34180 15804 34244 15808
rect 34180 15748 34184 15804
rect 34184 15748 34240 15804
rect 34240 15748 34244 15804
rect 34180 15744 34244 15748
rect 34260 15804 34324 15808
rect 34260 15748 34264 15804
rect 34264 15748 34320 15804
rect 34320 15748 34324 15804
rect 34260 15744 34324 15748
rect 10400 15260 10464 15264
rect 10400 15204 10404 15260
rect 10404 15204 10460 15260
rect 10460 15204 10464 15260
rect 10400 15200 10464 15204
rect 10480 15260 10544 15264
rect 10480 15204 10484 15260
rect 10484 15204 10540 15260
rect 10540 15204 10544 15260
rect 10480 15200 10544 15204
rect 10560 15260 10624 15264
rect 10560 15204 10564 15260
rect 10564 15204 10620 15260
rect 10620 15204 10624 15260
rect 10560 15200 10624 15204
rect 10640 15260 10704 15264
rect 10640 15204 10644 15260
rect 10644 15204 10700 15260
rect 10700 15204 10704 15260
rect 10640 15200 10704 15204
rect 19848 15260 19912 15264
rect 19848 15204 19852 15260
rect 19852 15204 19908 15260
rect 19908 15204 19912 15260
rect 19848 15200 19912 15204
rect 19928 15260 19992 15264
rect 19928 15204 19932 15260
rect 19932 15204 19988 15260
rect 19988 15204 19992 15260
rect 19928 15200 19992 15204
rect 20008 15260 20072 15264
rect 20008 15204 20012 15260
rect 20012 15204 20068 15260
rect 20068 15204 20072 15260
rect 20008 15200 20072 15204
rect 20088 15260 20152 15264
rect 20088 15204 20092 15260
rect 20092 15204 20148 15260
rect 20148 15204 20152 15260
rect 20088 15200 20152 15204
rect 29296 15260 29360 15264
rect 29296 15204 29300 15260
rect 29300 15204 29356 15260
rect 29356 15204 29360 15260
rect 29296 15200 29360 15204
rect 29376 15260 29440 15264
rect 29376 15204 29380 15260
rect 29380 15204 29436 15260
rect 29436 15204 29440 15260
rect 29376 15200 29440 15204
rect 29456 15260 29520 15264
rect 29456 15204 29460 15260
rect 29460 15204 29516 15260
rect 29516 15204 29520 15260
rect 29456 15200 29520 15204
rect 29536 15260 29600 15264
rect 29536 15204 29540 15260
rect 29540 15204 29596 15260
rect 29596 15204 29600 15260
rect 29536 15200 29600 15204
rect 5676 14716 5740 14720
rect 5676 14660 5680 14716
rect 5680 14660 5736 14716
rect 5736 14660 5740 14716
rect 5676 14656 5740 14660
rect 5756 14716 5820 14720
rect 5756 14660 5760 14716
rect 5760 14660 5816 14716
rect 5816 14660 5820 14716
rect 5756 14656 5820 14660
rect 5836 14716 5900 14720
rect 5836 14660 5840 14716
rect 5840 14660 5896 14716
rect 5896 14660 5900 14716
rect 5836 14656 5900 14660
rect 5916 14716 5980 14720
rect 5916 14660 5920 14716
rect 5920 14660 5976 14716
rect 5976 14660 5980 14716
rect 5916 14656 5980 14660
rect 15124 14716 15188 14720
rect 15124 14660 15128 14716
rect 15128 14660 15184 14716
rect 15184 14660 15188 14716
rect 15124 14656 15188 14660
rect 15204 14716 15268 14720
rect 15204 14660 15208 14716
rect 15208 14660 15264 14716
rect 15264 14660 15268 14716
rect 15204 14656 15268 14660
rect 15284 14716 15348 14720
rect 15284 14660 15288 14716
rect 15288 14660 15344 14716
rect 15344 14660 15348 14716
rect 15284 14656 15348 14660
rect 15364 14716 15428 14720
rect 15364 14660 15368 14716
rect 15368 14660 15424 14716
rect 15424 14660 15428 14716
rect 15364 14656 15428 14660
rect 24572 14716 24636 14720
rect 24572 14660 24576 14716
rect 24576 14660 24632 14716
rect 24632 14660 24636 14716
rect 24572 14656 24636 14660
rect 24652 14716 24716 14720
rect 24652 14660 24656 14716
rect 24656 14660 24712 14716
rect 24712 14660 24716 14716
rect 24652 14656 24716 14660
rect 24732 14716 24796 14720
rect 24732 14660 24736 14716
rect 24736 14660 24792 14716
rect 24792 14660 24796 14716
rect 24732 14656 24796 14660
rect 24812 14716 24876 14720
rect 24812 14660 24816 14716
rect 24816 14660 24872 14716
rect 24872 14660 24876 14716
rect 24812 14656 24876 14660
rect 34020 14716 34084 14720
rect 34020 14660 34024 14716
rect 34024 14660 34080 14716
rect 34080 14660 34084 14716
rect 34020 14656 34084 14660
rect 34100 14716 34164 14720
rect 34100 14660 34104 14716
rect 34104 14660 34160 14716
rect 34160 14660 34164 14716
rect 34100 14656 34164 14660
rect 34180 14716 34244 14720
rect 34180 14660 34184 14716
rect 34184 14660 34240 14716
rect 34240 14660 34244 14716
rect 34180 14656 34244 14660
rect 34260 14716 34324 14720
rect 34260 14660 34264 14716
rect 34264 14660 34320 14716
rect 34320 14660 34324 14716
rect 34260 14656 34324 14660
rect 10400 14172 10464 14176
rect 10400 14116 10404 14172
rect 10404 14116 10460 14172
rect 10460 14116 10464 14172
rect 10400 14112 10464 14116
rect 10480 14172 10544 14176
rect 10480 14116 10484 14172
rect 10484 14116 10540 14172
rect 10540 14116 10544 14172
rect 10480 14112 10544 14116
rect 10560 14172 10624 14176
rect 10560 14116 10564 14172
rect 10564 14116 10620 14172
rect 10620 14116 10624 14172
rect 10560 14112 10624 14116
rect 10640 14172 10704 14176
rect 10640 14116 10644 14172
rect 10644 14116 10700 14172
rect 10700 14116 10704 14172
rect 10640 14112 10704 14116
rect 19848 14172 19912 14176
rect 19848 14116 19852 14172
rect 19852 14116 19908 14172
rect 19908 14116 19912 14172
rect 19848 14112 19912 14116
rect 19928 14172 19992 14176
rect 19928 14116 19932 14172
rect 19932 14116 19988 14172
rect 19988 14116 19992 14172
rect 19928 14112 19992 14116
rect 20008 14172 20072 14176
rect 20008 14116 20012 14172
rect 20012 14116 20068 14172
rect 20068 14116 20072 14172
rect 20008 14112 20072 14116
rect 20088 14172 20152 14176
rect 20088 14116 20092 14172
rect 20092 14116 20148 14172
rect 20148 14116 20152 14172
rect 20088 14112 20152 14116
rect 29296 14172 29360 14176
rect 29296 14116 29300 14172
rect 29300 14116 29356 14172
rect 29356 14116 29360 14172
rect 29296 14112 29360 14116
rect 29376 14172 29440 14176
rect 29376 14116 29380 14172
rect 29380 14116 29436 14172
rect 29436 14116 29440 14172
rect 29376 14112 29440 14116
rect 29456 14172 29520 14176
rect 29456 14116 29460 14172
rect 29460 14116 29516 14172
rect 29516 14116 29520 14172
rect 29456 14112 29520 14116
rect 29536 14172 29600 14176
rect 29536 14116 29540 14172
rect 29540 14116 29596 14172
rect 29596 14116 29600 14172
rect 29536 14112 29600 14116
rect 5676 13628 5740 13632
rect 5676 13572 5680 13628
rect 5680 13572 5736 13628
rect 5736 13572 5740 13628
rect 5676 13568 5740 13572
rect 5756 13628 5820 13632
rect 5756 13572 5760 13628
rect 5760 13572 5816 13628
rect 5816 13572 5820 13628
rect 5756 13568 5820 13572
rect 5836 13628 5900 13632
rect 5836 13572 5840 13628
rect 5840 13572 5896 13628
rect 5896 13572 5900 13628
rect 5836 13568 5900 13572
rect 5916 13628 5980 13632
rect 5916 13572 5920 13628
rect 5920 13572 5976 13628
rect 5976 13572 5980 13628
rect 5916 13568 5980 13572
rect 15124 13628 15188 13632
rect 15124 13572 15128 13628
rect 15128 13572 15184 13628
rect 15184 13572 15188 13628
rect 15124 13568 15188 13572
rect 15204 13628 15268 13632
rect 15204 13572 15208 13628
rect 15208 13572 15264 13628
rect 15264 13572 15268 13628
rect 15204 13568 15268 13572
rect 15284 13628 15348 13632
rect 15284 13572 15288 13628
rect 15288 13572 15344 13628
rect 15344 13572 15348 13628
rect 15284 13568 15348 13572
rect 15364 13628 15428 13632
rect 15364 13572 15368 13628
rect 15368 13572 15424 13628
rect 15424 13572 15428 13628
rect 15364 13568 15428 13572
rect 24572 13628 24636 13632
rect 24572 13572 24576 13628
rect 24576 13572 24632 13628
rect 24632 13572 24636 13628
rect 24572 13568 24636 13572
rect 24652 13628 24716 13632
rect 24652 13572 24656 13628
rect 24656 13572 24712 13628
rect 24712 13572 24716 13628
rect 24652 13568 24716 13572
rect 24732 13628 24796 13632
rect 24732 13572 24736 13628
rect 24736 13572 24792 13628
rect 24792 13572 24796 13628
rect 24732 13568 24796 13572
rect 24812 13628 24876 13632
rect 24812 13572 24816 13628
rect 24816 13572 24872 13628
rect 24872 13572 24876 13628
rect 24812 13568 24876 13572
rect 34020 13628 34084 13632
rect 34020 13572 34024 13628
rect 34024 13572 34080 13628
rect 34080 13572 34084 13628
rect 34020 13568 34084 13572
rect 34100 13628 34164 13632
rect 34100 13572 34104 13628
rect 34104 13572 34160 13628
rect 34160 13572 34164 13628
rect 34100 13568 34164 13572
rect 34180 13628 34244 13632
rect 34180 13572 34184 13628
rect 34184 13572 34240 13628
rect 34240 13572 34244 13628
rect 34180 13568 34244 13572
rect 34260 13628 34324 13632
rect 34260 13572 34264 13628
rect 34264 13572 34320 13628
rect 34320 13572 34324 13628
rect 34260 13568 34324 13572
rect 10400 13084 10464 13088
rect 10400 13028 10404 13084
rect 10404 13028 10460 13084
rect 10460 13028 10464 13084
rect 10400 13024 10464 13028
rect 10480 13084 10544 13088
rect 10480 13028 10484 13084
rect 10484 13028 10540 13084
rect 10540 13028 10544 13084
rect 10480 13024 10544 13028
rect 10560 13084 10624 13088
rect 10560 13028 10564 13084
rect 10564 13028 10620 13084
rect 10620 13028 10624 13084
rect 10560 13024 10624 13028
rect 10640 13084 10704 13088
rect 10640 13028 10644 13084
rect 10644 13028 10700 13084
rect 10700 13028 10704 13084
rect 10640 13024 10704 13028
rect 19848 13084 19912 13088
rect 19848 13028 19852 13084
rect 19852 13028 19908 13084
rect 19908 13028 19912 13084
rect 19848 13024 19912 13028
rect 19928 13084 19992 13088
rect 19928 13028 19932 13084
rect 19932 13028 19988 13084
rect 19988 13028 19992 13084
rect 19928 13024 19992 13028
rect 20008 13084 20072 13088
rect 20008 13028 20012 13084
rect 20012 13028 20068 13084
rect 20068 13028 20072 13084
rect 20008 13024 20072 13028
rect 20088 13084 20152 13088
rect 20088 13028 20092 13084
rect 20092 13028 20148 13084
rect 20148 13028 20152 13084
rect 20088 13024 20152 13028
rect 29296 13084 29360 13088
rect 29296 13028 29300 13084
rect 29300 13028 29356 13084
rect 29356 13028 29360 13084
rect 29296 13024 29360 13028
rect 29376 13084 29440 13088
rect 29376 13028 29380 13084
rect 29380 13028 29436 13084
rect 29436 13028 29440 13084
rect 29376 13024 29440 13028
rect 29456 13084 29520 13088
rect 29456 13028 29460 13084
rect 29460 13028 29516 13084
rect 29516 13028 29520 13084
rect 29456 13024 29520 13028
rect 29536 13084 29600 13088
rect 29536 13028 29540 13084
rect 29540 13028 29596 13084
rect 29596 13028 29600 13084
rect 29536 13024 29600 13028
rect 5676 12540 5740 12544
rect 5676 12484 5680 12540
rect 5680 12484 5736 12540
rect 5736 12484 5740 12540
rect 5676 12480 5740 12484
rect 5756 12540 5820 12544
rect 5756 12484 5760 12540
rect 5760 12484 5816 12540
rect 5816 12484 5820 12540
rect 5756 12480 5820 12484
rect 5836 12540 5900 12544
rect 5836 12484 5840 12540
rect 5840 12484 5896 12540
rect 5896 12484 5900 12540
rect 5836 12480 5900 12484
rect 5916 12540 5980 12544
rect 5916 12484 5920 12540
rect 5920 12484 5976 12540
rect 5976 12484 5980 12540
rect 5916 12480 5980 12484
rect 15124 12540 15188 12544
rect 15124 12484 15128 12540
rect 15128 12484 15184 12540
rect 15184 12484 15188 12540
rect 15124 12480 15188 12484
rect 15204 12540 15268 12544
rect 15204 12484 15208 12540
rect 15208 12484 15264 12540
rect 15264 12484 15268 12540
rect 15204 12480 15268 12484
rect 15284 12540 15348 12544
rect 15284 12484 15288 12540
rect 15288 12484 15344 12540
rect 15344 12484 15348 12540
rect 15284 12480 15348 12484
rect 15364 12540 15428 12544
rect 15364 12484 15368 12540
rect 15368 12484 15424 12540
rect 15424 12484 15428 12540
rect 15364 12480 15428 12484
rect 24572 12540 24636 12544
rect 24572 12484 24576 12540
rect 24576 12484 24632 12540
rect 24632 12484 24636 12540
rect 24572 12480 24636 12484
rect 24652 12540 24716 12544
rect 24652 12484 24656 12540
rect 24656 12484 24712 12540
rect 24712 12484 24716 12540
rect 24652 12480 24716 12484
rect 24732 12540 24796 12544
rect 24732 12484 24736 12540
rect 24736 12484 24792 12540
rect 24792 12484 24796 12540
rect 24732 12480 24796 12484
rect 24812 12540 24876 12544
rect 24812 12484 24816 12540
rect 24816 12484 24872 12540
rect 24872 12484 24876 12540
rect 24812 12480 24876 12484
rect 34020 12540 34084 12544
rect 34020 12484 34024 12540
rect 34024 12484 34080 12540
rect 34080 12484 34084 12540
rect 34020 12480 34084 12484
rect 34100 12540 34164 12544
rect 34100 12484 34104 12540
rect 34104 12484 34160 12540
rect 34160 12484 34164 12540
rect 34100 12480 34164 12484
rect 34180 12540 34244 12544
rect 34180 12484 34184 12540
rect 34184 12484 34240 12540
rect 34240 12484 34244 12540
rect 34180 12480 34244 12484
rect 34260 12540 34324 12544
rect 34260 12484 34264 12540
rect 34264 12484 34320 12540
rect 34320 12484 34324 12540
rect 34260 12480 34324 12484
rect 10400 11996 10464 12000
rect 10400 11940 10404 11996
rect 10404 11940 10460 11996
rect 10460 11940 10464 11996
rect 10400 11936 10464 11940
rect 10480 11996 10544 12000
rect 10480 11940 10484 11996
rect 10484 11940 10540 11996
rect 10540 11940 10544 11996
rect 10480 11936 10544 11940
rect 10560 11996 10624 12000
rect 10560 11940 10564 11996
rect 10564 11940 10620 11996
rect 10620 11940 10624 11996
rect 10560 11936 10624 11940
rect 10640 11996 10704 12000
rect 10640 11940 10644 11996
rect 10644 11940 10700 11996
rect 10700 11940 10704 11996
rect 10640 11936 10704 11940
rect 19848 11996 19912 12000
rect 19848 11940 19852 11996
rect 19852 11940 19908 11996
rect 19908 11940 19912 11996
rect 19848 11936 19912 11940
rect 19928 11996 19992 12000
rect 19928 11940 19932 11996
rect 19932 11940 19988 11996
rect 19988 11940 19992 11996
rect 19928 11936 19992 11940
rect 20008 11996 20072 12000
rect 20008 11940 20012 11996
rect 20012 11940 20068 11996
rect 20068 11940 20072 11996
rect 20008 11936 20072 11940
rect 20088 11996 20152 12000
rect 20088 11940 20092 11996
rect 20092 11940 20148 11996
rect 20148 11940 20152 11996
rect 20088 11936 20152 11940
rect 29296 11996 29360 12000
rect 29296 11940 29300 11996
rect 29300 11940 29356 11996
rect 29356 11940 29360 11996
rect 29296 11936 29360 11940
rect 29376 11996 29440 12000
rect 29376 11940 29380 11996
rect 29380 11940 29436 11996
rect 29436 11940 29440 11996
rect 29376 11936 29440 11940
rect 29456 11996 29520 12000
rect 29456 11940 29460 11996
rect 29460 11940 29516 11996
rect 29516 11940 29520 11996
rect 29456 11936 29520 11940
rect 29536 11996 29600 12000
rect 29536 11940 29540 11996
rect 29540 11940 29596 11996
rect 29596 11940 29600 11996
rect 29536 11936 29600 11940
rect 5676 11452 5740 11456
rect 5676 11396 5680 11452
rect 5680 11396 5736 11452
rect 5736 11396 5740 11452
rect 5676 11392 5740 11396
rect 5756 11452 5820 11456
rect 5756 11396 5760 11452
rect 5760 11396 5816 11452
rect 5816 11396 5820 11452
rect 5756 11392 5820 11396
rect 5836 11452 5900 11456
rect 5836 11396 5840 11452
rect 5840 11396 5896 11452
rect 5896 11396 5900 11452
rect 5836 11392 5900 11396
rect 5916 11452 5980 11456
rect 5916 11396 5920 11452
rect 5920 11396 5976 11452
rect 5976 11396 5980 11452
rect 5916 11392 5980 11396
rect 15124 11452 15188 11456
rect 15124 11396 15128 11452
rect 15128 11396 15184 11452
rect 15184 11396 15188 11452
rect 15124 11392 15188 11396
rect 15204 11452 15268 11456
rect 15204 11396 15208 11452
rect 15208 11396 15264 11452
rect 15264 11396 15268 11452
rect 15204 11392 15268 11396
rect 15284 11452 15348 11456
rect 15284 11396 15288 11452
rect 15288 11396 15344 11452
rect 15344 11396 15348 11452
rect 15284 11392 15348 11396
rect 15364 11452 15428 11456
rect 15364 11396 15368 11452
rect 15368 11396 15424 11452
rect 15424 11396 15428 11452
rect 15364 11392 15428 11396
rect 24572 11452 24636 11456
rect 24572 11396 24576 11452
rect 24576 11396 24632 11452
rect 24632 11396 24636 11452
rect 24572 11392 24636 11396
rect 24652 11452 24716 11456
rect 24652 11396 24656 11452
rect 24656 11396 24712 11452
rect 24712 11396 24716 11452
rect 24652 11392 24716 11396
rect 24732 11452 24796 11456
rect 24732 11396 24736 11452
rect 24736 11396 24792 11452
rect 24792 11396 24796 11452
rect 24732 11392 24796 11396
rect 24812 11452 24876 11456
rect 24812 11396 24816 11452
rect 24816 11396 24872 11452
rect 24872 11396 24876 11452
rect 24812 11392 24876 11396
rect 34020 11452 34084 11456
rect 34020 11396 34024 11452
rect 34024 11396 34080 11452
rect 34080 11396 34084 11452
rect 34020 11392 34084 11396
rect 34100 11452 34164 11456
rect 34100 11396 34104 11452
rect 34104 11396 34160 11452
rect 34160 11396 34164 11452
rect 34100 11392 34164 11396
rect 34180 11452 34244 11456
rect 34180 11396 34184 11452
rect 34184 11396 34240 11452
rect 34240 11396 34244 11452
rect 34180 11392 34244 11396
rect 34260 11452 34324 11456
rect 34260 11396 34264 11452
rect 34264 11396 34320 11452
rect 34320 11396 34324 11452
rect 34260 11392 34324 11396
rect 10400 10908 10464 10912
rect 10400 10852 10404 10908
rect 10404 10852 10460 10908
rect 10460 10852 10464 10908
rect 10400 10848 10464 10852
rect 10480 10908 10544 10912
rect 10480 10852 10484 10908
rect 10484 10852 10540 10908
rect 10540 10852 10544 10908
rect 10480 10848 10544 10852
rect 10560 10908 10624 10912
rect 10560 10852 10564 10908
rect 10564 10852 10620 10908
rect 10620 10852 10624 10908
rect 10560 10848 10624 10852
rect 10640 10908 10704 10912
rect 10640 10852 10644 10908
rect 10644 10852 10700 10908
rect 10700 10852 10704 10908
rect 10640 10848 10704 10852
rect 19848 10908 19912 10912
rect 19848 10852 19852 10908
rect 19852 10852 19908 10908
rect 19908 10852 19912 10908
rect 19848 10848 19912 10852
rect 19928 10908 19992 10912
rect 19928 10852 19932 10908
rect 19932 10852 19988 10908
rect 19988 10852 19992 10908
rect 19928 10848 19992 10852
rect 20008 10908 20072 10912
rect 20008 10852 20012 10908
rect 20012 10852 20068 10908
rect 20068 10852 20072 10908
rect 20008 10848 20072 10852
rect 20088 10908 20152 10912
rect 20088 10852 20092 10908
rect 20092 10852 20148 10908
rect 20148 10852 20152 10908
rect 20088 10848 20152 10852
rect 29296 10908 29360 10912
rect 29296 10852 29300 10908
rect 29300 10852 29356 10908
rect 29356 10852 29360 10908
rect 29296 10848 29360 10852
rect 29376 10908 29440 10912
rect 29376 10852 29380 10908
rect 29380 10852 29436 10908
rect 29436 10852 29440 10908
rect 29376 10848 29440 10852
rect 29456 10908 29520 10912
rect 29456 10852 29460 10908
rect 29460 10852 29516 10908
rect 29516 10852 29520 10908
rect 29456 10848 29520 10852
rect 29536 10908 29600 10912
rect 29536 10852 29540 10908
rect 29540 10852 29596 10908
rect 29596 10852 29600 10908
rect 29536 10848 29600 10852
rect 5676 10364 5740 10368
rect 5676 10308 5680 10364
rect 5680 10308 5736 10364
rect 5736 10308 5740 10364
rect 5676 10304 5740 10308
rect 5756 10364 5820 10368
rect 5756 10308 5760 10364
rect 5760 10308 5816 10364
rect 5816 10308 5820 10364
rect 5756 10304 5820 10308
rect 5836 10364 5900 10368
rect 5836 10308 5840 10364
rect 5840 10308 5896 10364
rect 5896 10308 5900 10364
rect 5836 10304 5900 10308
rect 5916 10364 5980 10368
rect 5916 10308 5920 10364
rect 5920 10308 5976 10364
rect 5976 10308 5980 10364
rect 5916 10304 5980 10308
rect 15124 10364 15188 10368
rect 15124 10308 15128 10364
rect 15128 10308 15184 10364
rect 15184 10308 15188 10364
rect 15124 10304 15188 10308
rect 15204 10364 15268 10368
rect 15204 10308 15208 10364
rect 15208 10308 15264 10364
rect 15264 10308 15268 10364
rect 15204 10304 15268 10308
rect 15284 10364 15348 10368
rect 15284 10308 15288 10364
rect 15288 10308 15344 10364
rect 15344 10308 15348 10364
rect 15284 10304 15348 10308
rect 15364 10364 15428 10368
rect 15364 10308 15368 10364
rect 15368 10308 15424 10364
rect 15424 10308 15428 10364
rect 15364 10304 15428 10308
rect 24572 10364 24636 10368
rect 24572 10308 24576 10364
rect 24576 10308 24632 10364
rect 24632 10308 24636 10364
rect 24572 10304 24636 10308
rect 24652 10364 24716 10368
rect 24652 10308 24656 10364
rect 24656 10308 24712 10364
rect 24712 10308 24716 10364
rect 24652 10304 24716 10308
rect 24732 10364 24796 10368
rect 24732 10308 24736 10364
rect 24736 10308 24792 10364
rect 24792 10308 24796 10364
rect 24732 10304 24796 10308
rect 24812 10364 24876 10368
rect 24812 10308 24816 10364
rect 24816 10308 24872 10364
rect 24872 10308 24876 10364
rect 24812 10304 24876 10308
rect 34020 10364 34084 10368
rect 34020 10308 34024 10364
rect 34024 10308 34080 10364
rect 34080 10308 34084 10364
rect 34020 10304 34084 10308
rect 34100 10364 34164 10368
rect 34100 10308 34104 10364
rect 34104 10308 34160 10364
rect 34160 10308 34164 10364
rect 34100 10304 34164 10308
rect 34180 10364 34244 10368
rect 34180 10308 34184 10364
rect 34184 10308 34240 10364
rect 34240 10308 34244 10364
rect 34180 10304 34244 10308
rect 34260 10364 34324 10368
rect 34260 10308 34264 10364
rect 34264 10308 34320 10364
rect 34320 10308 34324 10364
rect 34260 10304 34324 10308
rect 10400 9820 10464 9824
rect 10400 9764 10404 9820
rect 10404 9764 10460 9820
rect 10460 9764 10464 9820
rect 10400 9760 10464 9764
rect 10480 9820 10544 9824
rect 10480 9764 10484 9820
rect 10484 9764 10540 9820
rect 10540 9764 10544 9820
rect 10480 9760 10544 9764
rect 10560 9820 10624 9824
rect 10560 9764 10564 9820
rect 10564 9764 10620 9820
rect 10620 9764 10624 9820
rect 10560 9760 10624 9764
rect 10640 9820 10704 9824
rect 10640 9764 10644 9820
rect 10644 9764 10700 9820
rect 10700 9764 10704 9820
rect 10640 9760 10704 9764
rect 19848 9820 19912 9824
rect 19848 9764 19852 9820
rect 19852 9764 19908 9820
rect 19908 9764 19912 9820
rect 19848 9760 19912 9764
rect 19928 9820 19992 9824
rect 19928 9764 19932 9820
rect 19932 9764 19988 9820
rect 19988 9764 19992 9820
rect 19928 9760 19992 9764
rect 20008 9820 20072 9824
rect 20008 9764 20012 9820
rect 20012 9764 20068 9820
rect 20068 9764 20072 9820
rect 20008 9760 20072 9764
rect 20088 9820 20152 9824
rect 20088 9764 20092 9820
rect 20092 9764 20148 9820
rect 20148 9764 20152 9820
rect 20088 9760 20152 9764
rect 29296 9820 29360 9824
rect 29296 9764 29300 9820
rect 29300 9764 29356 9820
rect 29356 9764 29360 9820
rect 29296 9760 29360 9764
rect 29376 9820 29440 9824
rect 29376 9764 29380 9820
rect 29380 9764 29436 9820
rect 29436 9764 29440 9820
rect 29376 9760 29440 9764
rect 29456 9820 29520 9824
rect 29456 9764 29460 9820
rect 29460 9764 29516 9820
rect 29516 9764 29520 9820
rect 29456 9760 29520 9764
rect 29536 9820 29600 9824
rect 29536 9764 29540 9820
rect 29540 9764 29596 9820
rect 29596 9764 29600 9820
rect 29536 9760 29600 9764
rect 5676 9276 5740 9280
rect 5676 9220 5680 9276
rect 5680 9220 5736 9276
rect 5736 9220 5740 9276
rect 5676 9216 5740 9220
rect 5756 9276 5820 9280
rect 5756 9220 5760 9276
rect 5760 9220 5816 9276
rect 5816 9220 5820 9276
rect 5756 9216 5820 9220
rect 5836 9276 5900 9280
rect 5836 9220 5840 9276
rect 5840 9220 5896 9276
rect 5896 9220 5900 9276
rect 5836 9216 5900 9220
rect 5916 9276 5980 9280
rect 5916 9220 5920 9276
rect 5920 9220 5976 9276
rect 5976 9220 5980 9276
rect 5916 9216 5980 9220
rect 15124 9276 15188 9280
rect 15124 9220 15128 9276
rect 15128 9220 15184 9276
rect 15184 9220 15188 9276
rect 15124 9216 15188 9220
rect 15204 9276 15268 9280
rect 15204 9220 15208 9276
rect 15208 9220 15264 9276
rect 15264 9220 15268 9276
rect 15204 9216 15268 9220
rect 15284 9276 15348 9280
rect 15284 9220 15288 9276
rect 15288 9220 15344 9276
rect 15344 9220 15348 9276
rect 15284 9216 15348 9220
rect 15364 9276 15428 9280
rect 15364 9220 15368 9276
rect 15368 9220 15424 9276
rect 15424 9220 15428 9276
rect 15364 9216 15428 9220
rect 24572 9276 24636 9280
rect 24572 9220 24576 9276
rect 24576 9220 24632 9276
rect 24632 9220 24636 9276
rect 24572 9216 24636 9220
rect 24652 9276 24716 9280
rect 24652 9220 24656 9276
rect 24656 9220 24712 9276
rect 24712 9220 24716 9276
rect 24652 9216 24716 9220
rect 24732 9276 24796 9280
rect 24732 9220 24736 9276
rect 24736 9220 24792 9276
rect 24792 9220 24796 9276
rect 24732 9216 24796 9220
rect 24812 9276 24876 9280
rect 24812 9220 24816 9276
rect 24816 9220 24872 9276
rect 24872 9220 24876 9276
rect 24812 9216 24876 9220
rect 34020 9276 34084 9280
rect 34020 9220 34024 9276
rect 34024 9220 34080 9276
rect 34080 9220 34084 9276
rect 34020 9216 34084 9220
rect 34100 9276 34164 9280
rect 34100 9220 34104 9276
rect 34104 9220 34160 9276
rect 34160 9220 34164 9276
rect 34100 9216 34164 9220
rect 34180 9276 34244 9280
rect 34180 9220 34184 9276
rect 34184 9220 34240 9276
rect 34240 9220 34244 9276
rect 34180 9216 34244 9220
rect 34260 9276 34324 9280
rect 34260 9220 34264 9276
rect 34264 9220 34320 9276
rect 34320 9220 34324 9276
rect 34260 9216 34324 9220
rect 10400 8732 10464 8736
rect 10400 8676 10404 8732
rect 10404 8676 10460 8732
rect 10460 8676 10464 8732
rect 10400 8672 10464 8676
rect 10480 8732 10544 8736
rect 10480 8676 10484 8732
rect 10484 8676 10540 8732
rect 10540 8676 10544 8732
rect 10480 8672 10544 8676
rect 10560 8732 10624 8736
rect 10560 8676 10564 8732
rect 10564 8676 10620 8732
rect 10620 8676 10624 8732
rect 10560 8672 10624 8676
rect 10640 8732 10704 8736
rect 10640 8676 10644 8732
rect 10644 8676 10700 8732
rect 10700 8676 10704 8732
rect 10640 8672 10704 8676
rect 19848 8732 19912 8736
rect 19848 8676 19852 8732
rect 19852 8676 19908 8732
rect 19908 8676 19912 8732
rect 19848 8672 19912 8676
rect 19928 8732 19992 8736
rect 19928 8676 19932 8732
rect 19932 8676 19988 8732
rect 19988 8676 19992 8732
rect 19928 8672 19992 8676
rect 20008 8732 20072 8736
rect 20008 8676 20012 8732
rect 20012 8676 20068 8732
rect 20068 8676 20072 8732
rect 20008 8672 20072 8676
rect 20088 8732 20152 8736
rect 20088 8676 20092 8732
rect 20092 8676 20148 8732
rect 20148 8676 20152 8732
rect 20088 8672 20152 8676
rect 29296 8732 29360 8736
rect 29296 8676 29300 8732
rect 29300 8676 29356 8732
rect 29356 8676 29360 8732
rect 29296 8672 29360 8676
rect 29376 8732 29440 8736
rect 29376 8676 29380 8732
rect 29380 8676 29436 8732
rect 29436 8676 29440 8732
rect 29376 8672 29440 8676
rect 29456 8732 29520 8736
rect 29456 8676 29460 8732
rect 29460 8676 29516 8732
rect 29516 8676 29520 8732
rect 29456 8672 29520 8676
rect 29536 8732 29600 8736
rect 29536 8676 29540 8732
rect 29540 8676 29596 8732
rect 29596 8676 29600 8732
rect 29536 8672 29600 8676
rect 5676 8188 5740 8192
rect 5676 8132 5680 8188
rect 5680 8132 5736 8188
rect 5736 8132 5740 8188
rect 5676 8128 5740 8132
rect 5756 8188 5820 8192
rect 5756 8132 5760 8188
rect 5760 8132 5816 8188
rect 5816 8132 5820 8188
rect 5756 8128 5820 8132
rect 5836 8188 5900 8192
rect 5836 8132 5840 8188
rect 5840 8132 5896 8188
rect 5896 8132 5900 8188
rect 5836 8128 5900 8132
rect 5916 8188 5980 8192
rect 5916 8132 5920 8188
rect 5920 8132 5976 8188
rect 5976 8132 5980 8188
rect 5916 8128 5980 8132
rect 15124 8188 15188 8192
rect 15124 8132 15128 8188
rect 15128 8132 15184 8188
rect 15184 8132 15188 8188
rect 15124 8128 15188 8132
rect 15204 8188 15268 8192
rect 15204 8132 15208 8188
rect 15208 8132 15264 8188
rect 15264 8132 15268 8188
rect 15204 8128 15268 8132
rect 15284 8188 15348 8192
rect 15284 8132 15288 8188
rect 15288 8132 15344 8188
rect 15344 8132 15348 8188
rect 15284 8128 15348 8132
rect 15364 8188 15428 8192
rect 15364 8132 15368 8188
rect 15368 8132 15424 8188
rect 15424 8132 15428 8188
rect 15364 8128 15428 8132
rect 24572 8188 24636 8192
rect 24572 8132 24576 8188
rect 24576 8132 24632 8188
rect 24632 8132 24636 8188
rect 24572 8128 24636 8132
rect 24652 8188 24716 8192
rect 24652 8132 24656 8188
rect 24656 8132 24712 8188
rect 24712 8132 24716 8188
rect 24652 8128 24716 8132
rect 24732 8188 24796 8192
rect 24732 8132 24736 8188
rect 24736 8132 24792 8188
rect 24792 8132 24796 8188
rect 24732 8128 24796 8132
rect 24812 8188 24876 8192
rect 24812 8132 24816 8188
rect 24816 8132 24872 8188
rect 24872 8132 24876 8188
rect 24812 8128 24876 8132
rect 34020 8188 34084 8192
rect 34020 8132 34024 8188
rect 34024 8132 34080 8188
rect 34080 8132 34084 8188
rect 34020 8128 34084 8132
rect 34100 8188 34164 8192
rect 34100 8132 34104 8188
rect 34104 8132 34160 8188
rect 34160 8132 34164 8188
rect 34100 8128 34164 8132
rect 34180 8188 34244 8192
rect 34180 8132 34184 8188
rect 34184 8132 34240 8188
rect 34240 8132 34244 8188
rect 34180 8128 34244 8132
rect 34260 8188 34324 8192
rect 34260 8132 34264 8188
rect 34264 8132 34320 8188
rect 34320 8132 34324 8188
rect 34260 8128 34324 8132
rect 10400 7644 10464 7648
rect 10400 7588 10404 7644
rect 10404 7588 10460 7644
rect 10460 7588 10464 7644
rect 10400 7584 10464 7588
rect 10480 7644 10544 7648
rect 10480 7588 10484 7644
rect 10484 7588 10540 7644
rect 10540 7588 10544 7644
rect 10480 7584 10544 7588
rect 10560 7644 10624 7648
rect 10560 7588 10564 7644
rect 10564 7588 10620 7644
rect 10620 7588 10624 7644
rect 10560 7584 10624 7588
rect 10640 7644 10704 7648
rect 10640 7588 10644 7644
rect 10644 7588 10700 7644
rect 10700 7588 10704 7644
rect 10640 7584 10704 7588
rect 19848 7644 19912 7648
rect 19848 7588 19852 7644
rect 19852 7588 19908 7644
rect 19908 7588 19912 7644
rect 19848 7584 19912 7588
rect 19928 7644 19992 7648
rect 19928 7588 19932 7644
rect 19932 7588 19988 7644
rect 19988 7588 19992 7644
rect 19928 7584 19992 7588
rect 20008 7644 20072 7648
rect 20008 7588 20012 7644
rect 20012 7588 20068 7644
rect 20068 7588 20072 7644
rect 20008 7584 20072 7588
rect 20088 7644 20152 7648
rect 20088 7588 20092 7644
rect 20092 7588 20148 7644
rect 20148 7588 20152 7644
rect 20088 7584 20152 7588
rect 29296 7644 29360 7648
rect 29296 7588 29300 7644
rect 29300 7588 29356 7644
rect 29356 7588 29360 7644
rect 29296 7584 29360 7588
rect 29376 7644 29440 7648
rect 29376 7588 29380 7644
rect 29380 7588 29436 7644
rect 29436 7588 29440 7644
rect 29376 7584 29440 7588
rect 29456 7644 29520 7648
rect 29456 7588 29460 7644
rect 29460 7588 29516 7644
rect 29516 7588 29520 7644
rect 29456 7584 29520 7588
rect 29536 7644 29600 7648
rect 29536 7588 29540 7644
rect 29540 7588 29596 7644
rect 29596 7588 29600 7644
rect 29536 7584 29600 7588
rect 5676 7100 5740 7104
rect 5676 7044 5680 7100
rect 5680 7044 5736 7100
rect 5736 7044 5740 7100
rect 5676 7040 5740 7044
rect 5756 7100 5820 7104
rect 5756 7044 5760 7100
rect 5760 7044 5816 7100
rect 5816 7044 5820 7100
rect 5756 7040 5820 7044
rect 5836 7100 5900 7104
rect 5836 7044 5840 7100
rect 5840 7044 5896 7100
rect 5896 7044 5900 7100
rect 5836 7040 5900 7044
rect 5916 7100 5980 7104
rect 5916 7044 5920 7100
rect 5920 7044 5976 7100
rect 5976 7044 5980 7100
rect 5916 7040 5980 7044
rect 15124 7100 15188 7104
rect 15124 7044 15128 7100
rect 15128 7044 15184 7100
rect 15184 7044 15188 7100
rect 15124 7040 15188 7044
rect 15204 7100 15268 7104
rect 15204 7044 15208 7100
rect 15208 7044 15264 7100
rect 15264 7044 15268 7100
rect 15204 7040 15268 7044
rect 15284 7100 15348 7104
rect 15284 7044 15288 7100
rect 15288 7044 15344 7100
rect 15344 7044 15348 7100
rect 15284 7040 15348 7044
rect 15364 7100 15428 7104
rect 15364 7044 15368 7100
rect 15368 7044 15424 7100
rect 15424 7044 15428 7100
rect 15364 7040 15428 7044
rect 24572 7100 24636 7104
rect 24572 7044 24576 7100
rect 24576 7044 24632 7100
rect 24632 7044 24636 7100
rect 24572 7040 24636 7044
rect 24652 7100 24716 7104
rect 24652 7044 24656 7100
rect 24656 7044 24712 7100
rect 24712 7044 24716 7100
rect 24652 7040 24716 7044
rect 24732 7100 24796 7104
rect 24732 7044 24736 7100
rect 24736 7044 24792 7100
rect 24792 7044 24796 7100
rect 24732 7040 24796 7044
rect 24812 7100 24876 7104
rect 24812 7044 24816 7100
rect 24816 7044 24872 7100
rect 24872 7044 24876 7100
rect 24812 7040 24876 7044
rect 34020 7100 34084 7104
rect 34020 7044 34024 7100
rect 34024 7044 34080 7100
rect 34080 7044 34084 7100
rect 34020 7040 34084 7044
rect 34100 7100 34164 7104
rect 34100 7044 34104 7100
rect 34104 7044 34160 7100
rect 34160 7044 34164 7100
rect 34100 7040 34164 7044
rect 34180 7100 34244 7104
rect 34180 7044 34184 7100
rect 34184 7044 34240 7100
rect 34240 7044 34244 7100
rect 34180 7040 34244 7044
rect 34260 7100 34324 7104
rect 34260 7044 34264 7100
rect 34264 7044 34320 7100
rect 34320 7044 34324 7100
rect 34260 7040 34324 7044
rect 10400 6556 10464 6560
rect 10400 6500 10404 6556
rect 10404 6500 10460 6556
rect 10460 6500 10464 6556
rect 10400 6496 10464 6500
rect 10480 6556 10544 6560
rect 10480 6500 10484 6556
rect 10484 6500 10540 6556
rect 10540 6500 10544 6556
rect 10480 6496 10544 6500
rect 10560 6556 10624 6560
rect 10560 6500 10564 6556
rect 10564 6500 10620 6556
rect 10620 6500 10624 6556
rect 10560 6496 10624 6500
rect 10640 6556 10704 6560
rect 10640 6500 10644 6556
rect 10644 6500 10700 6556
rect 10700 6500 10704 6556
rect 10640 6496 10704 6500
rect 19848 6556 19912 6560
rect 19848 6500 19852 6556
rect 19852 6500 19908 6556
rect 19908 6500 19912 6556
rect 19848 6496 19912 6500
rect 19928 6556 19992 6560
rect 19928 6500 19932 6556
rect 19932 6500 19988 6556
rect 19988 6500 19992 6556
rect 19928 6496 19992 6500
rect 20008 6556 20072 6560
rect 20008 6500 20012 6556
rect 20012 6500 20068 6556
rect 20068 6500 20072 6556
rect 20008 6496 20072 6500
rect 20088 6556 20152 6560
rect 20088 6500 20092 6556
rect 20092 6500 20148 6556
rect 20148 6500 20152 6556
rect 20088 6496 20152 6500
rect 29296 6556 29360 6560
rect 29296 6500 29300 6556
rect 29300 6500 29356 6556
rect 29356 6500 29360 6556
rect 29296 6496 29360 6500
rect 29376 6556 29440 6560
rect 29376 6500 29380 6556
rect 29380 6500 29436 6556
rect 29436 6500 29440 6556
rect 29376 6496 29440 6500
rect 29456 6556 29520 6560
rect 29456 6500 29460 6556
rect 29460 6500 29516 6556
rect 29516 6500 29520 6556
rect 29456 6496 29520 6500
rect 29536 6556 29600 6560
rect 29536 6500 29540 6556
rect 29540 6500 29596 6556
rect 29596 6500 29600 6556
rect 29536 6496 29600 6500
rect 5676 6012 5740 6016
rect 5676 5956 5680 6012
rect 5680 5956 5736 6012
rect 5736 5956 5740 6012
rect 5676 5952 5740 5956
rect 5756 6012 5820 6016
rect 5756 5956 5760 6012
rect 5760 5956 5816 6012
rect 5816 5956 5820 6012
rect 5756 5952 5820 5956
rect 5836 6012 5900 6016
rect 5836 5956 5840 6012
rect 5840 5956 5896 6012
rect 5896 5956 5900 6012
rect 5836 5952 5900 5956
rect 5916 6012 5980 6016
rect 5916 5956 5920 6012
rect 5920 5956 5976 6012
rect 5976 5956 5980 6012
rect 5916 5952 5980 5956
rect 15124 6012 15188 6016
rect 15124 5956 15128 6012
rect 15128 5956 15184 6012
rect 15184 5956 15188 6012
rect 15124 5952 15188 5956
rect 15204 6012 15268 6016
rect 15204 5956 15208 6012
rect 15208 5956 15264 6012
rect 15264 5956 15268 6012
rect 15204 5952 15268 5956
rect 15284 6012 15348 6016
rect 15284 5956 15288 6012
rect 15288 5956 15344 6012
rect 15344 5956 15348 6012
rect 15284 5952 15348 5956
rect 15364 6012 15428 6016
rect 15364 5956 15368 6012
rect 15368 5956 15424 6012
rect 15424 5956 15428 6012
rect 15364 5952 15428 5956
rect 24572 6012 24636 6016
rect 24572 5956 24576 6012
rect 24576 5956 24632 6012
rect 24632 5956 24636 6012
rect 24572 5952 24636 5956
rect 24652 6012 24716 6016
rect 24652 5956 24656 6012
rect 24656 5956 24712 6012
rect 24712 5956 24716 6012
rect 24652 5952 24716 5956
rect 24732 6012 24796 6016
rect 24732 5956 24736 6012
rect 24736 5956 24792 6012
rect 24792 5956 24796 6012
rect 24732 5952 24796 5956
rect 24812 6012 24876 6016
rect 24812 5956 24816 6012
rect 24816 5956 24872 6012
rect 24872 5956 24876 6012
rect 24812 5952 24876 5956
rect 34020 6012 34084 6016
rect 34020 5956 34024 6012
rect 34024 5956 34080 6012
rect 34080 5956 34084 6012
rect 34020 5952 34084 5956
rect 34100 6012 34164 6016
rect 34100 5956 34104 6012
rect 34104 5956 34160 6012
rect 34160 5956 34164 6012
rect 34100 5952 34164 5956
rect 34180 6012 34244 6016
rect 34180 5956 34184 6012
rect 34184 5956 34240 6012
rect 34240 5956 34244 6012
rect 34180 5952 34244 5956
rect 34260 6012 34324 6016
rect 34260 5956 34264 6012
rect 34264 5956 34320 6012
rect 34320 5956 34324 6012
rect 34260 5952 34324 5956
rect 10400 5468 10464 5472
rect 10400 5412 10404 5468
rect 10404 5412 10460 5468
rect 10460 5412 10464 5468
rect 10400 5408 10464 5412
rect 10480 5468 10544 5472
rect 10480 5412 10484 5468
rect 10484 5412 10540 5468
rect 10540 5412 10544 5468
rect 10480 5408 10544 5412
rect 10560 5468 10624 5472
rect 10560 5412 10564 5468
rect 10564 5412 10620 5468
rect 10620 5412 10624 5468
rect 10560 5408 10624 5412
rect 10640 5468 10704 5472
rect 10640 5412 10644 5468
rect 10644 5412 10700 5468
rect 10700 5412 10704 5468
rect 10640 5408 10704 5412
rect 19848 5468 19912 5472
rect 19848 5412 19852 5468
rect 19852 5412 19908 5468
rect 19908 5412 19912 5468
rect 19848 5408 19912 5412
rect 19928 5468 19992 5472
rect 19928 5412 19932 5468
rect 19932 5412 19988 5468
rect 19988 5412 19992 5468
rect 19928 5408 19992 5412
rect 20008 5468 20072 5472
rect 20008 5412 20012 5468
rect 20012 5412 20068 5468
rect 20068 5412 20072 5468
rect 20008 5408 20072 5412
rect 20088 5468 20152 5472
rect 20088 5412 20092 5468
rect 20092 5412 20148 5468
rect 20148 5412 20152 5468
rect 20088 5408 20152 5412
rect 29296 5468 29360 5472
rect 29296 5412 29300 5468
rect 29300 5412 29356 5468
rect 29356 5412 29360 5468
rect 29296 5408 29360 5412
rect 29376 5468 29440 5472
rect 29376 5412 29380 5468
rect 29380 5412 29436 5468
rect 29436 5412 29440 5468
rect 29376 5408 29440 5412
rect 29456 5468 29520 5472
rect 29456 5412 29460 5468
rect 29460 5412 29516 5468
rect 29516 5412 29520 5468
rect 29456 5408 29520 5412
rect 29536 5468 29600 5472
rect 29536 5412 29540 5468
rect 29540 5412 29596 5468
rect 29596 5412 29600 5468
rect 29536 5408 29600 5412
rect 5676 4924 5740 4928
rect 5676 4868 5680 4924
rect 5680 4868 5736 4924
rect 5736 4868 5740 4924
rect 5676 4864 5740 4868
rect 5756 4924 5820 4928
rect 5756 4868 5760 4924
rect 5760 4868 5816 4924
rect 5816 4868 5820 4924
rect 5756 4864 5820 4868
rect 5836 4924 5900 4928
rect 5836 4868 5840 4924
rect 5840 4868 5896 4924
rect 5896 4868 5900 4924
rect 5836 4864 5900 4868
rect 5916 4924 5980 4928
rect 5916 4868 5920 4924
rect 5920 4868 5976 4924
rect 5976 4868 5980 4924
rect 5916 4864 5980 4868
rect 15124 4924 15188 4928
rect 15124 4868 15128 4924
rect 15128 4868 15184 4924
rect 15184 4868 15188 4924
rect 15124 4864 15188 4868
rect 15204 4924 15268 4928
rect 15204 4868 15208 4924
rect 15208 4868 15264 4924
rect 15264 4868 15268 4924
rect 15204 4864 15268 4868
rect 15284 4924 15348 4928
rect 15284 4868 15288 4924
rect 15288 4868 15344 4924
rect 15344 4868 15348 4924
rect 15284 4864 15348 4868
rect 15364 4924 15428 4928
rect 15364 4868 15368 4924
rect 15368 4868 15424 4924
rect 15424 4868 15428 4924
rect 15364 4864 15428 4868
rect 24572 4924 24636 4928
rect 24572 4868 24576 4924
rect 24576 4868 24632 4924
rect 24632 4868 24636 4924
rect 24572 4864 24636 4868
rect 24652 4924 24716 4928
rect 24652 4868 24656 4924
rect 24656 4868 24712 4924
rect 24712 4868 24716 4924
rect 24652 4864 24716 4868
rect 24732 4924 24796 4928
rect 24732 4868 24736 4924
rect 24736 4868 24792 4924
rect 24792 4868 24796 4924
rect 24732 4864 24796 4868
rect 24812 4924 24876 4928
rect 24812 4868 24816 4924
rect 24816 4868 24872 4924
rect 24872 4868 24876 4924
rect 24812 4864 24876 4868
rect 34020 4924 34084 4928
rect 34020 4868 34024 4924
rect 34024 4868 34080 4924
rect 34080 4868 34084 4924
rect 34020 4864 34084 4868
rect 34100 4924 34164 4928
rect 34100 4868 34104 4924
rect 34104 4868 34160 4924
rect 34160 4868 34164 4924
rect 34100 4864 34164 4868
rect 34180 4924 34244 4928
rect 34180 4868 34184 4924
rect 34184 4868 34240 4924
rect 34240 4868 34244 4924
rect 34180 4864 34244 4868
rect 34260 4924 34324 4928
rect 34260 4868 34264 4924
rect 34264 4868 34320 4924
rect 34320 4868 34324 4924
rect 34260 4864 34324 4868
rect 10400 4380 10464 4384
rect 10400 4324 10404 4380
rect 10404 4324 10460 4380
rect 10460 4324 10464 4380
rect 10400 4320 10464 4324
rect 10480 4380 10544 4384
rect 10480 4324 10484 4380
rect 10484 4324 10540 4380
rect 10540 4324 10544 4380
rect 10480 4320 10544 4324
rect 10560 4380 10624 4384
rect 10560 4324 10564 4380
rect 10564 4324 10620 4380
rect 10620 4324 10624 4380
rect 10560 4320 10624 4324
rect 10640 4380 10704 4384
rect 10640 4324 10644 4380
rect 10644 4324 10700 4380
rect 10700 4324 10704 4380
rect 10640 4320 10704 4324
rect 19848 4380 19912 4384
rect 19848 4324 19852 4380
rect 19852 4324 19908 4380
rect 19908 4324 19912 4380
rect 19848 4320 19912 4324
rect 19928 4380 19992 4384
rect 19928 4324 19932 4380
rect 19932 4324 19988 4380
rect 19988 4324 19992 4380
rect 19928 4320 19992 4324
rect 20008 4380 20072 4384
rect 20008 4324 20012 4380
rect 20012 4324 20068 4380
rect 20068 4324 20072 4380
rect 20008 4320 20072 4324
rect 20088 4380 20152 4384
rect 20088 4324 20092 4380
rect 20092 4324 20148 4380
rect 20148 4324 20152 4380
rect 20088 4320 20152 4324
rect 29296 4380 29360 4384
rect 29296 4324 29300 4380
rect 29300 4324 29356 4380
rect 29356 4324 29360 4380
rect 29296 4320 29360 4324
rect 29376 4380 29440 4384
rect 29376 4324 29380 4380
rect 29380 4324 29436 4380
rect 29436 4324 29440 4380
rect 29376 4320 29440 4324
rect 29456 4380 29520 4384
rect 29456 4324 29460 4380
rect 29460 4324 29516 4380
rect 29516 4324 29520 4380
rect 29456 4320 29520 4324
rect 29536 4380 29600 4384
rect 29536 4324 29540 4380
rect 29540 4324 29596 4380
rect 29596 4324 29600 4380
rect 29536 4320 29600 4324
rect 5676 3836 5740 3840
rect 5676 3780 5680 3836
rect 5680 3780 5736 3836
rect 5736 3780 5740 3836
rect 5676 3776 5740 3780
rect 5756 3836 5820 3840
rect 5756 3780 5760 3836
rect 5760 3780 5816 3836
rect 5816 3780 5820 3836
rect 5756 3776 5820 3780
rect 5836 3836 5900 3840
rect 5836 3780 5840 3836
rect 5840 3780 5896 3836
rect 5896 3780 5900 3836
rect 5836 3776 5900 3780
rect 5916 3836 5980 3840
rect 5916 3780 5920 3836
rect 5920 3780 5976 3836
rect 5976 3780 5980 3836
rect 5916 3776 5980 3780
rect 15124 3836 15188 3840
rect 15124 3780 15128 3836
rect 15128 3780 15184 3836
rect 15184 3780 15188 3836
rect 15124 3776 15188 3780
rect 15204 3836 15268 3840
rect 15204 3780 15208 3836
rect 15208 3780 15264 3836
rect 15264 3780 15268 3836
rect 15204 3776 15268 3780
rect 15284 3836 15348 3840
rect 15284 3780 15288 3836
rect 15288 3780 15344 3836
rect 15344 3780 15348 3836
rect 15284 3776 15348 3780
rect 15364 3836 15428 3840
rect 15364 3780 15368 3836
rect 15368 3780 15424 3836
rect 15424 3780 15428 3836
rect 15364 3776 15428 3780
rect 24572 3836 24636 3840
rect 24572 3780 24576 3836
rect 24576 3780 24632 3836
rect 24632 3780 24636 3836
rect 24572 3776 24636 3780
rect 24652 3836 24716 3840
rect 24652 3780 24656 3836
rect 24656 3780 24712 3836
rect 24712 3780 24716 3836
rect 24652 3776 24716 3780
rect 24732 3836 24796 3840
rect 24732 3780 24736 3836
rect 24736 3780 24792 3836
rect 24792 3780 24796 3836
rect 24732 3776 24796 3780
rect 24812 3836 24876 3840
rect 24812 3780 24816 3836
rect 24816 3780 24872 3836
rect 24872 3780 24876 3836
rect 24812 3776 24876 3780
rect 34020 3836 34084 3840
rect 34020 3780 34024 3836
rect 34024 3780 34080 3836
rect 34080 3780 34084 3836
rect 34020 3776 34084 3780
rect 34100 3836 34164 3840
rect 34100 3780 34104 3836
rect 34104 3780 34160 3836
rect 34160 3780 34164 3836
rect 34100 3776 34164 3780
rect 34180 3836 34244 3840
rect 34180 3780 34184 3836
rect 34184 3780 34240 3836
rect 34240 3780 34244 3836
rect 34180 3776 34244 3780
rect 34260 3836 34324 3840
rect 34260 3780 34264 3836
rect 34264 3780 34320 3836
rect 34320 3780 34324 3836
rect 34260 3776 34324 3780
rect 10400 3292 10464 3296
rect 10400 3236 10404 3292
rect 10404 3236 10460 3292
rect 10460 3236 10464 3292
rect 10400 3232 10464 3236
rect 10480 3292 10544 3296
rect 10480 3236 10484 3292
rect 10484 3236 10540 3292
rect 10540 3236 10544 3292
rect 10480 3232 10544 3236
rect 10560 3292 10624 3296
rect 10560 3236 10564 3292
rect 10564 3236 10620 3292
rect 10620 3236 10624 3292
rect 10560 3232 10624 3236
rect 10640 3292 10704 3296
rect 10640 3236 10644 3292
rect 10644 3236 10700 3292
rect 10700 3236 10704 3292
rect 10640 3232 10704 3236
rect 19848 3292 19912 3296
rect 19848 3236 19852 3292
rect 19852 3236 19908 3292
rect 19908 3236 19912 3292
rect 19848 3232 19912 3236
rect 19928 3292 19992 3296
rect 19928 3236 19932 3292
rect 19932 3236 19988 3292
rect 19988 3236 19992 3292
rect 19928 3232 19992 3236
rect 20008 3292 20072 3296
rect 20008 3236 20012 3292
rect 20012 3236 20068 3292
rect 20068 3236 20072 3292
rect 20008 3232 20072 3236
rect 20088 3292 20152 3296
rect 20088 3236 20092 3292
rect 20092 3236 20148 3292
rect 20148 3236 20152 3292
rect 20088 3232 20152 3236
rect 29296 3292 29360 3296
rect 29296 3236 29300 3292
rect 29300 3236 29356 3292
rect 29356 3236 29360 3292
rect 29296 3232 29360 3236
rect 29376 3292 29440 3296
rect 29376 3236 29380 3292
rect 29380 3236 29436 3292
rect 29436 3236 29440 3292
rect 29376 3232 29440 3236
rect 29456 3292 29520 3296
rect 29456 3236 29460 3292
rect 29460 3236 29516 3292
rect 29516 3236 29520 3292
rect 29456 3232 29520 3236
rect 29536 3292 29600 3296
rect 29536 3236 29540 3292
rect 29540 3236 29596 3292
rect 29596 3236 29600 3292
rect 29536 3232 29600 3236
rect 5676 2748 5740 2752
rect 5676 2692 5680 2748
rect 5680 2692 5736 2748
rect 5736 2692 5740 2748
rect 5676 2688 5740 2692
rect 5756 2748 5820 2752
rect 5756 2692 5760 2748
rect 5760 2692 5816 2748
rect 5816 2692 5820 2748
rect 5756 2688 5820 2692
rect 5836 2748 5900 2752
rect 5836 2692 5840 2748
rect 5840 2692 5896 2748
rect 5896 2692 5900 2748
rect 5836 2688 5900 2692
rect 5916 2748 5980 2752
rect 5916 2692 5920 2748
rect 5920 2692 5976 2748
rect 5976 2692 5980 2748
rect 5916 2688 5980 2692
rect 15124 2748 15188 2752
rect 15124 2692 15128 2748
rect 15128 2692 15184 2748
rect 15184 2692 15188 2748
rect 15124 2688 15188 2692
rect 15204 2748 15268 2752
rect 15204 2692 15208 2748
rect 15208 2692 15264 2748
rect 15264 2692 15268 2748
rect 15204 2688 15268 2692
rect 15284 2748 15348 2752
rect 15284 2692 15288 2748
rect 15288 2692 15344 2748
rect 15344 2692 15348 2748
rect 15284 2688 15348 2692
rect 15364 2748 15428 2752
rect 15364 2692 15368 2748
rect 15368 2692 15424 2748
rect 15424 2692 15428 2748
rect 15364 2688 15428 2692
rect 24572 2748 24636 2752
rect 24572 2692 24576 2748
rect 24576 2692 24632 2748
rect 24632 2692 24636 2748
rect 24572 2688 24636 2692
rect 24652 2748 24716 2752
rect 24652 2692 24656 2748
rect 24656 2692 24712 2748
rect 24712 2692 24716 2748
rect 24652 2688 24716 2692
rect 24732 2748 24796 2752
rect 24732 2692 24736 2748
rect 24736 2692 24792 2748
rect 24792 2692 24796 2748
rect 24732 2688 24796 2692
rect 24812 2748 24876 2752
rect 24812 2692 24816 2748
rect 24816 2692 24872 2748
rect 24872 2692 24876 2748
rect 24812 2688 24876 2692
rect 34020 2748 34084 2752
rect 34020 2692 34024 2748
rect 34024 2692 34080 2748
rect 34080 2692 34084 2748
rect 34020 2688 34084 2692
rect 34100 2748 34164 2752
rect 34100 2692 34104 2748
rect 34104 2692 34160 2748
rect 34160 2692 34164 2748
rect 34100 2688 34164 2692
rect 34180 2748 34244 2752
rect 34180 2692 34184 2748
rect 34184 2692 34240 2748
rect 34240 2692 34244 2748
rect 34180 2688 34244 2692
rect 34260 2748 34324 2752
rect 34260 2692 34264 2748
rect 34264 2692 34320 2748
rect 34320 2692 34324 2748
rect 34260 2688 34324 2692
rect 10400 2204 10464 2208
rect 10400 2148 10404 2204
rect 10404 2148 10460 2204
rect 10460 2148 10464 2204
rect 10400 2144 10464 2148
rect 10480 2204 10544 2208
rect 10480 2148 10484 2204
rect 10484 2148 10540 2204
rect 10540 2148 10544 2204
rect 10480 2144 10544 2148
rect 10560 2204 10624 2208
rect 10560 2148 10564 2204
rect 10564 2148 10620 2204
rect 10620 2148 10624 2204
rect 10560 2144 10624 2148
rect 10640 2204 10704 2208
rect 10640 2148 10644 2204
rect 10644 2148 10700 2204
rect 10700 2148 10704 2204
rect 10640 2144 10704 2148
rect 19848 2204 19912 2208
rect 19848 2148 19852 2204
rect 19852 2148 19908 2204
rect 19908 2148 19912 2204
rect 19848 2144 19912 2148
rect 19928 2204 19992 2208
rect 19928 2148 19932 2204
rect 19932 2148 19988 2204
rect 19988 2148 19992 2204
rect 19928 2144 19992 2148
rect 20008 2204 20072 2208
rect 20008 2148 20012 2204
rect 20012 2148 20068 2204
rect 20068 2148 20072 2204
rect 20008 2144 20072 2148
rect 20088 2204 20152 2208
rect 20088 2148 20092 2204
rect 20092 2148 20148 2204
rect 20148 2148 20152 2204
rect 20088 2144 20152 2148
rect 29296 2204 29360 2208
rect 29296 2148 29300 2204
rect 29300 2148 29356 2204
rect 29356 2148 29360 2204
rect 29296 2144 29360 2148
rect 29376 2204 29440 2208
rect 29376 2148 29380 2204
rect 29380 2148 29436 2204
rect 29436 2148 29440 2204
rect 29376 2144 29440 2148
rect 29456 2204 29520 2208
rect 29456 2148 29460 2204
rect 29460 2148 29516 2204
rect 29516 2148 29520 2204
rect 29456 2144 29520 2148
rect 29536 2204 29600 2208
rect 29536 2148 29540 2204
rect 29540 2148 29596 2204
rect 29596 2148 29600 2204
rect 29536 2144 29600 2148
<< metal4 >>
rect 5668 33216 5988 33776
rect 5668 33152 5676 33216
rect 5740 33152 5756 33216
rect 5820 33152 5836 33216
rect 5900 33152 5916 33216
rect 5980 33152 5988 33216
rect 5668 32128 5988 33152
rect 5668 32064 5676 32128
rect 5740 32064 5756 32128
rect 5820 32064 5836 32128
rect 5900 32064 5916 32128
rect 5980 32064 5988 32128
rect 5668 31040 5988 32064
rect 5668 30976 5676 31040
rect 5740 30976 5756 31040
rect 5820 30976 5836 31040
rect 5900 30976 5916 31040
rect 5980 30976 5988 31040
rect 5668 29952 5988 30976
rect 5668 29888 5676 29952
rect 5740 29888 5756 29952
rect 5820 29888 5836 29952
rect 5900 29888 5916 29952
rect 5980 29888 5988 29952
rect 5668 28864 5988 29888
rect 5668 28800 5676 28864
rect 5740 28800 5756 28864
rect 5820 28800 5836 28864
rect 5900 28800 5916 28864
rect 5980 28800 5988 28864
rect 5668 27776 5988 28800
rect 5668 27712 5676 27776
rect 5740 27712 5756 27776
rect 5820 27712 5836 27776
rect 5900 27712 5916 27776
rect 5980 27712 5988 27776
rect 5668 26688 5988 27712
rect 5668 26624 5676 26688
rect 5740 26624 5756 26688
rect 5820 26624 5836 26688
rect 5900 26624 5916 26688
rect 5980 26624 5988 26688
rect 5668 25600 5988 26624
rect 5668 25536 5676 25600
rect 5740 25536 5756 25600
rect 5820 25536 5836 25600
rect 5900 25536 5916 25600
rect 5980 25536 5988 25600
rect 5668 24512 5988 25536
rect 5668 24448 5676 24512
rect 5740 24448 5756 24512
rect 5820 24448 5836 24512
rect 5900 24448 5916 24512
rect 5980 24448 5988 24512
rect 5668 23424 5988 24448
rect 5668 23360 5676 23424
rect 5740 23360 5756 23424
rect 5820 23360 5836 23424
rect 5900 23360 5916 23424
rect 5980 23360 5988 23424
rect 5668 22336 5988 23360
rect 5668 22272 5676 22336
rect 5740 22272 5756 22336
rect 5820 22272 5836 22336
rect 5900 22272 5916 22336
rect 5980 22272 5988 22336
rect 5668 21248 5988 22272
rect 5668 21184 5676 21248
rect 5740 21184 5756 21248
rect 5820 21184 5836 21248
rect 5900 21184 5916 21248
rect 5980 21184 5988 21248
rect 5668 20160 5988 21184
rect 5668 20096 5676 20160
rect 5740 20096 5756 20160
rect 5820 20096 5836 20160
rect 5900 20096 5916 20160
rect 5980 20096 5988 20160
rect 5668 19072 5988 20096
rect 5668 19008 5676 19072
rect 5740 19008 5756 19072
rect 5820 19008 5836 19072
rect 5900 19008 5916 19072
rect 5980 19008 5988 19072
rect 5668 17984 5988 19008
rect 5668 17920 5676 17984
rect 5740 17920 5756 17984
rect 5820 17920 5836 17984
rect 5900 17920 5916 17984
rect 5980 17920 5988 17984
rect 5668 16896 5988 17920
rect 5668 16832 5676 16896
rect 5740 16832 5756 16896
rect 5820 16832 5836 16896
rect 5900 16832 5916 16896
rect 5980 16832 5988 16896
rect 5668 15808 5988 16832
rect 5668 15744 5676 15808
rect 5740 15744 5756 15808
rect 5820 15744 5836 15808
rect 5900 15744 5916 15808
rect 5980 15744 5988 15808
rect 5668 14720 5988 15744
rect 5668 14656 5676 14720
rect 5740 14656 5756 14720
rect 5820 14656 5836 14720
rect 5900 14656 5916 14720
rect 5980 14656 5988 14720
rect 5668 13632 5988 14656
rect 5668 13568 5676 13632
rect 5740 13568 5756 13632
rect 5820 13568 5836 13632
rect 5900 13568 5916 13632
rect 5980 13568 5988 13632
rect 5668 12544 5988 13568
rect 5668 12480 5676 12544
rect 5740 12480 5756 12544
rect 5820 12480 5836 12544
rect 5900 12480 5916 12544
rect 5980 12480 5988 12544
rect 5668 11456 5988 12480
rect 5668 11392 5676 11456
rect 5740 11392 5756 11456
rect 5820 11392 5836 11456
rect 5900 11392 5916 11456
rect 5980 11392 5988 11456
rect 5668 10368 5988 11392
rect 5668 10304 5676 10368
rect 5740 10304 5756 10368
rect 5820 10304 5836 10368
rect 5900 10304 5916 10368
rect 5980 10304 5988 10368
rect 5668 9280 5988 10304
rect 5668 9216 5676 9280
rect 5740 9216 5756 9280
rect 5820 9216 5836 9280
rect 5900 9216 5916 9280
rect 5980 9216 5988 9280
rect 5668 8192 5988 9216
rect 5668 8128 5676 8192
rect 5740 8128 5756 8192
rect 5820 8128 5836 8192
rect 5900 8128 5916 8192
rect 5980 8128 5988 8192
rect 5668 7104 5988 8128
rect 5668 7040 5676 7104
rect 5740 7040 5756 7104
rect 5820 7040 5836 7104
rect 5900 7040 5916 7104
rect 5980 7040 5988 7104
rect 5668 6016 5988 7040
rect 5668 5952 5676 6016
rect 5740 5952 5756 6016
rect 5820 5952 5836 6016
rect 5900 5952 5916 6016
rect 5980 5952 5988 6016
rect 5668 4928 5988 5952
rect 5668 4864 5676 4928
rect 5740 4864 5756 4928
rect 5820 4864 5836 4928
rect 5900 4864 5916 4928
rect 5980 4864 5988 4928
rect 5668 3840 5988 4864
rect 5668 3776 5676 3840
rect 5740 3776 5756 3840
rect 5820 3776 5836 3840
rect 5900 3776 5916 3840
rect 5980 3776 5988 3840
rect 5668 2752 5988 3776
rect 5668 2688 5676 2752
rect 5740 2688 5756 2752
rect 5820 2688 5836 2752
rect 5900 2688 5916 2752
rect 5980 2688 5988 2752
rect 5668 2128 5988 2688
rect 10392 33760 10712 33776
rect 10392 33696 10400 33760
rect 10464 33696 10480 33760
rect 10544 33696 10560 33760
rect 10624 33696 10640 33760
rect 10704 33696 10712 33760
rect 10392 32672 10712 33696
rect 10392 32608 10400 32672
rect 10464 32608 10480 32672
rect 10544 32608 10560 32672
rect 10624 32608 10640 32672
rect 10704 32608 10712 32672
rect 10392 31584 10712 32608
rect 10392 31520 10400 31584
rect 10464 31520 10480 31584
rect 10544 31520 10560 31584
rect 10624 31520 10640 31584
rect 10704 31520 10712 31584
rect 10392 30496 10712 31520
rect 10392 30432 10400 30496
rect 10464 30432 10480 30496
rect 10544 30432 10560 30496
rect 10624 30432 10640 30496
rect 10704 30432 10712 30496
rect 10392 29408 10712 30432
rect 10392 29344 10400 29408
rect 10464 29344 10480 29408
rect 10544 29344 10560 29408
rect 10624 29344 10640 29408
rect 10704 29344 10712 29408
rect 10392 28320 10712 29344
rect 10392 28256 10400 28320
rect 10464 28256 10480 28320
rect 10544 28256 10560 28320
rect 10624 28256 10640 28320
rect 10704 28256 10712 28320
rect 10392 27232 10712 28256
rect 10392 27168 10400 27232
rect 10464 27168 10480 27232
rect 10544 27168 10560 27232
rect 10624 27168 10640 27232
rect 10704 27168 10712 27232
rect 10392 26144 10712 27168
rect 10392 26080 10400 26144
rect 10464 26080 10480 26144
rect 10544 26080 10560 26144
rect 10624 26080 10640 26144
rect 10704 26080 10712 26144
rect 10392 25056 10712 26080
rect 10392 24992 10400 25056
rect 10464 24992 10480 25056
rect 10544 24992 10560 25056
rect 10624 24992 10640 25056
rect 10704 24992 10712 25056
rect 10392 23968 10712 24992
rect 10392 23904 10400 23968
rect 10464 23904 10480 23968
rect 10544 23904 10560 23968
rect 10624 23904 10640 23968
rect 10704 23904 10712 23968
rect 10392 22880 10712 23904
rect 10392 22816 10400 22880
rect 10464 22816 10480 22880
rect 10544 22816 10560 22880
rect 10624 22816 10640 22880
rect 10704 22816 10712 22880
rect 10392 21792 10712 22816
rect 10392 21728 10400 21792
rect 10464 21728 10480 21792
rect 10544 21728 10560 21792
rect 10624 21728 10640 21792
rect 10704 21728 10712 21792
rect 10392 20704 10712 21728
rect 10392 20640 10400 20704
rect 10464 20640 10480 20704
rect 10544 20640 10560 20704
rect 10624 20640 10640 20704
rect 10704 20640 10712 20704
rect 10392 19616 10712 20640
rect 10392 19552 10400 19616
rect 10464 19552 10480 19616
rect 10544 19552 10560 19616
rect 10624 19552 10640 19616
rect 10704 19552 10712 19616
rect 10392 18528 10712 19552
rect 10392 18464 10400 18528
rect 10464 18464 10480 18528
rect 10544 18464 10560 18528
rect 10624 18464 10640 18528
rect 10704 18464 10712 18528
rect 10392 17440 10712 18464
rect 10392 17376 10400 17440
rect 10464 17376 10480 17440
rect 10544 17376 10560 17440
rect 10624 17376 10640 17440
rect 10704 17376 10712 17440
rect 10392 16352 10712 17376
rect 10392 16288 10400 16352
rect 10464 16288 10480 16352
rect 10544 16288 10560 16352
rect 10624 16288 10640 16352
rect 10704 16288 10712 16352
rect 10392 15264 10712 16288
rect 10392 15200 10400 15264
rect 10464 15200 10480 15264
rect 10544 15200 10560 15264
rect 10624 15200 10640 15264
rect 10704 15200 10712 15264
rect 10392 14176 10712 15200
rect 10392 14112 10400 14176
rect 10464 14112 10480 14176
rect 10544 14112 10560 14176
rect 10624 14112 10640 14176
rect 10704 14112 10712 14176
rect 10392 13088 10712 14112
rect 10392 13024 10400 13088
rect 10464 13024 10480 13088
rect 10544 13024 10560 13088
rect 10624 13024 10640 13088
rect 10704 13024 10712 13088
rect 10392 12000 10712 13024
rect 10392 11936 10400 12000
rect 10464 11936 10480 12000
rect 10544 11936 10560 12000
rect 10624 11936 10640 12000
rect 10704 11936 10712 12000
rect 10392 10912 10712 11936
rect 10392 10848 10400 10912
rect 10464 10848 10480 10912
rect 10544 10848 10560 10912
rect 10624 10848 10640 10912
rect 10704 10848 10712 10912
rect 10392 9824 10712 10848
rect 10392 9760 10400 9824
rect 10464 9760 10480 9824
rect 10544 9760 10560 9824
rect 10624 9760 10640 9824
rect 10704 9760 10712 9824
rect 10392 8736 10712 9760
rect 10392 8672 10400 8736
rect 10464 8672 10480 8736
rect 10544 8672 10560 8736
rect 10624 8672 10640 8736
rect 10704 8672 10712 8736
rect 10392 7648 10712 8672
rect 10392 7584 10400 7648
rect 10464 7584 10480 7648
rect 10544 7584 10560 7648
rect 10624 7584 10640 7648
rect 10704 7584 10712 7648
rect 10392 6560 10712 7584
rect 10392 6496 10400 6560
rect 10464 6496 10480 6560
rect 10544 6496 10560 6560
rect 10624 6496 10640 6560
rect 10704 6496 10712 6560
rect 10392 5472 10712 6496
rect 10392 5408 10400 5472
rect 10464 5408 10480 5472
rect 10544 5408 10560 5472
rect 10624 5408 10640 5472
rect 10704 5408 10712 5472
rect 10392 4384 10712 5408
rect 10392 4320 10400 4384
rect 10464 4320 10480 4384
rect 10544 4320 10560 4384
rect 10624 4320 10640 4384
rect 10704 4320 10712 4384
rect 10392 3296 10712 4320
rect 10392 3232 10400 3296
rect 10464 3232 10480 3296
rect 10544 3232 10560 3296
rect 10624 3232 10640 3296
rect 10704 3232 10712 3296
rect 10392 2208 10712 3232
rect 10392 2144 10400 2208
rect 10464 2144 10480 2208
rect 10544 2144 10560 2208
rect 10624 2144 10640 2208
rect 10704 2144 10712 2208
rect 10392 2128 10712 2144
rect 15116 33216 15436 33776
rect 15116 33152 15124 33216
rect 15188 33152 15204 33216
rect 15268 33152 15284 33216
rect 15348 33152 15364 33216
rect 15428 33152 15436 33216
rect 15116 32128 15436 33152
rect 15116 32064 15124 32128
rect 15188 32064 15204 32128
rect 15268 32064 15284 32128
rect 15348 32064 15364 32128
rect 15428 32064 15436 32128
rect 15116 31040 15436 32064
rect 15116 30976 15124 31040
rect 15188 30976 15204 31040
rect 15268 30976 15284 31040
rect 15348 30976 15364 31040
rect 15428 30976 15436 31040
rect 15116 29952 15436 30976
rect 15116 29888 15124 29952
rect 15188 29888 15204 29952
rect 15268 29888 15284 29952
rect 15348 29888 15364 29952
rect 15428 29888 15436 29952
rect 15116 28864 15436 29888
rect 15116 28800 15124 28864
rect 15188 28800 15204 28864
rect 15268 28800 15284 28864
rect 15348 28800 15364 28864
rect 15428 28800 15436 28864
rect 15116 27776 15436 28800
rect 15116 27712 15124 27776
rect 15188 27712 15204 27776
rect 15268 27712 15284 27776
rect 15348 27712 15364 27776
rect 15428 27712 15436 27776
rect 15116 26688 15436 27712
rect 15116 26624 15124 26688
rect 15188 26624 15204 26688
rect 15268 26624 15284 26688
rect 15348 26624 15364 26688
rect 15428 26624 15436 26688
rect 15116 25600 15436 26624
rect 15116 25536 15124 25600
rect 15188 25536 15204 25600
rect 15268 25536 15284 25600
rect 15348 25536 15364 25600
rect 15428 25536 15436 25600
rect 15116 24512 15436 25536
rect 15116 24448 15124 24512
rect 15188 24448 15204 24512
rect 15268 24448 15284 24512
rect 15348 24448 15364 24512
rect 15428 24448 15436 24512
rect 15116 23424 15436 24448
rect 15116 23360 15124 23424
rect 15188 23360 15204 23424
rect 15268 23360 15284 23424
rect 15348 23360 15364 23424
rect 15428 23360 15436 23424
rect 15116 22336 15436 23360
rect 15116 22272 15124 22336
rect 15188 22272 15204 22336
rect 15268 22272 15284 22336
rect 15348 22272 15364 22336
rect 15428 22272 15436 22336
rect 15116 21248 15436 22272
rect 15116 21184 15124 21248
rect 15188 21184 15204 21248
rect 15268 21184 15284 21248
rect 15348 21184 15364 21248
rect 15428 21184 15436 21248
rect 15116 20160 15436 21184
rect 15116 20096 15124 20160
rect 15188 20096 15204 20160
rect 15268 20096 15284 20160
rect 15348 20096 15364 20160
rect 15428 20096 15436 20160
rect 15116 19072 15436 20096
rect 15116 19008 15124 19072
rect 15188 19008 15204 19072
rect 15268 19008 15284 19072
rect 15348 19008 15364 19072
rect 15428 19008 15436 19072
rect 15116 17984 15436 19008
rect 15116 17920 15124 17984
rect 15188 17920 15204 17984
rect 15268 17920 15284 17984
rect 15348 17920 15364 17984
rect 15428 17920 15436 17984
rect 15116 16896 15436 17920
rect 15116 16832 15124 16896
rect 15188 16832 15204 16896
rect 15268 16832 15284 16896
rect 15348 16832 15364 16896
rect 15428 16832 15436 16896
rect 15116 15808 15436 16832
rect 15116 15744 15124 15808
rect 15188 15744 15204 15808
rect 15268 15744 15284 15808
rect 15348 15744 15364 15808
rect 15428 15744 15436 15808
rect 15116 14720 15436 15744
rect 15116 14656 15124 14720
rect 15188 14656 15204 14720
rect 15268 14656 15284 14720
rect 15348 14656 15364 14720
rect 15428 14656 15436 14720
rect 15116 13632 15436 14656
rect 15116 13568 15124 13632
rect 15188 13568 15204 13632
rect 15268 13568 15284 13632
rect 15348 13568 15364 13632
rect 15428 13568 15436 13632
rect 15116 12544 15436 13568
rect 15116 12480 15124 12544
rect 15188 12480 15204 12544
rect 15268 12480 15284 12544
rect 15348 12480 15364 12544
rect 15428 12480 15436 12544
rect 15116 11456 15436 12480
rect 15116 11392 15124 11456
rect 15188 11392 15204 11456
rect 15268 11392 15284 11456
rect 15348 11392 15364 11456
rect 15428 11392 15436 11456
rect 15116 10368 15436 11392
rect 15116 10304 15124 10368
rect 15188 10304 15204 10368
rect 15268 10304 15284 10368
rect 15348 10304 15364 10368
rect 15428 10304 15436 10368
rect 15116 9280 15436 10304
rect 15116 9216 15124 9280
rect 15188 9216 15204 9280
rect 15268 9216 15284 9280
rect 15348 9216 15364 9280
rect 15428 9216 15436 9280
rect 15116 8192 15436 9216
rect 15116 8128 15124 8192
rect 15188 8128 15204 8192
rect 15268 8128 15284 8192
rect 15348 8128 15364 8192
rect 15428 8128 15436 8192
rect 15116 7104 15436 8128
rect 15116 7040 15124 7104
rect 15188 7040 15204 7104
rect 15268 7040 15284 7104
rect 15348 7040 15364 7104
rect 15428 7040 15436 7104
rect 15116 6016 15436 7040
rect 15116 5952 15124 6016
rect 15188 5952 15204 6016
rect 15268 5952 15284 6016
rect 15348 5952 15364 6016
rect 15428 5952 15436 6016
rect 15116 4928 15436 5952
rect 15116 4864 15124 4928
rect 15188 4864 15204 4928
rect 15268 4864 15284 4928
rect 15348 4864 15364 4928
rect 15428 4864 15436 4928
rect 15116 3840 15436 4864
rect 15116 3776 15124 3840
rect 15188 3776 15204 3840
rect 15268 3776 15284 3840
rect 15348 3776 15364 3840
rect 15428 3776 15436 3840
rect 15116 2752 15436 3776
rect 15116 2688 15124 2752
rect 15188 2688 15204 2752
rect 15268 2688 15284 2752
rect 15348 2688 15364 2752
rect 15428 2688 15436 2752
rect 15116 2128 15436 2688
rect 19840 33760 20160 33776
rect 19840 33696 19848 33760
rect 19912 33696 19928 33760
rect 19992 33696 20008 33760
rect 20072 33696 20088 33760
rect 20152 33696 20160 33760
rect 19840 32672 20160 33696
rect 19840 32608 19848 32672
rect 19912 32608 19928 32672
rect 19992 32608 20008 32672
rect 20072 32608 20088 32672
rect 20152 32608 20160 32672
rect 19840 31584 20160 32608
rect 19840 31520 19848 31584
rect 19912 31520 19928 31584
rect 19992 31520 20008 31584
rect 20072 31520 20088 31584
rect 20152 31520 20160 31584
rect 19840 30496 20160 31520
rect 19840 30432 19848 30496
rect 19912 30432 19928 30496
rect 19992 30432 20008 30496
rect 20072 30432 20088 30496
rect 20152 30432 20160 30496
rect 19840 29408 20160 30432
rect 19840 29344 19848 29408
rect 19912 29344 19928 29408
rect 19992 29344 20008 29408
rect 20072 29344 20088 29408
rect 20152 29344 20160 29408
rect 19840 28320 20160 29344
rect 19840 28256 19848 28320
rect 19912 28256 19928 28320
rect 19992 28256 20008 28320
rect 20072 28256 20088 28320
rect 20152 28256 20160 28320
rect 19840 27232 20160 28256
rect 19840 27168 19848 27232
rect 19912 27168 19928 27232
rect 19992 27168 20008 27232
rect 20072 27168 20088 27232
rect 20152 27168 20160 27232
rect 19840 26144 20160 27168
rect 19840 26080 19848 26144
rect 19912 26080 19928 26144
rect 19992 26080 20008 26144
rect 20072 26080 20088 26144
rect 20152 26080 20160 26144
rect 19840 25056 20160 26080
rect 19840 24992 19848 25056
rect 19912 24992 19928 25056
rect 19992 24992 20008 25056
rect 20072 24992 20088 25056
rect 20152 24992 20160 25056
rect 19840 23968 20160 24992
rect 19840 23904 19848 23968
rect 19912 23904 19928 23968
rect 19992 23904 20008 23968
rect 20072 23904 20088 23968
rect 20152 23904 20160 23968
rect 19840 22880 20160 23904
rect 19840 22816 19848 22880
rect 19912 22816 19928 22880
rect 19992 22816 20008 22880
rect 20072 22816 20088 22880
rect 20152 22816 20160 22880
rect 19840 21792 20160 22816
rect 19840 21728 19848 21792
rect 19912 21728 19928 21792
rect 19992 21728 20008 21792
rect 20072 21728 20088 21792
rect 20152 21728 20160 21792
rect 19840 20704 20160 21728
rect 19840 20640 19848 20704
rect 19912 20640 19928 20704
rect 19992 20640 20008 20704
rect 20072 20640 20088 20704
rect 20152 20640 20160 20704
rect 19840 19616 20160 20640
rect 19840 19552 19848 19616
rect 19912 19552 19928 19616
rect 19992 19552 20008 19616
rect 20072 19552 20088 19616
rect 20152 19552 20160 19616
rect 19840 18528 20160 19552
rect 19840 18464 19848 18528
rect 19912 18464 19928 18528
rect 19992 18464 20008 18528
rect 20072 18464 20088 18528
rect 20152 18464 20160 18528
rect 19840 17440 20160 18464
rect 19840 17376 19848 17440
rect 19912 17376 19928 17440
rect 19992 17376 20008 17440
rect 20072 17376 20088 17440
rect 20152 17376 20160 17440
rect 19840 16352 20160 17376
rect 19840 16288 19848 16352
rect 19912 16288 19928 16352
rect 19992 16288 20008 16352
rect 20072 16288 20088 16352
rect 20152 16288 20160 16352
rect 19840 15264 20160 16288
rect 19840 15200 19848 15264
rect 19912 15200 19928 15264
rect 19992 15200 20008 15264
rect 20072 15200 20088 15264
rect 20152 15200 20160 15264
rect 19840 14176 20160 15200
rect 19840 14112 19848 14176
rect 19912 14112 19928 14176
rect 19992 14112 20008 14176
rect 20072 14112 20088 14176
rect 20152 14112 20160 14176
rect 19840 13088 20160 14112
rect 19840 13024 19848 13088
rect 19912 13024 19928 13088
rect 19992 13024 20008 13088
rect 20072 13024 20088 13088
rect 20152 13024 20160 13088
rect 19840 12000 20160 13024
rect 19840 11936 19848 12000
rect 19912 11936 19928 12000
rect 19992 11936 20008 12000
rect 20072 11936 20088 12000
rect 20152 11936 20160 12000
rect 19840 10912 20160 11936
rect 19840 10848 19848 10912
rect 19912 10848 19928 10912
rect 19992 10848 20008 10912
rect 20072 10848 20088 10912
rect 20152 10848 20160 10912
rect 19840 9824 20160 10848
rect 19840 9760 19848 9824
rect 19912 9760 19928 9824
rect 19992 9760 20008 9824
rect 20072 9760 20088 9824
rect 20152 9760 20160 9824
rect 19840 8736 20160 9760
rect 19840 8672 19848 8736
rect 19912 8672 19928 8736
rect 19992 8672 20008 8736
rect 20072 8672 20088 8736
rect 20152 8672 20160 8736
rect 19840 7648 20160 8672
rect 19840 7584 19848 7648
rect 19912 7584 19928 7648
rect 19992 7584 20008 7648
rect 20072 7584 20088 7648
rect 20152 7584 20160 7648
rect 19840 6560 20160 7584
rect 19840 6496 19848 6560
rect 19912 6496 19928 6560
rect 19992 6496 20008 6560
rect 20072 6496 20088 6560
rect 20152 6496 20160 6560
rect 19840 5472 20160 6496
rect 19840 5408 19848 5472
rect 19912 5408 19928 5472
rect 19992 5408 20008 5472
rect 20072 5408 20088 5472
rect 20152 5408 20160 5472
rect 19840 4384 20160 5408
rect 19840 4320 19848 4384
rect 19912 4320 19928 4384
rect 19992 4320 20008 4384
rect 20072 4320 20088 4384
rect 20152 4320 20160 4384
rect 19840 3296 20160 4320
rect 19840 3232 19848 3296
rect 19912 3232 19928 3296
rect 19992 3232 20008 3296
rect 20072 3232 20088 3296
rect 20152 3232 20160 3296
rect 19840 2208 20160 3232
rect 19840 2144 19848 2208
rect 19912 2144 19928 2208
rect 19992 2144 20008 2208
rect 20072 2144 20088 2208
rect 20152 2144 20160 2208
rect 19840 2128 20160 2144
rect 24564 33216 24884 33776
rect 24564 33152 24572 33216
rect 24636 33152 24652 33216
rect 24716 33152 24732 33216
rect 24796 33152 24812 33216
rect 24876 33152 24884 33216
rect 24564 32128 24884 33152
rect 24564 32064 24572 32128
rect 24636 32064 24652 32128
rect 24716 32064 24732 32128
rect 24796 32064 24812 32128
rect 24876 32064 24884 32128
rect 24564 31040 24884 32064
rect 24564 30976 24572 31040
rect 24636 30976 24652 31040
rect 24716 30976 24732 31040
rect 24796 30976 24812 31040
rect 24876 30976 24884 31040
rect 24564 29952 24884 30976
rect 24564 29888 24572 29952
rect 24636 29888 24652 29952
rect 24716 29888 24732 29952
rect 24796 29888 24812 29952
rect 24876 29888 24884 29952
rect 24564 28864 24884 29888
rect 24564 28800 24572 28864
rect 24636 28800 24652 28864
rect 24716 28800 24732 28864
rect 24796 28800 24812 28864
rect 24876 28800 24884 28864
rect 24564 27776 24884 28800
rect 24564 27712 24572 27776
rect 24636 27712 24652 27776
rect 24716 27712 24732 27776
rect 24796 27712 24812 27776
rect 24876 27712 24884 27776
rect 24564 26688 24884 27712
rect 24564 26624 24572 26688
rect 24636 26624 24652 26688
rect 24716 26624 24732 26688
rect 24796 26624 24812 26688
rect 24876 26624 24884 26688
rect 24564 25600 24884 26624
rect 24564 25536 24572 25600
rect 24636 25536 24652 25600
rect 24716 25536 24732 25600
rect 24796 25536 24812 25600
rect 24876 25536 24884 25600
rect 24564 24512 24884 25536
rect 24564 24448 24572 24512
rect 24636 24448 24652 24512
rect 24716 24448 24732 24512
rect 24796 24448 24812 24512
rect 24876 24448 24884 24512
rect 24564 23424 24884 24448
rect 24564 23360 24572 23424
rect 24636 23360 24652 23424
rect 24716 23360 24732 23424
rect 24796 23360 24812 23424
rect 24876 23360 24884 23424
rect 24564 22336 24884 23360
rect 24564 22272 24572 22336
rect 24636 22272 24652 22336
rect 24716 22272 24732 22336
rect 24796 22272 24812 22336
rect 24876 22272 24884 22336
rect 24564 21248 24884 22272
rect 24564 21184 24572 21248
rect 24636 21184 24652 21248
rect 24716 21184 24732 21248
rect 24796 21184 24812 21248
rect 24876 21184 24884 21248
rect 24564 20160 24884 21184
rect 24564 20096 24572 20160
rect 24636 20096 24652 20160
rect 24716 20096 24732 20160
rect 24796 20096 24812 20160
rect 24876 20096 24884 20160
rect 24564 19072 24884 20096
rect 24564 19008 24572 19072
rect 24636 19008 24652 19072
rect 24716 19008 24732 19072
rect 24796 19008 24812 19072
rect 24876 19008 24884 19072
rect 24564 17984 24884 19008
rect 24564 17920 24572 17984
rect 24636 17920 24652 17984
rect 24716 17920 24732 17984
rect 24796 17920 24812 17984
rect 24876 17920 24884 17984
rect 24564 16896 24884 17920
rect 24564 16832 24572 16896
rect 24636 16832 24652 16896
rect 24716 16832 24732 16896
rect 24796 16832 24812 16896
rect 24876 16832 24884 16896
rect 24564 15808 24884 16832
rect 24564 15744 24572 15808
rect 24636 15744 24652 15808
rect 24716 15744 24732 15808
rect 24796 15744 24812 15808
rect 24876 15744 24884 15808
rect 24564 14720 24884 15744
rect 24564 14656 24572 14720
rect 24636 14656 24652 14720
rect 24716 14656 24732 14720
rect 24796 14656 24812 14720
rect 24876 14656 24884 14720
rect 24564 13632 24884 14656
rect 24564 13568 24572 13632
rect 24636 13568 24652 13632
rect 24716 13568 24732 13632
rect 24796 13568 24812 13632
rect 24876 13568 24884 13632
rect 24564 12544 24884 13568
rect 24564 12480 24572 12544
rect 24636 12480 24652 12544
rect 24716 12480 24732 12544
rect 24796 12480 24812 12544
rect 24876 12480 24884 12544
rect 24564 11456 24884 12480
rect 24564 11392 24572 11456
rect 24636 11392 24652 11456
rect 24716 11392 24732 11456
rect 24796 11392 24812 11456
rect 24876 11392 24884 11456
rect 24564 10368 24884 11392
rect 24564 10304 24572 10368
rect 24636 10304 24652 10368
rect 24716 10304 24732 10368
rect 24796 10304 24812 10368
rect 24876 10304 24884 10368
rect 24564 9280 24884 10304
rect 24564 9216 24572 9280
rect 24636 9216 24652 9280
rect 24716 9216 24732 9280
rect 24796 9216 24812 9280
rect 24876 9216 24884 9280
rect 24564 8192 24884 9216
rect 24564 8128 24572 8192
rect 24636 8128 24652 8192
rect 24716 8128 24732 8192
rect 24796 8128 24812 8192
rect 24876 8128 24884 8192
rect 24564 7104 24884 8128
rect 24564 7040 24572 7104
rect 24636 7040 24652 7104
rect 24716 7040 24732 7104
rect 24796 7040 24812 7104
rect 24876 7040 24884 7104
rect 24564 6016 24884 7040
rect 24564 5952 24572 6016
rect 24636 5952 24652 6016
rect 24716 5952 24732 6016
rect 24796 5952 24812 6016
rect 24876 5952 24884 6016
rect 24564 4928 24884 5952
rect 24564 4864 24572 4928
rect 24636 4864 24652 4928
rect 24716 4864 24732 4928
rect 24796 4864 24812 4928
rect 24876 4864 24884 4928
rect 24564 3840 24884 4864
rect 24564 3776 24572 3840
rect 24636 3776 24652 3840
rect 24716 3776 24732 3840
rect 24796 3776 24812 3840
rect 24876 3776 24884 3840
rect 24564 2752 24884 3776
rect 24564 2688 24572 2752
rect 24636 2688 24652 2752
rect 24716 2688 24732 2752
rect 24796 2688 24812 2752
rect 24876 2688 24884 2752
rect 24564 2128 24884 2688
rect 29288 33760 29608 33776
rect 29288 33696 29296 33760
rect 29360 33696 29376 33760
rect 29440 33696 29456 33760
rect 29520 33696 29536 33760
rect 29600 33696 29608 33760
rect 29288 32672 29608 33696
rect 29288 32608 29296 32672
rect 29360 32608 29376 32672
rect 29440 32608 29456 32672
rect 29520 32608 29536 32672
rect 29600 32608 29608 32672
rect 29288 31584 29608 32608
rect 29288 31520 29296 31584
rect 29360 31520 29376 31584
rect 29440 31520 29456 31584
rect 29520 31520 29536 31584
rect 29600 31520 29608 31584
rect 29288 30496 29608 31520
rect 29288 30432 29296 30496
rect 29360 30432 29376 30496
rect 29440 30432 29456 30496
rect 29520 30432 29536 30496
rect 29600 30432 29608 30496
rect 29288 29408 29608 30432
rect 29288 29344 29296 29408
rect 29360 29344 29376 29408
rect 29440 29344 29456 29408
rect 29520 29344 29536 29408
rect 29600 29344 29608 29408
rect 29288 28320 29608 29344
rect 29288 28256 29296 28320
rect 29360 28256 29376 28320
rect 29440 28256 29456 28320
rect 29520 28256 29536 28320
rect 29600 28256 29608 28320
rect 29288 27232 29608 28256
rect 29288 27168 29296 27232
rect 29360 27168 29376 27232
rect 29440 27168 29456 27232
rect 29520 27168 29536 27232
rect 29600 27168 29608 27232
rect 29288 26144 29608 27168
rect 29288 26080 29296 26144
rect 29360 26080 29376 26144
rect 29440 26080 29456 26144
rect 29520 26080 29536 26144
rect 29600 26080 29608 26144
rect 29288 25056 29608 26080
rect 29288 24992 29296 25056
rect 29360 24992 29376 25056
rect 29440 24992 29456 25056
rect 29520 24992 29536 25056
rect 29600 24992 29608 25056
rect 29288 23968 29608 24992
rect 29288 23904 29296 23968
rect 29360 23904 29376 23968
rect 29440 23904 29456 23968
rect 29520 23904 29536 23968
rect 29600 23904 29608 23968
rect 29288 22880 29608 23904
rect 29288 22816 29296 22880
rect 29360 22816 29376 22880
rect 29440 22816 29456 22880
rect 29520 22816 29536 22880
rect 29600 22816 29608 22880
rect 29288 21792 29608 22816
rect 29288 21728 29296 21792
rect 29360 21728 29376 21792
rect 29440 21728 29456 21792
rect 29520 21728 29536 21792
rect 29600 21728 29608 21792
rect 29288 20704 29608 21728
rect 29288 20640 29296 20704
rect 29360 20640 29376 20704
rect 29440 20640 29456 20704
rect 29520 20640 29536 20704
rect 29600 20640 29608 20704
rect 29288 19616 29608 20640
rect 29288 19552 29296 19616
rect 29360 19552 29376 19616
rect 29440 19552 29456 19616
rect 29520 19552 29536 19616
rect 29600 19552 29608 19616
rect 29288 18528 29608 19552
rect 29288 18464 29296 18528
rect 29360 18464 29376 18528
rect 29440 18464 29456 18528
rect 29520 18464 29536 18528
rect 29600 18464 29608 18528
rect 29288 17440 29608 18464
rect 29288 17376 29296 17440
rect 29360 17376 29376 17440
rect 29440 17376 29456 17440
rect 29520 17376 29536 17440
rect 29600 17376 29608 17440
rect 29288 16352 29608 17376
rect 29288 16288 29296 16352
rect 29360 16288 29376 16352
rect 29440 16288 29456 16352
rect 29520 16288 29536 16352
rect 29600 16288 29608 16352
rect 29288 15264 29608 16288
rect 29288 15200 29296 15264
rect 29360 15200 29376 15264
rect 29440 15200 29456 15264
rect 29520 15200 29536 15264
rect 29600 15200 29608 15264
rect 29288 14176 29608 15200
rect 29288 14112 29296 14176
rect 29360 14112 29376 14176
rect 29440 14112 29456 14176
rect 29520 14112 29536 14176
rect 29600 14112 29608 14176
rect 29288 13088 29608 14112
rect 29288 13024 29296 13088
rect 29360 13024 29376 13088
rect 29440 13024 29456 13088
rect 29520 13024 29536 13088
rect 29600 13024 29608 13088
rect 29288 12000 29608 13024
rect 29288 11936 29296 12000
rect 29360 11936 29376 12000
rect 29440 11936 29456 12000
rect 29520 11936 29536 12000
rect 29600 11936 29608 12000
rect 29288 10912 29608 11936
rect 29288 10848 29296 10912
rect 29360 10848 29376 10912
rect 29440 10848 29456 10912
rect 29520 10848 29536 10912
rect 29600 10848 29608 10912
rect 29288 9824 29608 10848
rect 29288 9760 29296 9824
rect 29360 9760 29376 9824
rect 29440 9760 29456 9824
rect 29520 9760 29536 9824
rect 29600 9760 29608 9824
rect 29288 8736 29608 9760
rect 29288 8672 29296 8736
rect 29360 8672 29376 8736
rect 29440 8672 29456 8736
rect 29520 8672 29536 8736
rect 29600 8672 29608 8736
rect 29288 7648 29608 8672
rect 29288 7584 29296 7648
rect 29360 7584 29376 7648
rect 29440 7584 29456 7648
rect 29520 7584 29536 7648
rect 29600 7584 29608 7648
rect 29288 6560 29608 7584
rect 29288 6496 29296 6560
rect 29360 6496 29376 6560
rect 29440 6496 29456 6560
rect 29520 6496 29536 6560
rect 29600 6496 29608 6560
rect 29288 5472 29608 6496
rect 29288 5408 29296 5472
rect 29360 5408 29376 5472
rect 29440 5408 29456 5472
rect 29520 5408 29536 5472
rect 29600 5408 29608 5472
rect 29288 4384 29608 5408
rect 29288 4320 29296 4384
rect 29360 4320 29376 4384
rect 29440 4320 29456 4384
rect 29520 4320 29536 4384
rect 29600 4320 29608 4384
rect 29288 3296 29608 4320
rect 29288 3232 29296 3296
rect 29360 3232 29376 3296
rect 29440 3232 29456 3296
rect 29520 3232 29536 3296
rect 29600 3232 29608 3296
rect 29288 2208 29608 3232
rect 29288 2144 29296 2208
rect 29360 2144 29376 2208
rect 29440 2144 29456 2208
rect 29520 2144 29536 2208
rect 29600 2144 29608 2208
rect 29288 2128 29608 2144
rect 34012 33216 34332 33776
rect 34012 33152 34020 33216
rect 34084 33152 34100 33216
rect 34164 33152 34180 33216
rect 34244 33152 34260 33216
rect 34324 33152 34332 33216
rect 34012 32128 34332 33152
rect 34012 32064 34020 32128
rect 34084 32064 34100 32128
rect 34164 32064 34180 32128
rect 34244 32064 34260 32128
rect 34324 32064 34332 32128
rect 34012 31040 34332 32064
rect 34012 30976 34020 31040
rect 34084 30976 34100 31040
rect 34164 30976 34180 31040
rect 34244 30976 34260 31040
rect 34324 30976 34332 31040
rect 34012 29952 34332 30976
rect 34012 29888 34020 29952
rect 34084 29888 34100 29952
rect 34164 29888 34180 29952
rect 34244 29888 34260 29952
rect 34324 29888 34332 29952
rect 34012 28864 34332 29888
rect 34012 28800 34020 28864
rect 34084 28800 34100 28864
rect 34164 28800 34180 28864
rect 34244 28800 34260 28864
rect 34324 28800 34332 28864
rect 34012 27776 34332 28800
rect 34012 27712 34020 27776
rect 34084 27712 34100 27776
rect 34164 27712 34180 27776
rect 34244 27712 34260 27776
rect 34324 27712 34332 27776
rect 34012 26688 34332 27712
rect 34012 26624 34020 26688
rect 34084 26624 34100 26688
rect 34164 26624 34180 26688
rect 34244 26624 34260 26688
rect 34324 26624 34332 26688
rect 34012 25600 34332 26624
rect 34012 25536 34020 25600
rect 34084 25536 34100 25600
rect 34164 25536 34180 25600
rect 34244 25536 34260 25600
rect 34324 25536 34332 25600
rect 34012 24512 34332 25536
rect 34012 24448 34020 24512
rect 34084 24448 34100 24512
rect 34164 24448 34180 24512
rect 34244 24448 34260 24512
rect 34324 24448 34332 24512
rect 34012 23424 34332 24448
rect 34012 23360 34020 23424
rect 34084 23360 34100 23424
rect 34164 23360 34180 23424
rect 34244 23360 34260 23424
rect 34324 23360 34332 23424
rect 34012 22336 34332 23360
rect 34012 22272 34020 22336
rect 34084 22272 34100 22336
rect 34164 22272 34180 22336
rect 34244 22272 34260 22336
rect 34324 22272 34332 22336
rect 34012 21248 34332 22272
rect 34012 21184 34020 21248
rect 34084 21184 34100 21248
rect 34164 21184 34180 21248
rect 34244 21184 34260 21248
rect 34324 21184 34332 21248
rect 34012 20160 34332 21184
rect 34012 20096 34020 20160
rect 34084 20096 34100 20160
rect 34164 20096 34180 20160
rect 34244 20096 34260 20160
rect 34324 20096 34332 20160
rect 34012 19072 34332 20096
rect 34012 19008 34020 19072
rect 34084 19008 34100 19072
rect 34164 19008 34180 19072
rect 34244 19008 34260 19072
rect 34324 19008 34332 19072
rect 34012 17984 34332 19008
rect 34012 17920 34020 17984
rect 34084 17920 34100 17984
rect 34164 17920 34180 17984
rect 34244 17920 34260 17984
rect 34324 17920 34332 17984
rect 34012 16896 34332 17920
rect 34012 16832 34020 16896
rect 34084 16832 34100 16896
rect 34164 16832 34180 16896
rect 34244 16832 34260 16896
rect 34324 16832 34332 16896
rect 34012 15808 34332 16832
rect 34012 15744 34020 15808
rect 34084 15744 34100 15808
rect 34164 15744 34180 15808
rect 34244 15744 34260 15808
rect 34324 15744 34332 15808
rect 34012 14720 34332 15744
rect 34012 14656 34020 14720
rect 34084 14656 34100 14720
rect 34164 14656 34180 14720
rect 34244 14656 34260 14720
rect 34324 14656 34332 14720
rect 34012 13632 34332 14656
rect 34012 13568 34020 13632
rect 34084 13568 34100 13632
rect 34164 13568 34180 13632
rect 34244 13568 34260 13632
rect 34324 13568 34332 13632
rect 34012 12544 34332 13568
rect 34012 12480 34020 12544
rect 34084 12480 34100 12544
rect 34164 12480 34180 12544
rect 34244 12480 34260 12544
rect 34324 12480 34332 12544
rect 34012 11456 34332 12480
rect 34012 11392 34020 11456
rect 34084 11392 34100 11456
rect 34164 11392 34180 11456
rect 34244 11392 34260 11456
rect 34324 11392 34332 11456
rect 34012 10368 34332 11392
rect 34012 10304 34020 10368
rect 34084 10304 34100 10368
rect 34164 10304 34180 10368
rect 34244 10304 34260 10368
rect 34324 10304 34332 10368
rect 34012 9280 34332 10304
rect 34012 9216 34020 9280
rect 34084 9216 34100 9280
rect 34164 9216 34180 9280
rect 34244 9216 34260 9280
rect 34324 9216 34332 9280
rect 34012 8192 34332 9216
rect 34012 8128 34020 8192
rect 34084 8128 34100 8192
rect 34164 8128 34180 8192
rect 34244 8128 34260 8192
rect 34324 8128 34332 8192
rect 34012 7104 34332 8128
rect 34012 7040 34020 7104
rect 34084 7040 34100 7104
rect 34164 7040 34180 7104
rect 34244 7040 34260 7104
rect 34324 7040 34332 7104
rect 34012 6016 34332 7040
rect 34012 5952 34020 6016
rect 34084 5952 34100 6016
rect 34164 5952 34180 6016
rect 34244 5952 34260 6016
rect 34324 5952 34332 6016
rect 34012 4928 34332 5952
rect 34012 4864 34020 4928
rect 34084 4864 34100 4928
rect 34164 4864 34180 4928
rect 34244 4864 34260 4928
rect 34324 4864 34332 4928
rect 34012 3840 34332 4864
rect 34012 3776 34020 3840
rect 34084 3776 34100 3840
rect 34164 3776 34180 3840
rect 34244 3776 34260 3840
rect 34324 3776 34332 3840
rect 34012 2752 34332 3776
rect 34012 2688 34020 2752
rect 34084 2688 34100 2752
rect 34164 2688 34180 2752
rect 34244 2688 34260 2752
rect 34324 2688 34332 2752
rect 34012 2128 34332 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__293__A dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2392 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__302__A
timestamp 1649977179
transform 1 0 11500 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__309__B
timestamp 1649977179
transform -1 0 15548 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__310__A1
timestamp 1649977179
transform 1 0 13524 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__310__C1
timestamp 1649977179
transform 1 0 12972 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__314__A4
timestamp 1649977179
transform 1 0 15180 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__314__B1
timestamp 1649977179
transform 1 0 13248 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__315__A3
timestamp 1649977179
transform 1 0 14812 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__320__A2
timestamp 1649977179
transform 1 0 17204 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__321__A3
timestamp 1649977179
transform 1 0 15088 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__321__C1
timestamp 1649977179
transform -1 0 13616 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__322__A2
timestamp 1649977179
transform 1 0 2852 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__322__B1
timestamp 1649977179
transform 1 0 4140 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__323__A2
timestamp 1649977179
transform -1 0 2944 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__337__A
timestamp 1649977179
transform 1 0 13432 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__345__B_N
timestamp 1649977179
transform 1 0 8832 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__346__C
timestamp 1649977179
transform -1 0 11500 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__370__A
timestamp 1649977179
transform 1 0 26312 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__383__A
timestamp 1649977179
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__384__A
timestamp 1649977179
transform 1 0 2760 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__386__A
timestamp 1649977179
transform -1 0 23092 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__388__C
timestamp 1649977179
transform 1 0 18860 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__389__A
timestamp 1649977179
transform -1 0 3496 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__397__A1
timestamp 1649977179
transform 1 0 14812 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__398__B1
timestamp 1649977179
transform 1 0 12880 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__402__A
timestamp 1649977179
transform 1 0 17848 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__403__A
timestamp 1649977179
transform 1 0 9752 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__406__A
timestamp 1649977179
transform 1 0 9752 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__411__A
timestamp 1649977179
transform -1 0 22172 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__412__A
timestamp 1649977179
transform 1 0 19504 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__417__A
timestamp 1649977179
transform 1 0 15364 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__420__A
timestamp 1649977179
transform 1 0 19320 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__424__A
timestamp 1649977179
transform 1 0 34500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__426__A
timestamp 1649977179
transform -1 0 19136 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__427__A
timestamp 1649977179
transform 1 0 4600 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__430__A
timestamp 1649977179
transform -1 0 4232 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__432__A
timestamp 1649977179
transform 1 0 20516 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__434__A
timestamp 1649977179
transform 1 0 20240 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__436__A
timestamp 1649977179
transform 1 0 7360 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__438__A
timestamp 1649977179
transform 1 0 28980 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__442__A
timestamp 1649977179
transform 1 0 34040 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__446__A
timestamp 1649977179
transform 1 0 23368 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__450__A
timestamp 1649977179
transform 1 0 24012 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__452__A
timestamp 1649977179
transform 1 0 3772 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__454__A
timestamp 1649977179
transform 1 0 30912 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__456__A
timestamp 1649977179
transform 1 0 32292 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__457__A
timestamp 1649977179
transform -1 0 21988 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__459__A
timestamp 1649977179
transform 1 0 4876 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__459__B
timestamp 1649977179
transform 1 0 4324 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__461__A
timestamp 1649977179
transform 1 0 17480 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__463__A
timestamp 1649977179
transform 1 0 34776 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__465__A
timestamp 1649977179
transform -1 0 31556 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__465__B
timestamp 1649977179
transform 1 0 30820 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__467__A
timestamp 1649977179
transform 1 0 25576 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__469__A
timestamp 1649977179
transform -1 0 34132 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__471__A
timestamp 1649977179
transform 1 0 13892 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__472__A
timestamp 1649977179
transform 1 0 3496 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__474__A
timestamp 1649977179
transform 1 0 3772 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__476__A
timestamp 1649977179
transform -1 0 3956 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__478__A
timestamp 1649977179
transform 1 0 32108 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__480__A
timestamp 1649977179
transform 1 0 15456 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__482__A
timestamp 1649977179
transform -1 0 3312 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__482__B
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__484__A
timestamp 1649977179
transform 1 0 14352 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__486__A
timestamp 1649977179
transform 1 0 30176 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__493__A
timestamp 1649977179
transform 1 0 31924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__493__B
timestamp 1649977179
transform -1 0 31924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__499__A
timestamp 1649977179
transform 1 0 13340 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__506__A
timestamp 1649977179
transform 1 0 30636 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__511__A
timestamp 1649977179
transform 1 0 7360 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__511__B
timestamp 1649977179
transform 1 0 6808 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__515__A
timestamp 1649977179
transform -1 0 31924 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__522__A
timestamp 1649977179
transform -1 0 30636 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__522__B
timestamp 1649977179
transform 1 0 30084 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__528__A
timestamp 1649977179
transform 1 0 15364 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__529__B
timestamp 1649977179
transform 1 0 12328 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__535__A
timestamp 1649977179
transform 1 0 31924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__539__A
timestamp 1649977179
transform -1 0 7452 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__539__B
timestamp 1649977179
transform -1 0 7636 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__543__A
timestamp 1649977179
transform 1 0 31556 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__544__A
timestamp 1649977179
transform -1 0 27508 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__546__A
timestamp 1649977179
transform 1 0 26956 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__548__A
timestamp 1649977179
transform 1 0 31648 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__550__A
timestamp 1649977179
transform 1 0 29900 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__550__B
timestamp 1649977179
transform 1 0 30452 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__552__A
timestamp 1649977179
transform -1 0 29716 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__554__A
timestamp 1649977179
transform -1 0 32660 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__556__A
timestamp 1649977179
transform 1 0 12788 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__556__B
timestamp 1649977179
transform 1 0 13340 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__558__A
timestamp 1649977179
transform 1 0 9936 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__560__A
timestamp 1649977179
transform 1 0 4600 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__562__A
timestamp 1649977179
transform 1 0 26312 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__564__A
timestamp 1649977179
transform 1 0 19412 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__564__B
timestamp 1649977179
transform 1 0 20424 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__566__A
timestamp 1649977179
transform 1 0 8740 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__566__B
timestamp 1649977179
transform 1 0 9292 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__568__A
timestamp 1649977179
transform 1 0 18216 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__577__B
timestamp 1649977179
transform 1 0 23276 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__581__A
timestamp 1649977179
transform 1 0 31464 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__583__A
timestamp 1649977179
transform 1 0 9844 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__589__A
timestamp 1649977179
transform 1 0 8280 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__590__A
timestamp 1649977179
transform -1 0 10856 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__601__CLK
timestamp 1649977179
transform -1 0 11776 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__603__CLK
timestamp 1649977179
transform -1 0 12328 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__604__CLK
timestamp 1649977179
transform 1 0 10856 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__612__CLK
timestamp 1649977179
transform -1 0 8648 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__693__A
timestamp 1649977179
transform 1 0 2484 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__695__A
timestamp 1649977179
transform 1 0 2852 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1649977179
transform -1 0 7912 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 28428 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 30452 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 31648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 32292 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 34040 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 34684 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 36432 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 37444 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 36800 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 38180 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 12880 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 13800 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 14904 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 16192 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 17664 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 18768 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 20056 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 21344 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 23276 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 23644 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 3312 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 9292 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output23_A
timestamp 1649977179
transform 1 0 25576 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output26_A
timestamp 1649977179
transform 1 0 2116 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output27_A
timestamp 1649977179
transform -1 0 2300 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output28_A
timestamp 1649977179
transform 1 0 2116 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output29_A
timestamp 1649977179
transform -1 0 2300 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output30_A
timestamp 1649977179
transform -1 0 1932 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output33_A
timestamp 1649977179
transform -1 0 2300 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output34_A
timestamp 1649977179
transform -1 0 2300 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output35_A
timestamp 1649977179
transform 1 0 2116 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output36_A
timestamp 1649977179
transform 1 0 2116 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output37_A
timestamp 1649977179
transform 1 0 2116 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output38_A
timestamp 1649977179
transform -1 0 2300 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output39_A
timestamp 1649977179
transform 1 0 2116 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output40_A
timestamp 1649977179
transform -1 0 2300 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output41_A
timestamp 1649977179
transform 1 0 10028 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output43_A
timestamp 1649977179
transform 1 0 2116 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output44_A
timestamp 1649977179
transform 1 0 4876 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output49_A
timestamp 1649977179
transform -1 0 2300 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output51_A
timestamp 1649977179
transform 1 0 2116 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output52_A
timestamp 1649977179
transform 1 0 2116 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output54_A
timestamp 1649977179
transform -1 0 2300 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output55_A
timestamp 1649977179
transform 1 0 2116 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_repeater67_A
timestamp 1649977179
transform 1 0 30360 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_repeater68_A
timestamp 1649977179
transform 1 0 19688 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_repeater69_A
timestamp 1649977179
transform -1 0 20332 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_repeater71_A
timestamp 1649977179
transform -1 0 28612 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_repeater72_A
timestamp 1649977179
transform -1 0 31188 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2484 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3036 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24
timestamp 1649977179
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32
timestamp 1649977179
transform 1 0 4048 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36
timestamp 1649977179
transform 1 0 4416 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41
timestamp 1649977179
transform 1 0 4876 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47
timestamp 1649977179
transform 1 0 5428 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1649977179
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7268 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75
timestamp 1649977179
transform 1 0 8004 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80
timestamp 1649977179
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_93
timestamp 1649977179
transform 1 0 9660 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1649977179
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_119
timestamp 1649977179
transform 1 0 12052 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_127
timestamp 1649977179
transform 1 0 12788 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_131
timestamp 1649977179
transform 1 0 13156 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1649977179
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_144
timestamp 1649977179
transform 1 0 14352 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_150
timestamp 1649977179
transform 1 0 14904 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_157
timestamp 1649977179
transform 1 0 15548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_161
timestamp 1649977179
transform 1 0 15916 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_164
timestamp 1649977179
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_172
timestamp 1649977179
transform 1 0 16928 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_183
timestamp 1649977179
transform 1 0 17940 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_189
timestamp 1649977179
transform 1 0 18492 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_192
timestamp 1649977179
transform 1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_200
timestamp 1649977179
transform 1 0 19504 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_209
timestamp 1649977179
transform 1 0 20332 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_217
timestamp 1649977179
transform 1 0 21068 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_220
timestamp 1649977179
transform 1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_228
timestamp 1649977179
transform 1 0 22080 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_235
timestamp 1649977179
transform 1 0 22724 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_241
timestamp 1649977179
transform 1 0 23276 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_248
timestamp 1649977179
transform 1 0 23920 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_253
timestamp 1649977179
transform 1 0 24380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_257
timestamp 1649977179
transform 1 0 24748 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_262
timestamp 1649977179
transform 1 0 25208 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_268
timestamp 1649977179
transform 1 0 25760 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_281 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 26956 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_288
timestamp 1649977179
transform 1 0 27600 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_296
timestamp 1649977179
transform 1 0 28336 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_300
timestamp 1649977179
transform 1 0 28704 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_309
timestamp 1649977179
transform 1 0 29532 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_313
timestamp 1649977179
transform 1 0 29900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_319
timestamp 1649977179
transform 1 0 30452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_326
timestamp 1649977179
transform 1 0 31096 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_332
timestamp 1649977179
transform 1 0 31648 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_340
timestamp 1649977179
transform 1 0 32384 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_348
timestamp 1649977179
transform 1 0 33120 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_352
timestamp 1649977179
transform 1 0 33488 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_358
timestamp 1649977179
transform 1 0 34040 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_368
timestamp 1649977179
transform 1 0 34960 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_374
timestamp 1649977179
transform 1 0 35512 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_378
timestamp 1649977179
transform 1 0 35880 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_384
timestamp 1649977179
transform 1 0 36432 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_396
timestamp 1649977179
transform 1 0 37536 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_403
timestamp 1649977179
transform 1 0 38180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_13
timestamp 1649977179
transform 1 0 2300 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_20
timestamp 1649977179
transform 1 0 2944 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_26
timestamp 1649977179
transform 1 0 3496 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_38
timestamp 1649977179
transform 1 0 4600 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_43
timestamp 1649977179
transform 1 0 5060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1649977179
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1649977179
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1649977179
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1649977179
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1649977179
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1649977179
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_125
timestamp 1649977179
transform 1 0 12604 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_128
timestamp 1649977179
transform 1 0 12880 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_138
timestamp 1649977179
transform 1 0 13800 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_147
timestamp 1649977179
transform 1 0 14628 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_159
timestamp 1649977179
transform 1 0 15732 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1649977179
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_169
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_177
timestamp 1649977179
transform 1 0 17388 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_180
timestamp 1649977179
transform 1 0 17664 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_192
timestamp 1649977179
transform 1 0 18768 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_206
timestamp 1649977179
transform 1 0 20056 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_218
timestamp 1649977179
transform 1 0 21160 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1649977179
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_237
timestamp 1649977179
transform 1 0 22908 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_256
timestamp 1649977179
transform 1 0 24656 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_268
timestamp 1649977179
transform 1 0 25760 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1649977179
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_293
timestamp 1649977179
transform 1 0 28060 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_297
timestamp 1649977179
transform 1 0 28428 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_309
timestamp 1649977179
transform 1 0 29532 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_321
timestamp 1649977179
transform 1 0 30636 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_327
timestamp 1649977179
transform 1 0 31188 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_332
timestamp 1649977179
transform 1 0 31648 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_339
timestamp 1649977179
transform 1 0 32292 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_351
timestamp 1649977179
transform 1 0 33396 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_365
timestamp 1649977179
transform 1 0 34684 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_377
timestamp 1649977179
transform 1 0 35788 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_385
timestamp 1649977179
transform 1 0 36524 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_388
timestamp 1649977179
transform 1 0 36800 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_395
timestamp 1649977179
transform 1 0 37444 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_399
timestamp 1649977179
transform 1 0 37812 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_403
timestamp 1649977179
transform 1 0 38180 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_7
timestamp 1649977179
transform 1 0 1748 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_15
timestamp 1649977179
transform 1 0 2484 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_20
timestamp 1649977179
transform 1 0 2944 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1649977179
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1649977179
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1649977179
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1649977179
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_97
timestamp 1649977179
transform 1 0 10028 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_101
timestamp 1649977179
transform 1 0 10396 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_114
timestamp 1649977179
transform 1 0 11592 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_124
timestamp 1649977179
transform 1 0 12512 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_130
timestamp 1649977179
transform 1 0 13064 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1649977179
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1649977179
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_165
timestamp 1649977179
transform 1 0 16284 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_172
timestamp 1649977179
transform 1 0 16928 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_184
timestamp 1649977179
transform 1 0 18032 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_209
timestamp 1649977179
transform 1 0 20332 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_217
timestamp 1649977179
transform 1 0 21068 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_224
timestamp 1649977179
transform 1 0 21712 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_236
timestamp 1649977179
transform 1 0 22816 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_242
timestamp 1649977179
transform 1 0 23368 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1649977179
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1649977179
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1649977179
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1649977179
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_277
timestamp 1649977179
transform 1 0 26588 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_293
timestamp 1649977179
transform 1 0 28060 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_299
timestamp 1649977179
transform 1 0 28612 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1649977179
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_309
timestamp 1649977179
transform 1 0 29532 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_317
timestamp 1649977179
transform 1 0 30268 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_334
timestamp 1649977179
transform 1 0 31832 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_344
timestamp 1649977179
transform 1 0 32752 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_356
timestamp 1649977179
transform 1 0 33856 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1649977179
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_377
timestamp 1649977179
transform 1 0 35788 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_385
timestamp 1649977179
transform 1 0 36524 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_392
timestamp 1649977179
transform 1 0 37168 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_400
timestamp 1649977179
transform 1 0 37904 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_403
timestamp 1649977179
transform 1 0 38180 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_11
timestamp 1649977179
transform 1 0 2116 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_18
timestamp 1649977179
transform 1 0 2760 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_34
timestamp 1649977179
transform 1 0 4232 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 1649977179
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_70
timestamp 1649977179
transform 1 0 7544 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_82
timestamp 1649977179
transform 1 0 8648 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_90
timestamp 1649977179
transform 1 0 9384 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_103
timestamp 1649977179
transform 1 0 10580 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1649977179
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1649977179
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_137
timestamp 1649977179
transform 1 0 13708 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_145
timestamp 1649977179
transform 1 0 14444 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_151
timestamp 1649977179
transform 1 0 14996 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_163
timestamp 1649977179
transform 1 0 16100 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1649977179
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_181
timestamp 1649977179
transform 1 0 17756 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_196
timestamp 1649977179
transform 1 0 19136 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_204
timestamp 1649977179
transform 1 0 19872 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_211
timestamp 1649977179
transform 1 0 20516 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1649977179
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1649977179
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_237
timestamp 1649977179
transform 1 0 22908 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_246
timestamp 1649977179
transform 1 0 23736 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_258
timestamp 1649977179
transform 1 0 24840 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_270
timestamp 1649977179
transform 1 0 25944 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_278
timestamp 1649977179
transform 1 0 26680 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_281
timestamp 1649977179
transform 1 0 26956 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_289
timestamp 1649977179
transform 1 0 27692 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_299
timestamp 1649977179
transform 1 0 28612 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_311
timestamp 1649977179
transform 1 0 29716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_323
timestamp 1649977179
transform 1 0 30820 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1649977179
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1649977179
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1649977179
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1649977179
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1649977179
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1649977179
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1649977179
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1649977179
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_405
timestamp 1649977179
transform 1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_7
timestamp 1649977179
transform 1 0 1748 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_15
timestamp 1649977179
transform 1 0 2484 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_20
timestamp 1649977179
transform 1 0 2944 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_41
timestamp 1649977179
transform 1 0 4876 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_49
timestamp 1649977179
transform 1 0 5612 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_55
timestamp 1649977179
transform 1 0 6164 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_67
timestamp 1649977179
transform 1 0 7268 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_73
timestamp 1649977179
transform 1 0 7820 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_81
timestamp 1649977179
transform 1 0 8556 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1649977179
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1649977179
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1649977179
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1649977179
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1649977179
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_153
timestamp 1649977179
transform 1 0 15180 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_160
timestamp 1649977179
transform 1 0 15824 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_172
timestamp 1649977179
transform 1 0 16928 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_184
timestamp 1649977179
transform 1 0 18032 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_197
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_201
timestamp 1649977179
transform 1 0 19596 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_210
timestamp 1649977179
transform 1 0 20424 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_222
timestamp 1649977179
transform 1 0 21528 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_230
timestamp 1649977179
transform 1 0 22264 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_240
timestamp 1649977179
transform 1 0 23184 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1649977179
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1649977179
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_277
timestamp 1649977179
transform 1 0 26588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_281
timestamp 1649977179
transform 1 0 26956 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_289
timestamp 1649977179
transform 1 0 27692 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_296
timestamp 1649977179
transform 1 0 28336 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1649977179
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1649977179
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1649977179
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1649977179
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1649977179
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1649977179
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1649977179
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1649977179
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1649977179
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_401
timestamp 1649977179
transform 1 0 37996 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1649977179
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1649977179
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1649977179
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1649977179
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1649977179
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1649977179
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1649977179
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1649977179
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1649977179
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1649977179
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1649977179
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1649977179
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1649977179
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1649977179
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1649977179
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1649977179
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_193
timestamp 1649977179
transform 1 0 18860 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_197
timestamp 1649977179
transform 1 0 19228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_202
timestamp 1649977179
transform 1 0 19688 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_213
timestamp 1649977179
transform 1 0 20700 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_221
timestamp 1649977179
transform 1 0 21436 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_225
timestamp 1649977179
transform 1 0 21804 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_234
timestamp 1649977179
transform 1 0 22632 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_246
timestamp 1649977179
transform 1 0 23736 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_258
timestamp 1649977179
transform 1 0 24840 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_270
timestamp 1649977179
transform 1 0 25944 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_278
timestamp 1649977179
transform 1 0 26680 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_284
timestamp 1649977179
transform 1 0 27232 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_296
timestamp 1649977179
transform 1 0 28336 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_308
timestamp 1649977179
transform 1 0 29440 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_320
timestamp 1649977179
transform 1 0 30544 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_332
timestamp 1649977179
transform 1 0 31648 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1649977179
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1649977179
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1649977179
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1649977179
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1649977179
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1649977179
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1649977179
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_405
timestamp 1649977179
transform 1 0 38364 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1649977179
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1649977179
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_53
timestamp 1649977179
transform 1 0 5980 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_58
timestamp 1649977179
transform 1 0 6440 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_70
timestamp 1649977179
transform 1 0 7544 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1649977179
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1649977179
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1649977179
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1649977179
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1649977179
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1649977179
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1649977179
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1649977179
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1649977179
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1649977179
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_197
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1649977179
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_221
timestamp 1649977179
transform 1 0 21436 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_233
timestamp 1649977179
transform 1 0 22540 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_243
timestamp 1649977179
transform 1 0 23460 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1649977179
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1649977179
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1649977179
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_277
timestamp 1649977179
transform 1 0 26588 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_297
timestamp 1649977179
transform 1 0 28428 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_305
timestamp 1649977179
transform 1 0 29164 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1649977179
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1649977179
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1649977179
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1649977179
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1649977179
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1649977179
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1649977179
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1649977179
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1649977179
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_401
timestamp 1649977179
transform 1 0 37996 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_7
timestamp 1649977179
transform 1 0 1748 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_13
timestamp 1649977179
transform 1 0 2300 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_31
timestamp 1649977179
transform 1 0 3956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_43
timestamp 1649977179
transform 1 0 5060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1649977179
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1649977179
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1649977179
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1649977179
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1649977179
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1649977179
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1649977179
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1649977179
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1649977179
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1649977179
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1649977179
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1649977179
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_197
timestamp 1649977179
transform 1 0 19228 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_209
timestamp 1649977179
transform 1 0 20332 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_221
timestamp 1649977179
transform 1 0 21436 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1649977179
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1649977179
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1649977179
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1649977179
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1649977179
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1649977179
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1649977179
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1649977179
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1649977179
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_317
timestamp 1649977179
transform 1 0 30268 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_325
timestamp 1649977179
transform 1 0 31004 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_331
timestamp 1649977179
transform 1 0 31556 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1649977179
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1649977179
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1649977179
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1649977179
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1649977179
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1649977179
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_405
timestamp 1649977179
transform 1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1649977179
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1649977179
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_53
timestamp 1649977179
transform 1 0 5980 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_64
timestamp 1649977179
transform 1 0 6992 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_76
timestamp 1649977179
transform 1 0 8096 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1649977179
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1649977179
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1649977179
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1649977179
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1649977179
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1649977179
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1649977179
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_177
timestamp 1649977179
transform 1 0 17388 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_184
timestamp 1649977179
transform 1 0 18032 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_191
timestamp 1649977179
transform 1 0 18676 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1649977179
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_207
timestamp 1649977179
transform 1 0 20148 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_219
timestamp 1649977179
transform 1 0 21252 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_231
timestamp 1649977179
transform 1 0 22356 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_243
timestamp 1649977179
transform 1 0 23460 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1649977179
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1649977179
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_265
timestamp 1649977179
transform 1 0 25484 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_280
timestamp 1649977179
transform 1 0 26864 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_292
timestamp 1649977179
transform 1 0 27968 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_304
timestamp 1649977179
transform 1 0 29072 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_309
timestamp 1649977179
transform 1 0 29532 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_317
timestamp 1649977179
transform 1 0 30268 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_321
timestamp 1649977179
transform 1 0 30636 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_332
timestamp 1649977179
transform 1 0 31648 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_339
timestamp 1649977179
transform 1 0 32292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_351
timestamp 1649977179
transform 1 0 33396 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1649977179
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_368
timestamp 1649977179
transform 1 0 34960 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_380
timestamp 1649977179
transform 1 0 36064 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_392
timestamp 1649977179
transform 1 0 37168 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_404
timestamp 1649977179
transform 1 0 38272 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_7
timestamp 1649977179
transform 1 0 1748 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_13
timestamp 1649977179
transform 1 0 2300 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_25
timestamp 1649977179
transform 1 0 3404 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_37
timestamp 1649977179
transform 1 0 4508 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_49
timestamp 1649977179
transform 1 0 5612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1649977179
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_61
timestamp 1649977179
transform 1 0 6716 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_64
timestamp 1649977179
transform 1 0 6992 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_70
timestamp 1649977179
transform 1 0 7544 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_82
timestamp 1649977179
transform 1 0 8648 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_94
timestamp 1649977179
transform 1 0 9752 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_98
timestamp 1649977179
transform 1 0 10120 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1649977179
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_116
timestamp 1649977179
transform 1 0 11776 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_122
timestamp 1649977179
transform 1 0 12328 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_146
timestamp 1649977179
transform 1 0 14536 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_158
timestamp 1649977179
transform 1 0 15640 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1649977179
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_169
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_177
timestamp 1649977179
transform 1 0 17388 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_187
timestamp 1649977179
transform 1 0 18308 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_199
timestamp 1649977179
transform 1 0 19412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_211
timestamp 1649977179
transform 1 0 20516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1649977179
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1649977179
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1649977179
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1649977179
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1649977179
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1649977179
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1649977179
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1649977179
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1649977179
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_305
timestamp 1649977179
transform 1 0 29164 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_313
timestamp 1649977179
transform 1 0 29900 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_317
timestamp 1649977179
transform 1 0 30268 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_326
timestamp 1649977179
transform 1 0 31096 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_334
timestamp 1649977179
transform 1 0 31832 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1649977179
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1649977179
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1649977179
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1649977179
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1649977179
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1649977179
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_405
timestamp 1649977179
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_15
timestamp 1649977179
transform 1 0 2484 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_24
timestamp 1649977179
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1649977179
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_53
timestamp 1649977179
transform 1 0 5980 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_60
timestamp 1649977179
transform 1 0 6624 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_68
timestamp 1649977179
transform 1 0 7360 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_71
timestamp 1649977179
transform 1 0 7636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1649977179
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_85
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_107
timestamp 1649977179
transform 1 0 10948 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_115
timestamp 1649977179
transform 1 0 11684 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_136
timestamp 1649977179
transform 1 0 13616 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_144
timestamp 1649977179
transform 1 0 14352 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_156
timestamp 1649977179
transform 1 0 15456 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_168
timestamp 1649977179
transform 1 0 16560 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_180
timestamp 1649977179
transform 1 0 17664 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_192
timestamp 1649977179
transform 1 0 18768 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1649977179
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1649977179
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_233
timestamp 1649977179
transform 1 0 22540 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_241
timestamp 1649977179
transform 1 0 23276 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_244
timestamp 1649977179
transform 1 0 23552 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1649977179
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1649977179
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1649977179
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_292
timestamp 1649977179
transform 1 0 27968 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_304
timestamp 1649977179
transform 1 0 29072 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_309
timestamp 1649977179
transform 1 0 29532 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_317
timestamp 1649977179
transform 1 0 30268 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_320
timestamp 1649977179
transform 1 0 30544 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_328
timestamp 1649977179
transform 1 0 31280 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_332
timestamp 1649977179
transform 1 0 31648 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_335
timestamp 1649977179
transform 1 0 31924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_347
timestamp 1649977179
transform 1 0 33028 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_10_358
timestamp 1649977179
transform 1 0 34040 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_368
timestamp 1649977179
transform 1 0 34960 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_388
timestamp 1649977179
transform 1 0 36800 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_400
timestamp 1649977179
transform 1 0 37904 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_406
timestamp 1649977179
transform 1 0 38456 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_15
timestamp 1649977179
transform 1 0 2484 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_24
timestamp 1649977179
transform 1 0 3312 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_31
timestamp 1649977179
transform 1 0 3956 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_37
timestamp 1649977179
transform 1 0 4508 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_43
timestamp 1649977179
transform 1 0 5060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1649977179
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_57
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_61
timestamp 1649977179
transform 1 0 6716 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_67
timestamp 1649977179
transform 1 0 7268 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_73
timestamp 1649977179
transform 1 0 7820 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_79
timestamp 1649977179
transform 1 0 8372 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_85
timestamp 1649977179
transform 1 0 8924 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_91
timestamp 1649977179
transform 1 0 9476 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_103
timestamp 1649977179
transform 1 0 10580 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1649977179
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_125
timestamp 1649977179
transform 1 0 12604 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_132
timestamp 1649977179
transform 1 0 13248 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_144
timestamp 1649977179
transform 1 0 14352 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_156
timestamp 1649977179
transform 1 0 15456 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_169
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_177
timestamp 1649977179
transform 1 0 17388 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_190
timestamp 1649977179
transform 1 0 18584 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_198
timestamp 1649977179
transform 1 0 19320 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_204
timestamp 1649977179
transform 1 0 19872 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_216
timestamp 1649977179
transform 1 0 20976 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_225
timestamp 1649977179
transform 1 0 21804 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_239
timestamp 1649977179
transform 1 0 23092 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_243
timestamp 1649977179
transform 1 0 23460 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1649977179
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1649977179
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1649977179
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1649977179
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_284
timestamp 1649977179
transform 1 0 27232 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_300
timestamp 1649977179
transform 1 0 28704 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_312
timestamp 1649977179
transform 1 0 29808 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_315
timestamp 1649977179
transform 1 0 30084 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_321
timestamp 1649977179
transform 1 0 30636 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_330
timestamp 1649977179
transform 1 0 31464 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_342
timestamp 1649977179
transform 1 0 32568 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_354
timestamp 1649977179
transform 1 0 33672 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_366
timestamp 1649977179
transform 1 0 34776 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_378
timestamp 1649977179
transform 1 0 35880 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_390
timestamp 1649977179
transform 1 0 36984 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1649977179
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_405
timestamp 1649977179
transform 1 0 38364 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_7
timestamp 1649977179
transform 1 0 1748 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_13
timestamp 1649977179
transform 1 0 2300 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_22
timestamp 1649977179
transform 1 0 3128 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_31
timestamp 1649977179
transform 1 0 3956 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_43
timestamp 1649977179
transform 1 0 5060 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_55
timestamp 1649977179
transform 1 0 6164 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_62
timestamp 1649977179
transform 1 0 6808 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_66
timestamp 1649977179
transform 1 0 7176 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_69
timestamp 1649977179
transform 1 0 7452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_81
timestamp 1649977179
transform 1 0 8556 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1649977179
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1649977179
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1649977179
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1649977179
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1649977179
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1649977179
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1649977179
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1649977179
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1649977179
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1649977179
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_209
timestamp 1649977179
transform 1 0 20332 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_213
timestamp 1649977179
transform 1 0 20700 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_218
timestamp 1649977179
transform 1 0 21160 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_228
timestamp 1649977179
transform 1 0 22080 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_237
timestamp 1649977179
transform 1 0 22908 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_243
timestamp 1649977179
transform 1 0 23460 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1649977179
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1649977179
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_265
timestamp 1649977179
transform 1 0 25484 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_273
timestamp 1649977179
transform 1 0 26220 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_287
timestamp 1649977179
transform 1 0 27508 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_299
timestamp 1649977179
transform 1 0 28612 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1649977179
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_309
timestamp 1649977179
transform 1 0 29532 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_317
timestamp 1649977179
transform 1 0 30268 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_323
timestamp 1649977179
transform 1 0 30820 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_331
timestamp 1649977179
transform 1 0 31556 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_337
timestamp 1649977179
transform 1 0 32108 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_349
timestamp 1649977179
transform 1 0 33212 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_361
timestamp 1649977179
transform 1 0 34316 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1649977179
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1649977179
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1649977179
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_401
timestamp 1649977179
transform 1 0 37996 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_15
timestamp 1649977179
transform 1 0 2484 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_21
timestamp 1649977179
transform 1 0 3036 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_24
timestamp 1649977179
transform 1 0 3312 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_36
timestamp 1649977179
transform 1 0 4416 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_48
timestamp 1649977179
transform 1 0 5520 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_67
timestamp 1649977179
transform 1 0 7268 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_79
timestamp 1649977179
transform 1 0 8372 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_91
timestamp 1649977179
transform 1 0 9476 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_103
timestamp 1649977179
transform 1 0 10580 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1649977179
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1649977179
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1649977179
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1649977179
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1649977179
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1649977179
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1649977179
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1649977179
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1649977179
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1649977179
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1649977179
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_238
timestamp 1649977179
transform 1 0 23000 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_250
timestamp 1649977179
transform 1 0 24104 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_256
timestamp 1649977179
transform 1 0 24656 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_268
timestamp 1649977179
transform 1 0 25760 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1649977179
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1649977179
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1649977179
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_317
timestamp 1649977179
transform 1 0 30268 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_327
timestamp 1649977179
transform 1 0 31188 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1649977179
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1649977179
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1649977179
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1649977179
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1649977179
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1649977179
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1649977179
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1649977179
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_405
timestamp 1649977179
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_7
timestamp 1649977179
transform 1 0 1748 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_13
timestamp 1649977179
transform 1 0 2300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_25
timestamp 1649977179
transform 1 0 3404 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_37
timestamp 1649977179
transform 1 0 4508 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_42
timestamp 1649977179
transform 1 0 4968 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_54
timestamp 1649977179
transform 1 0 6072 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_66
timestamp 1649977179
transform 1 0 7176 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_78
timestamp 1649977179
transform 1 0 8280 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1649977179
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1649977179
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1649977179
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1649977179
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1649977179
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_153
timestamp 1649977179
transform 1 0 15180 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_161
timestamp 1649977179
transform 1 0 15916 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_172
timestamp 1649977179
transform 1 0 16928 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_184
timestamp 1649977179
transform 1 0 18032 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1649977179
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1649977179
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1649977179
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1649977179
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1649977179
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1649977179
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1649977179
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_277
timestamp 1649977179
transform 1 0 26588 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_283
timestamp 1649977179
transform 1 0 27140 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_287
timestamp 1649977179
transform 1 0 27508 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_299
timestamp 1649977179
transform 1 0 28612 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1649977179
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1649977179
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1649977179
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1649977179
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1649977179
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1649977179
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1649977179
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_365
timestamp 1649977179
transform 1 0 34684 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_373
timestamp 1649977179
transform 1 0 35420 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_386
timestamp 1649977179
transform 1 0 36616 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_398
timestamp 1649977179
transform 1 0 37720 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_406
timestamp 1649977179
transform 1 0 38456 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1649977179
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1649977179
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1649977179
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1649977179
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_57
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_68
timestamp 1649977179
transform 1 0 7360 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_80
timestamp 1649977179
transform 1 0 8464 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_92
timestamp 1649977179
transform 1 0 9568 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_104
timestamp 1649977179
transform 1 0 10672 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1649977179
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1649977179
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1649977179
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1649977179
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1649977179
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_181
timestamp 1649977179
transform 1 0 17756 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_189
timestamp 1649977179
transform 1 0 18492 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_195
timestamp 1649977179
transform 1 0 19044 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_207
timestamp 1649977179
transform 1 0 20148 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_219
timestamp 1649977179
transform 1 0 21252 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1649977179
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_225
timestamp 1649977179
transform 1 0 21804 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_233
timestamp 1649977179
transform 1 0 22540 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_239
timestamp 1649977179
transform 1 0 23092 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_251
timestamp 1649977179
transform 1 0 24196 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_263
timestamp 1649977179
transform 1 0 25300 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_275
timestamp 1649977179
transform 1 0 26404 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1649977179
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1649977179
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1649977179
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1649977179
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1649977179
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1649977179
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1649977179
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_339
timestamp 1649977179
transform 1 0 32292 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_350
timestamp 1649977179
transform 1 0 33304 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_357
timestamp 1649977179
transform 1 0 33948 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_365
timestamp 1649977179
transform 1 0 34684 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_378
timestamp 1649977179
transform 1 0 35880 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_390
timestamp 1649977179
transform 1 0 36984 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1649977179
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_405
timestamp 1649977179
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1649977179
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1649977179
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1649977179
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1649977179
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1649977179
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1649977179
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1649977179
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_85
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_93
timestamp 1649977179
transform 1 0 9660 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_99
timestamp 1649977179
transform 1 0 10212 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_111
timestamp 1649977179
transform 1 0 11316 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_123
timestamp 1649977179
transform 1 0 12420 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_131
timestamp 1649977179
transform 1 0 13156 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_136
timestamp 1649977179
transform 1 0 13616 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_149
timestamp 1649977179
transform 1 0 14812 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_161
timestamp 1649977179
transform 1 0 15916 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_171
timestamp 1649977179
transform 1 0 16836 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1649977179
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1649977179
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1649977179
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1649977179
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1649977179
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1649977179
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1649977179
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1649977179
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_258
timestamp 1649977179
transform 1 0 24840 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_270
timestamp 1649977179
transform 1 0 25944 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_278
timestamp 1649977179
transform 1 0 26680 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_282
timestamp 1649977179
transform 1 0 27048 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_294
timestamp 1649977179
transform 1 0 28152 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_306
timestamp 1649977179
transform 1 0 29256 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1649977179
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_321
timestamp 1649977179
transform 1 0 30636 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_326
timestamp 1649977179
transform 1 0 31096 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_335
timestamp 1649977179
transform 1 0 31924 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_344
timestamp 1649977179
transform 1 0 32752 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_356
timestamp 1649977179
transform 1 0 33856 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1649977179
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1649977179
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1649977179
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_401
timestamp 1649977179
transform 1 0 37996 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_7
timestamp 1649977179
transform 1 0 1748 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_13
timestamp 1649977179
transform 1 0 2300 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_17
timestamp 1649977179
transform 1 0 2668 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_20
timestamp 1649977179
transform 1 0 2944 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_30
timestamp 1649977179
transform 1 0 3864 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_42
timestamp 1649977179
transform 1 0 4968 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1649977179
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_60
timestamp 1649977179
transform 1 0 6624 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_72
timestamp 1649977179
transform 1 0 7728 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_82
timestamp 1649977179
transform 1 0 8648 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_106
timestamp 1649977179
transform 1 0 10856 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_125
timestamp 1649977179
transform 1 0 12604 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_132
timestamp 1649977179
transform 1 0 13248 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_140
timestamp 1649977179
transform 1 0 13984 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_148
timestamp 1649977179
transform 1 0 14720 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_154
timestamp 1649977179
transform 1 0 15272 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1649977179
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_181
timestamp 1649977179
transform 1 0 17756 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_187
timestamp 1649977179
transform 1 0 18308 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_199
timestamp 1649977179
transform 1 0 19412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_211
timestamp 1649977179
transform 1 0 20516 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1649977179
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1649977179
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1649977179
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1649977179
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1649977179
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1649977179
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1649977179
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_293
timestamp 1649977179
transform 1 0 28060 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_309
timestamp 1649977179
transform 1 0 29532 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_321
timestamp 1649977179
transform 1 0 30636 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_333
timestamp 1649977179
transform 1 0 31740 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1649977179
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1649977179
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1649977179
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1649977179
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1649977179
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1649977179
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1649977179
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_405
timestamp 1649977179
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_11
timestamp 1649977179
transform 1 0 2116 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_16
timestamp 1649977179
transform 1 0 2576 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_24
timestamp 1649977179
transform 1 0 3312 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_50
timestamp 1649977179
transform 1 0 5704 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_62
timestamp 1649977179
transform 1 0 6808 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_74
timestamp 1649977179
transform 1 0 7912 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1649977179
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_91
timestamp 1649977179
transform 1 0 9476 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1649977179
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1649977179
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_121
timestamp 1649977179
transform 1 0 12236 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_125
timestamp 1649977179
transform 1 0 12604 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_136
timestamp 1649977179
transform 1 0 13616 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_149
timestamp 1649977179
transform 1 0 14812 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_155
timestamp 1649977179
transform 1 0 15364 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_167
timestamp 1649977179
transform 1 0 16468 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_179
timestamp 1649977179
transform 1 0 17572 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_191
timestamp 1649977179
transform 1 0 18676 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1649977179
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1649977179
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1649977179
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1649977179
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1649977179
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1649977179
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_253
timestamp 1649977179
transform 1 0 24380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_259
timestamp 1649977179
transform 1 0 24932 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_263
timestamp 1649977179
transform 1 0 25300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_275
timestamp 1649977179
transform 1 0 26404 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_286
timestamp 1649977179
transform 1 0 27416 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_298
timestamp 1649977179
transform 1 0 28520 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_306
timestamp 1649977179
transform 1 0 29256 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1649977179
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1649977179
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_333
timestamp 1649977179
transform 1 0 31740 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_337
timestamp 1649977179
transform 1 0 32108 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_349
timestamp 1649977179
transform 1 0 33212 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_361
timestamp 1649977179
transform 1 0 34316 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1649977179
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1649977179
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_401
timestamp 1649977179
transform 1 0 37996 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_7
timestamp 1649977179
transform 1 0 1748 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_13
timestamp 1649977179
transform 1 0 2300 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_21
timestamp 1649977179
transform 1 0 3036 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_29
timestamp 1649977179
transform 1 0 3772 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_35
timestamp 1649977179
transform 1 0 4324 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_47
timestamp 1649977179
transform 1 0 5428 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1649977179
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1649977179
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1649977179
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1649977179
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1649977179
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1649977179
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_125
timestamp 1649977179
transform 1 0 12604 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_131
timestamp 1649977179
transform 1 0 13156 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_134
timestamp 1649977179
transform 1 0 13432 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_145
timestamp 1649977179
transform 1 0 14444 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_151
timestamp 1649977179
transform 1 0 14996 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_163
timestamp 1649977179
transform 1 0 16100 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1649977179
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_181
timestamp 1649977179
transform 1 0 17756 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_184
timestamp 1649977179
transform 1 0 18032 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_192
timestamp 1649977179
transform 1 0 18768 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_199
timestamp 1649977179
transform 1 0 19412 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_209
timestamp 1649977179
transform 1 0 20332 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_221
timestamp 1649977179
transform 1 0 21436 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_228
timestamp 1649977179
transform 1 0 22080 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_240
timestamp 1649977179
transform 1 0 23184 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1649977179
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1649977179
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_273
timestamp 1649977179
transform 1 0 26220 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_276
timestamp 1649977179
transform 1 0 26496 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_286
timestamp 1649977179
transform 1 0 27416 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_298
timestamp 1649977179
transform 1 0 28520 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_310
timestamp 1649977179
transform 1 0 29624 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_318
timestamp 1649977179
transform 1 0 30360 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_323
timestamp 1649977179
transform 1 0 30820 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_332
timestamp 1649977179
transform 1 0 31648 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_342
timestamp 1649977179
transform 1 0 32568 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_353
timestamp 1649977179
transform 1 0 33580 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_361
timestamp 1649977179
transform 1 0 34316 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_367
timestamp 1649977179
transform 1 0 34868 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_371
timestamp 1649977179
transform 1 0 35236 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_384
timestamp 1649977179
transform 1 0 36432 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1649977179
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_405
timestamp 1649977179
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1649977179
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1649977179
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1649977179
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_53
timestamp 1649977179
transform 1 0 5980 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_60
timestamp 1649977179
transform 1 0 6624 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_69
timestamp 1649977179
transform 1 0 7452 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_76
timestamp 1649977179
transform 1 0 8096 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_90
timestamp 1649977179
transform 1 0 9384 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_102
timestamp 1649977179
transform 1 0 10488 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_110
timestamp 1649977179
transform 1 0 11224 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_115
timestamp 1649977179
transform 1 0 11684 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_123
timestamp 1649977179
transform 1 0 12420 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_135
timestamp 1649977179
transform 1 0 13524 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1649977179
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1649977179
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_165
timestamp 1649977179
transform 1 0 16284 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_174
timestamp 1649977179
transform 1 0 17112 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_188
timestamp 1649977179
transform 1 0 18400 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_207
timestamp 1649977179
transform 1 0 20148 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_20_220
timestamp 1649977179
transform 1 0 21344 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_226
timestamp 1649977179
transform 1 0 21896 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_235
timestamp 1649977179
transform 1 0 22724 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_247
timestamp 1649977179
transform 1 0 23828 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1649977179
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_253
timestamp 1649977179
transform 1 0 24380 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_261
timestamp 1649977179
transform 1 0 25116 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_273
timestamp 1649977179
transform 1 0 26220 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_285
timestamp 1649977179
transform 1 0 27324 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_297
timestamp 1649977179
transform 1 0 28428 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_305
timestamp 1649977179
transform 1 0 29164 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1649977179
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1649977179
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1649977179
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1649977179
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1649977179
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1649977179
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1649977179
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1649977179
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1649977179
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_401
timestamp 1649977179
transform 1 0 37996 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1649977179
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1649977179
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1649977179
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1649977179
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1649977179
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_69
timestamp 1649977179
transform 1 0 7452 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_74
timestamp 1649977179
transform 1 0 7912 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_80
timestamp 1649977179
transform 1 0 8464 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_92
timestamp 1649977179
transform 1 0 9568 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_104
timestamp 1649977179
transform 1 0 10672 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1649977179
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1649977179
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1649977179
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1649977179
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1649977179
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_169
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_177
timestamp 1649977179
transform 1 0 17388 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_189
timestamp 1649977179
transform 1 0 18492 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_201
timestamp 1649977179
transform 1 0 19596 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_213
timestamp 1649977179
transform 1 0 20700 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_221
timestamp 1649977179
transform 1 0 21436 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_233
timestamp 1649977179
transform 1 0 22540 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_244
timestamp 1649977179
transform 1 0 23552 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_256
timestamp 1649977179
transform 1 0 24656 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_268
timestamp 1649977179
transform 1 0 25760 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_276
timestamp 1649977179
transform 1 0 26496 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_287
timestamp 1649977179
transform 1 0 27508 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_299
timestamp 1649977179
transform 1 0 28612 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_311
timestamp 1649977179
transform 1 0 29716 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_323
timestamp 1649977179
transform 1 0 30820 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_329
timestamp 1649977179
transform 1 0 31372 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_332
timestamp 1649977179
transform 1 0 31648 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_342
timestamp 1649977179
transform 1 0 32568 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_354
timestamp 1649977179
transform 1 0 33672 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_366
timestamp 1649977179
transform 1 0 34776 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_378
timestamp 1649977179
transform 1 0 35880 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_390
timestamp 1649977179
transform 1 0 36984 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1649977179
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_405
timestamp 1649977179
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_7
timestamp 1649977179
transform 1 0 1748 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_13
timestamp 1649977179
transform 1 0 2300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_25
timestamp 1649977179
transform 1 0 3404 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_41
timestamp 1649977179
transform 1 0 4876 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_67
timestamp 1649977179
transform 1 0 7268 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_79
timestamp 1649977179
transform 1 0 8372 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1649977179
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_103
timestamp 1649977179
transform 1 0 10580 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_115
timestamp 1649977179
transform 1 0 11684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_127
timestamp 1649977179
transform 1 0 12788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1649977179
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_163
timestamp 1649977179
transform 1 0 16100 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_177
timestamp 1649977179
transform 1 0 17388 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_181
timestamp 1649977179
transform 1 0 17756 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_192
timestamp 1649977179
transform 1 0 18768 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1649977179
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_221
timestamp 1649977179
transform 1 0 21436 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1649977179
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1649977179
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1649977179
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1649977179
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1649977179
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_277
timestamp 1649977179
transform 1 0 26588 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_282
timestamp 1649977179
transform 1 0 27048 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_294
timestamp 1649977179
transform 1 0 28152 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_306
timestamp 1649977179
transform 1 0 29256 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1649977179
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_321
timestamp 1649977179
transform 1 0 30636 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_325
timestamp 1649977179
transform 1 0 31004 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_331
timestamp 1649977179
transform 1 0 31556 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_338
timestamp 1649977179
transform 1 0 32200 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_350
timestamp 1649977179
transform 1 0 33304 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_355
timestamp 1649977179
transform 1 0 33764 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1649977179
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1649977179
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1649977179
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1649977179
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_401
timestamp 1649977179
transform 1 0 37996 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1649977179
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1649977179
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1649977179
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1649977179
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1649977179
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1649977179
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_81
timestamp 1649977179
transform 1 0 8556 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_86
timestamp 1649977179
transform 1 0 9016 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_108
timestamp 1649977179
transform 1 0 11040 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1649977179
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1649977179
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_149
timestamp 1649977179
transform 1 0 14812 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_163
timestamp 1649977179
transform 1 0 16100 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1649977179
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_169
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_177
timestamp 1649977179
transform 1 0 17388 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_188
timestamp 1649977179
transform 1 0 18400 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_195
timestamp 1649977179
transform 1 0 19044 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_207
timestamp 1649977179
transform 1 0 20148 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_219
timestamp 1649977179
transform 1 0 21252 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1649977179
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1649977179
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1649977179
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_249
timestamp 1649977179
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_261
timestamp 1649977179
transform 1 0 25116 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_267
timestamp 1649977179
transform 1 0 25668 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_274
timestamp 1649977179
transform 1 0 26312 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_291
timestamp 1649977179
transform 1 0 27876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_303
timestamp 1649977179
transform 1 0 28980 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_311
timestamp 1649977179
transform 1 0 29716 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1649977179
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1649977179
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1649977179
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_337
timestamp 1649977179
transform 1 0 32108 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_23_348
timestamp 1649977179
transform 1 0 33120 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_360
timestamp 1649977179
transform 1 0 34224 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_375
timestamp 1649977179
transform 1 0 35604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_387
timestamp 1649977179
transform 1 0 36708 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1649977179
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1649977179
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_405
timestamp 1649977179
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_7
timestamp 1649977179
transform 1 0 1748 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_13
timestamp 1649977179
transform 1 0 2300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_25
timestamp 1649977179
transform 1 0 3404 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1649977179
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1649977179
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1649977179
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1649977179
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1649977179
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_96
timestamp 1649977179
transform 1 0 9936 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_108
timestamp 1649977179
transform 1 0 11040 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_116
timestamp 1649977179
transform 1 0 11776 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_128
timestamp 1649977179
transform 1 0 12880 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1649977179
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1649977179
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1649977179
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1649977179
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1649977179
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1649977179
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1649977179
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1649977179
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1649977179
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1649977179
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_253
timestamp 1649977179
transform 1 0 24380 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_259
timestamp 1649977179
transform 1 0 24932 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_271
timestamp 1649977179
transform 1 0 26036 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_283
timestamp 1649977179
transform 1 0 27140 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_295
timestamp 1649977179
transform 1 0 28244 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1649977179
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_309
timestamp 1649977179
transform 1 0 29532 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_323
timestamp 1649977179
transform 1 0 30820 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_335
timestamp 1649977179
transform 1 0 31924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_347
timestamp 1649977179
transform 1 0 33028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_359
timestamp 1649977179
transform 1 0 34132 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1649977179
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1649977179
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_377
timestamp 1649977179
transform 1 0 35788 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_383
timestamp 1649977179
transform 1 0 36340 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_396
timestamp 1649977179
transform 1 0 37536 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_404
timestamp 1649977179
transform 1 0 38272 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_15
timestamp 1649977179
transform 1 0 2484 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_21
timestamp 1649977179
transform 1 0 3036 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_33
timestamp 1649977179
transform 1 0 4140 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_45
timestamp 1649977179
transform 1 0 5244 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 1649977179
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_69
timestamp 1649977179
transform 1 0 7452 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_93
timestamp 1649977179
transform 1 0 9660 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_103
timestamp 1649977179
transform 1 0 10580 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1649977179
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_123
timestamp 1649977179
transform 1 0 12420 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_135
timestamp 1649977179
transform 1 0 13524 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_147
timestamp 1649977179
transform 1 0 14628 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_159
timestamp 1649977179
transform 1 0 15732 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1649977179
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1649977179
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_193
timestamp 1649977179
transform 1 0 18860 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_25_204
timestamp 1649977179
transform 1 0 19872 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_216
timestamp 1649977179
transform 1 0 20976 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1649977179
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1649977179
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1649977179
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_261
timestamp 1649977179
transform 1 0 25116 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_276
timestamp 1649977179
transform 1 0 26496 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1649977179
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_293
timestamp 1649977179
transform 1 0 28060 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_301
timestamp 1649977179
transform 1 0 28796 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_305
timestamp 1649977179
transform 1 0 29164 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_314
timestamp 1649977179
transform 1 0 29992 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_326
timestamp 1649977179
transform 1 0 31096 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_334
timestamp 1649977179
transform 1 0 31832 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1649977179
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1649977179
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_361
timestamp 1649977179
transform 1 0 34316 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_365
timestamp 1649977179
transform 1 0 34684 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_373
timestamp 1649977179
transform 1 0 35420 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_379
timestamp 1649977179
transform 1 0 35972 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1649977179
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1649977179
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_405
timestamp 1649977179
transform 1 0 38364 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_11
timestamp 1649977179
transform 1 0 2116 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_24
timestamp 1649977179
transform 1 0 3312 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_34
timestamp 1649977179
transform 1 0 4232 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_40
timestamp 1649977179
transform 1 0 4784 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_52
timestamp 1649977179
transform 1 0 5888 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_59
timestamp 1649977179
transform 1 0 6532 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_67
timestamp 1649977179
transform 1 0 7268 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_79
timestamp 1649977179
transform 1 0 8372 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1649977179
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_85
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_98
timestamp 1649977179
transform 1 0 10120 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_110
timestamp 1649977179
transform 1 0 11224 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_113
timestamp 1649977179
transform 1 0 11500 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_123
timestamp 1649977179
transform 1 0 12420 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_135
timestamp 1649977179
transform 1 0 13524 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1649977179
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_153
timestamp 1649977179
transform 1 0 15180 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_159
timestamp 1649977179
transform 1 0 15732 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_166
timestamp 1649977179
transform 1 0 16376 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_178
timestamp 1649977179
transform 1 0 17480 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_190
timestamp 1649977179
transform 1 0 18584 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_26_197
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_213
timestamp 1649977179
transform 1 0 20700 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_224
timestamp 1649977179
transform 1 0 21712 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_232
timestamp 1649977179
transform 1 0 22448 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_239
timestamp 1649977179
transform 1 0 23092 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1649977179
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1649977179
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1649977179
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1649977179
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_289
timestamp 1649977179
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1649977179
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1649977179
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1649977179
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1649977179
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_333
timestamp 1649977179
transform 1 0 31740 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_344
timestamp 1649977179
transform 1 0 32752 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_356
timestamp 1649977179
transform 1 0 33856 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_360
timestamp 1649977179
transform 1 0 34224 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_370
timestamp 1649977179
transform 1 0 35144 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_388
timestamp 1649977179
transform 1 0 36800 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_400
timestamp 1649977179
transform 1 0 37904 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_406
timestamp 1649977179
transform 1 0 38456 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_7
timestamp 1649977179
transform 1 0 1748 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_13
timestamp 1649977179
transform 1 0 2300 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_25
timestamp 1649977179
transform 1 0 3404 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_37
timestamp 1649977179
transform 1 0 4508 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_49
timestamp 1649977179
transform 1 0 5612 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1649977179
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1649977179
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1649977179
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1649977179
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1649977179
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1649977179
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1649977179
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1649977179
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1649977179
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1649977179
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1649977179
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_169
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_177
timestamp 1649977179
transform 1 0 17388 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_186
timestamp 1649977179
transform 1 0 18216 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_195
timestamp 1649977179
transform 1 0 19044 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_207
timestamp 1649977179
transform 1 0 20148 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_219
timestamp 1649977179
transform 1 0 21252 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1649977179
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_225
timestamp 1649977179
transform 1 0 21804 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_233
timestamp 1649977179
transform 1 0 22540 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_245
timestamp 1649977179
transform 1 0 23644 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_257
timestamp 1649977179
transform 1 0 24748 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_269
timestamp 1649977179
transform 1 0 25852 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_277
timestamp 1649977179
transform 1 0 26588 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_281
timestamp 1649977179
transform 1 0 26956 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_287
timestamp 1649977179
transform 1 0 27508 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_299
timestamp 1649977179
transform 1 0 28612 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_313
timestamp 1649977179
transform 1 0 29900 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_325
timestamp 1649977179
transform 1 0 31004 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_333
timestamp 1649977179
transform 1 0 31740 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_337
timestamp 1649977179
transform 1 0 32108 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_343
timestamp 1649977179
transform 1 0 32660 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_352
timestamp 1649977179
transform 1 0 33488 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_364
timestamp 1649977179
transform 1 0 34592 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_376
timestamp 1649977179
transform 1 0 35696 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_380
timestamp 1649977179
transform 1 0 36064 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1649977179
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_405
timestamp 1649977179
transform 1 0 38364 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1649977179
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1649977179
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1649977179
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_29
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_42
timestamp 1649977179
transform 1 0 4968 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_54
timestamp 1649977179
transform 1 0 6072 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_66
timestamp 1649977179
transform 1 0 7176 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_70
timestamp 1649977179
transform 1 0 7544 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1649977179
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_90
timestamp 1649977179
transform 1 0 9384 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_102
timestamp 1649977179
transform 1 0 10488 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_114
timestamp 1649977179
transform 1 0 11592 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_126
timestamp 1649977179
transform 1 0 12696 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1649977179
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_141
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_147
timestamp 1649977179
transform 1 0 14628 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_151
timestamp 1649977179
transform 1 0 14996 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_157
timestamp 1649977179
transform 1 0 15548 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_169
timestamp 1649977179
transform 1 0 16652 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_181
timestamp 1649977179
transform 1 0 17756 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_193
timestamp 1649977179
transform 1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1649977179
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1649977179
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_233
timestamp 1649977179
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1649977179
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1649977179
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_253
timestamp 1649977179
transform 1 0 24380 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_266
timestamp 1649977179
transform 1 0 25576 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_278
timestamp 1649977179
transform 1 0 26680 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_285
timestamp 1649977179
transform 1 0 27324 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_28_296
timestamp 1649977179
transform 1 0 28336 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1649977179
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1649977179
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1649977179
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1649977179
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1649977179
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1649977179
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1649977179
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1649977179
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1649977179
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_401
timestamp 1649977179
transform 1 0 37996 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_7
timestamp 1649977179
transform 1 0 1748 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_13
timestamp 1649977179
transform 1 0 2300 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_31
timestamp 1649977179
transform 1 0 3956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_43
timestamp 1649977179
transform 1 0 5060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1649977179
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_57
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_68
timestamp 1649977179
transform 1 0 7360 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_72
timestamp 1649977179
transform 1 0 7728 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1649977179
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1649977179
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1649977179
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_125
timestamp 1649977179
transform 1 0 12604 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_131
timestamp 1649977179
transform 1 0 13156 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_137
timestamp 1649977179
transform 1 0 13708 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_147
timestamp 1649977179
transform 1 0 14628 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_159
timestamp 1649977179
transform 1 0 15732 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1649977179
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1649977179
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1649977179
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1649977179
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1649977179
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1649977179
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1649977179
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1649977179
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1649977179
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_261
timestamp 1649977179
transform 1 0 25116 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_265
timestamp 1649977179
transform 1 0 25484 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_277
timestamp 1649977179
transform 1 0 26588 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1649977179
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1649977179
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1649977179
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1649977179
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1649977179
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1649977179
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1649977179
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1649977179
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1649977179
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1649977179
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1649977179
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1649977179
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1649977179
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_405
timestamp 1649977179
transform 1 0 38364 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1649977179
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1649977179
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1649977179
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_32
timestamp 1649977179
transform 1 0 4048 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_44
timestamp 1649977179
transform 1 0 5152 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_56
timestamp 1649977179
transform 1 0 6256 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_69
timestamp 1649977179
transform 1 0 7452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_81
timestamp 1649977179
transform 1 0 8556 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_85
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_93
timestamp 1649977179
transform 1 0 9660 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_98
timestamp 1649977179
transform 1 0 10120 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_102
timestamp 1649977179
transform 1 0 10488 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_123
timestamp 1649977179
transform 1 0 12420 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_135
timestamp 1649977179
transform 1 0 13524 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1649977179
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1649977179
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1649977179
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1649977179
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1649977179
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1649977179
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_209
timestamp 1649977179
transform 1 0 20332 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_227
timestamp 1649977179
transform 1 0 21988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_239
timestamp 1649977179
transform 1 0 23092 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1649977179
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_258
timestamp 1649977179
transform 1 0 24840 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_274
timestamp 1649977179
transform 1 0 26312 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_286
timestamp 1649977179
transform 1 0 27416 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_298
timestamp 1649977179
transform 1 0 28520 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_306
timestamp 1649977179
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1649977179
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1649977179
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1649977179
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1649977179
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1649977179
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1649977179
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1649977179
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_377
timestamp 1649977179
transform 1 0 35788 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_385
timestamp 1649977179
transform 1 0 36524 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_398
timestamp 1649977179
transform 1 0 37720 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_406
timestamp 1649977179
transform 1 0 38456 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1649977179
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_15
timestamp 1649977179
transform 1 0 2484 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_28
timestamp 1649977179
transform 1 0 3680 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_34
timestamp 1649977179
transform 1 0 4232 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_46
timestamp 1649977179
transform 1 0 5336 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1649977179
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_57
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_66
timestamp 1649977179
transform 1 0 7176 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_78
timestamp 1649977179
transform 1 0 8280 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_90
timestamp 1649977179
transform 1 0 9384 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_96
timestamp 1649977179
transform 1 0 9936 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_100
timestamp 1649977179
transform 1 0 10304 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_106
timestamp 1649977179
transform 1 0 10856 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1649977179
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1649977179
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1649977179
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1649977179
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1649977179
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_174
timestamp 1649977179
transform 1 0 17112 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_186
timestamp 1649977179
transform 1 0 18216 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_198
timestamp 1649977179
transform 1 0 19320 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_210
timestamp 1649977179
transform 1 0 20424 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1649977179
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_228
timestamp 1649977179
transform 1 0 22080 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_240
timestamp 1649977179
transform 1 0 23184 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_252
timestamp 1649977179
transform 1 0 24288 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_260
timestamp 1649977179
transform 1 0 25024 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_266
timestamp 1649977179
transform 1 0 25576 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1649977179
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1649977179
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1649977179
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1649977179
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_305
timestamp 1649977179
transform 1 0 29164 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_309
timestamp 1649977179
transform 1 0 29532 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_322
timestamp 1649977179
transform 1 0 30728 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_334
timestamp 1649977179
transform 1 0 31832 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1649977179
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_349
timestamp 1649977179
transform 1 0 33212 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_369
timestamp 1649977179
transform 1 0 35052 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_381
timestamp 1649977179
transform 1 0 36156 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_389
timestamp 1649977179
transform 1 0 36892 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1649977179
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_405
timestamp 1649977179
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_7
timestamp 1649977179
transform 1 0 1748 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_13
timestamp 1649977179
transform 1 0 2300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_25
timestamp 1649977179
transform 1 0 3404 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1649977179
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_53
timestamp 1649977179
transform 1 0 5980 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_57
timestamp 1649977179
transform 1 0 6348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_61
timestamp 1649977179
transform 1 0 6716 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_73
timestamp 1649977179
transform 1 0 7820 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_81
timestamp 1649977179
transform 1 0 8556 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1649977179
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1649977179
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1649977179
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1649977179
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1649977179
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_141
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_147
timestamp 1649977179
transform 1 0 14628 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_156
timestamp 1649977179
transform 1 0 15456 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_172
timestamp 1649977179
transform 1 0 16928 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_179
timestamp 1649977179
transform 1 0 17572 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_191
timestamp 1649977179
transform 1 0 18676 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1649977179
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_209
timestamp 1649977179
transform 1 0 20332 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_213
timestamp 1649977179
transform 1 0 20700 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_222
timestamp 1649977179
transform 1 0 21528 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_234
timestamp 1649977179
transform 1 0 22632 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_246
timestamp 1649977179
transform 1 0 23736 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1649977179
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1649977179
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1649977179
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1649977179
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1649977179
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1649977179
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_309
timestamp 1649977179
transform 1 0 29532 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_322
timestamp 1649977179
transform 1 0 30728 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_334
timestamp 1649977179
transform 1 0 31832 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_346
timestamp 1649977179
transform 1 0 32936 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_354
timestamp 1649977179
transform 1 0 33672 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_359
timestamp 1649977179
transform 1 0 34132 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1649977179
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_365
timestamp 1649977179
transform 1 0 34684 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_373
timestamp 1649977179
transform 1 0 35420 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_388
timestamp 1649977179
transform 1 0 36800 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_400
timestamp 1649977179
transform 1 0 37904 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_406
timestamp 1649977179
transform 1 0 38456 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_3
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_9
timestamp 1649977179
transform 1 0 1932 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_21
timestamp 1649977179
transform 1 0 3036 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_33
timestamp 1649977179
transform 1 0 4140 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_45
timestamp 1649977179
transform 1 0 5244 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_53
timestamp 1649977179
transform 1 0 5980 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_69
timestamp 1649977179
transform 1 0 7452 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_74
timestamp 1649977179
transform 1 0 7912 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_98
timestamp 1649977179
transform 1 0 10120 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1649977179
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1649977179
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1649977179
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1649977179
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1649977179
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1649977179
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_169
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_182
timestamp 1649977179
transform 1 0 17848 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_188
timestamp 1649977179
transform 1 0 18400 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_196
timestamp 1649977179
transform 1 0 19136 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_204
timestamp 1649977179
transform 1 0 19872 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_216
timestamp 1649977179
transform 1 0 20976 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1649977179
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1649977179
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1649977179
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_261
timestamp 1649977179
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1649977179
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1649977179
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1649977179
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1649977179
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_305
timestamp 1649977179
transform 1 0 29164 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_312
timestamp 1649977179
transform 1 0 29808 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_321
timestamp 1649977179
transform 1 0 30636 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_333
timestamp 1649977179
transform 1 0 31740 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_337
timestamp 1649977179
transform 1 0 32108 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_345
timestamp 1649977179
transform 1 0 32844 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_353
timestamp 1649977179
transform 1 0 33580 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_357
timestamp 1649977179
transform 1 0 33948 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_363
timestamp 1649977179
transform 1 0 34500 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_372
timestamp 1649977179
transform 1 0 35328 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_384
timestamp 1649977179
transform 1 0 36432 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1649977179
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_405
timestamp 1649977179
transform 1 0 38364 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_7
timestamp 1649977179
transform 1 0 1748 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_11
timestamp 1649977179
transform 1 0 2116 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_24
timestamp 1649977179
transform 1 0 3312 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1649977179
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_41
timestamp 1649977179
transform 1 0 4876 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_57
timestamp 1649977179
transform 1 0 6348 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_73
timestamp 1649977179
transform 1 0 7820 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_81
timestamp 1649977179
transform 1 0 8556 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1649977179
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1649977179
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1649977179
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1649977179
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1649977179
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1649977179
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1649977179
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1649977179
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1649977179
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1649977179
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1649977179
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1649977179
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_199
timestamp 1649977179
transform 1 0 19412 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_217
timestamp 1649977179
transform 1 0 21068 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_229
timestamp 1649977179
transform 1 0 22172 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_241
timestamp 1649977179
transform 1 0 23276 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_249
timestamp 1649977179
transform 1 0 24012 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1649977179
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1649977179
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1649977179
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_289
timestamp 1649977179
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1649977179
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1649977179
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_309
timestamp 1649977179
transform 1 0 29532 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_314
timestamp 1649977179
transform 1 0 29992 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1649977179
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1649977179
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1649977179
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1649977179
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1649977179
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1649977179
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_377
timestamp 1649977179
transform 1 0 35788 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_382
timestamp 1649977179
transform 1 0 36248 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_394
timestamp 1649977179
transform 1 0 37352 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_406
timestamp 1649977179
transform 1 0 38456 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1649977179
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_15
timestamp 1649977179
transform 1 0 2484 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_22
timestamp 1649977179
transform 1 0 3128 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_34
timestamp 1649977179
transform 1 0 4232 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_46
timestamp 1649977179
transform 1 0 5336 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1649977179
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1649977179
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1649977179
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1649977179
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1649977179
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1649977179
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1649977179
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1649977179
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1649977179
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1649977179
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1649977179
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1649977179
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1649977179
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1649977179
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_181
timestamp 1649977179
transform 1 0 17756 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_189
timestamp 1649977179
transform 1 0 18492 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_196
timestamp 1649977179
transform 1 0 19136 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_207
timestamp 1649977179
transform 1 0 20148 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_219
timestamp 1649977179
transform 1 0 21252 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1649977179
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_225
timestamp 1649977179
transform 1 0 21804 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_232
timestamp 1649977179
transform 1 0 22448 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_240
timestamp 1649977179
transform 1 0 23184 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_246
timestamp 1649977179
transform 1 0 23736 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_258
timestamp 1649977179
transform 1 0 24840 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_264
timestamp 1649977179
transform 1 0 25392 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_276
timestamp 1649977179
transform 1 0 26496 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1649977179
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1649977179
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1649977179
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1649977179
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1649977179
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1649977179
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1649977179
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_349
timestamp 1649977179
transform 1 0 33212 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_359
timestamp 1649977179
transform 1 0 34132 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_368
timestamp 1649977179
transform 1 0 34960 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_380
timestamp 1649977179
transform 1 0 36064 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1649977179
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_405
timestamp 1649977179
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1649977179
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1649977179
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1649977179
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1649977179
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_41
timestamp 1649977179
transform 1 0 4876 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_49
timestamp 1649977179
transform 1 0 5612 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_54
timestamp 1649977179
transform 1 0 6072 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_62
timestamp 1649977179
transform 1 0 6808 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_66
timestamp 1649977179
transform 1 0 7176 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_78
timestamp 1649977179
transform 1 0 8280 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1649977179
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_97
timestamp 1649977179
transform 1 0 10028 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_110
timestamp 1649977179
transform 1 0 11224 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_117
timestamp 1649977179
transform 1 0 11868 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1649977179
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1649977179
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_141
timestamp 1649977179
transform 1 0 14076 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_152
timestamp 1649977179
transform 1 0 15088 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_164
timestamp 1649977179
transform 1 0 16192 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_176
timestamp 1649977179
transform 1 0 17296 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_188
timestamp 1649977179
transform 1 0 18400 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1649977179
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1649977179
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1649977179
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1649977179
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_248
timestamp 1649977179
transform 1 0 23920 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_265
timestamp 1649977179
transform 1 0 25484 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_269
timestamp 1649977179
transform 1 0 25852 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_283
timestamp 1649977179
transform 1 0 27140 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_295
timestamp 1649977179
transform 1 0 28244 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1649977179
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1649977179
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1649977179
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1649977179
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1649977179
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1649977179
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1649977179
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1649977179
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1649977179
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1649977179
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_401
timestamp 1649977179
transform 1 0 37996 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_6
timestamp 1649977179
transform 1 0 1656 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_18
timestamp 1649977179
transform 1 0 2760 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_25
timestamp 1649977179
transform 1 0 3404 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_31
timestamp 1649977179
transform 1 0 3956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_43
timestamp 1649977179
transform 1 0 5060 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1649977179
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_57
timestamp 1649977179
transform 1 0 6348 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_61
timestamp 1649977179
transform 1 0 6716 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_67
timestamp 1649977179
transform 1 0 7268 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_79
timestamp 1649977179
transform 1 0 8372 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_91
timestamp 1649977179
transform 1 0 9476 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_95
timestamp 1649977179
transform 1 0 9844 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_99
timestamp 1649977179
transform 1 0 10212 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1649977179
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_113
timestamp 1649977179
transform 1 0 11500 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_121
timestamp 1649977179
transform 1 0 12236 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_128
timestamp 1649977179
transform 1 0 12880 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_135
timestamp 1649977179
transform 1 0 13524 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_147
timestamp 1649977179
transform 1 0 14628 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_159
timestamp 1649977179
transform 1 0 15732 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1649977179
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_174
timestamp 1649977179
transform 1 0 17112 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_180
timestamp 1649977179
transform 1 0 17664 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_192
timestamp 1649977179
transform 1 0 18768 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_204
timestamp 1649977179
transform 1 0 19872 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_216
timestamp 1649977179
transform 1 0 20976 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1649977179
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1649977179
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1649977179
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_261
timestamp 1649977179
transform 1 0 25116 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_37_270
timestamp 1649977179
transform 1 0 25944 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_278
timestamp 1649977179
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1649977179
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1649977179
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1649977179
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1649977179
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1649977179
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1649977179
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1649977179
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1649977179
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1649977179
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1649977179
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1649977179
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1649977179
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1649977179
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_405
timestamp 1649977179
transform 1 0 38364 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1649977179
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1649977179
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1649977179
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1649977179
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_41
timestamp 1649977179
transform 1 0 4876 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_47
timestamp 1649977179
transform 1 0 5428 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1649977179
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1649977179
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1649977179
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1649977179
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_85
timestamp 1649977179
transform 1 0 8924 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_91
timestamp 1649977179
transform 1 0 9476 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_98
timestamp 1649977179
transform 1 0 10120 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_110
timestamp 1649977179
transform 1 0 11224 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_122
timestamp 1649977179
transform 1 0 12328 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_134
timestamp 1649977179
transform 1 0 13432 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1649977179
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_153
timestamp 1649977179
transform 1 0 15180 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_158
timestamp 1649977179
transform 1 0 15640 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_174
timestamp 1649977179
transform 1 0 17112 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_186
timestamp 1649977179
transform 1 0 18216 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1649977179
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1649977179
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1649977179
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1649977179
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_233
timestamp 1649977179
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1649977179
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1649977179
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1649977179
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1649977179
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1649977179
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1649977179
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1649977179
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1649977179
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1649977179
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_321
timestamp 1649977179
transform 1 0 30636 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_334
timestamp 1649977179
transform 1 0 31832 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_346
timestamp 1649977179
transform 1 0 32936 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_358
timestamp 1649977179
transform 1 0 34040 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_365
timestamp 1649977179
transform 1 0 34684 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_373
timestamp 1649977179
transform 1 0 35420 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1649977179
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1649977179
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_401
timestamp 1649977179
transform 1 0 37996 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_7
timestamp 1649977179
transform 1 0 1748 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_31
timestamp 1649977179
transform 1 0 3956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_43
timestamp 1649977179
transform 1 0 5060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1649977179
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1649977179
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_69
timestamp 1649977179
transform 1 0 7452 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_76
timestamp 1649977179
transform 1 0 8096 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_92
timestamp 1649977179
transform 1 0 9568 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_98
timestamp 1649977179
transform 1 0 10120 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1649977179
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1649977179
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_125
timestamp 1649977179
transform 1 0 12604 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_135
timestamp 1649977179
transform 1 0 13524 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_141
timestamp 1649977179
transform 1 0 14076 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_153
timestamp 1649977179
transform 1 0 15180 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_165
timestamp 1649977179
transform 1 0 16284 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_172
timestamp 1649977179
transform 1 0 16928 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_184
timestamp 1649977179
transform 1 0 18032 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_196
timestamp 1649977179
transform 1 0 19136 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_39_216
timestamp 1649977179
transform 1 0 20976 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1649977179
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1649977179
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1649977179
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1649977179
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1649977179
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1649977179
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_281
timestamp 1649977179
transform 1 0 26956 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_301
timestamp 1649977179
transform 1 0 28796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_308
timestamp 1649977179
transform 1 0 29440 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_318
timestamp 1649977179
transform 1 0 30360 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_332
timestamp 1649977179
transform 1 0 31648 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_337
timestamp 1649977179
transform 1 0 32108 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_341
timestamp 1649977179
transform 1 0 32476 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_347
timestamp 1649977179
transform 1 0 33028 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_355
timestamp 1649977179
transform 1 0 33764 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_360
timestamp 1649977179
transform 1 0 34224 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_369
timestamp 1649977179
transform 1 0 35052 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_388
timestamp 1649977179
transform 1 0 36800 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1649977179
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_405
timestamp 1649977179
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1649977179
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_15
timestamp 1649977179
transform 1 0 2484 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_24
timestamp 1649977179
transform 1 0 3312 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_34
timestamp 1649977179
transform 1 0 4232 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_40
timestamp 1649977179
transform 1 0 4784 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_52
timestamp 1649977179
transform 1 0 5888 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_64
timestamp 1649977179
transform 1 0 6992 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_76
timestamp 1649977179
transform 1 0 8096 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_40_95
timestamp 1649977179
transform 1 0 9844 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_107
timestamp 1649977179
transform 1 0 10948 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_119
timestamp 1649977179
transform 1 0 12052 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_131
timestamp 1649977179
transform 1 0 13156 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1649977179
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1649977179
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1649977179
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1649977179
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1649977179
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1649977179
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1649977179
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_197
timestamp 1649977179
transform 1 0 19228 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_200
timestamp 1649977179
transform 1 0 19504 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_209
timestamp 1649977179
transform 1 0 20332 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_216
timestamp 1649977179
transform 1 0 20976 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_228
timestamp 1649977179
transform 1 0 22080 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_240
timestamp 1649977179
transform 1 0 23184 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1649977179
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1649977179
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1649977179
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_289
timestamp 1649977179
transform 1 0 27692 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_40_302
timestamp 1649977179
transform 1 0 28888 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1649977179
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_321
timestamp 1649977179
transform 1 0 30636 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_329
timestamp 1649977179
transform 1 0 31372 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_335
timestamp 1649977179
transform 1 0 31924 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_343
timestamp 1649977179
transform 1 0 32660 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_358
timestamp 1649977179
transform 1 0 34040 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1649977179
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1649977179
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1649977179
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_401
timestamp 1649977179
transform 1 0 37996 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1649977179
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1649977179
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1649977179
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1649977179
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1649977179
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1649977179
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1649977179
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1649977179
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1649977179
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1649977179
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1649977179
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1649977179
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1649977179
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_129
timestamp 1649977179
transform 1 0 12972 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_135
timestamp 1649977179
transform 1 0 13524 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_143
timestamp 1649977179
transform 1 0 14260 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_146
timestamp 1649977179
transform 1 0 14536 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_155
timestamp 1649977179
transform 1 0 15364 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_162
timestamp 1649977179
transform 1 0 16008 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1649977179
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1649977179
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1649977179
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_208
timestamp 1649977179
transform 1 0 20240 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_220
timestamp 1649977179
transform 1 0 21344 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_228
timestamp 1649977179
transform 1 0 22080 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_240
timestamp 1649977179
transform 1 0 23184 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_252
timestamp 1649977179
transform 1 0 24288 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_264
timestamp 1649977179
transform 1 0 25392 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_276
timestamp 1649977179
transform 1 0 26496 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1649977179
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_293
timestamp 1649977179
transform 1 0 28060 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_301
timestamp 1649977179
transform 1 0 28796 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_313
timestamp 1649977179
transform 1 0 29900 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_325
timestamp 1649977179
transform 1 0 31004 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_333
timestamp 1649977179
transform 1 0 31740 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_337
timestamp 1649977179
transform 1 0 32108 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_345
timestamp 1649977179
transform 1 0 32844 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_349
timestamp 1649977179
transform 1 0 33212 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_356
timestamp 1649977179
transform 1 0 33856 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_368
timestamp 1649977179
transform 1 0 34960 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_380
timestamp 1649977179
transform 1 0 36064 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1649977179
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_405
timestamp 1649977179
transform 1 0 38364 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_7
timestamp 1649977179
transform 1 0 1748 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_13
timestamp 1649977179
transform 1 0 2300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_25
timestamp 1649977179
transform 1 0 3404 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1649977179
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1649977179
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1649977179
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1649977179
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1649977179
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1649977179
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1649977179
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1649977179
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1649977179
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_126
timestamp 1649977179
transform 1 0 12696 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_138
timestamp 1649977179
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1649977179
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_153
timestamp 1649977179
transform 1 0 15180 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_169
timestamp 1649977179
transform 1 0 16652 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_181
timestamp 1649977179
transform 1 0 17756 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_193
timestamp 1649977179
transform 1 0 18860 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_197
timestamp 1649977179
transform 1 0 19228 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_205
timestamp 1649977179
transform 1 0 19964 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_210
timestamp 1649977179
transform 1 0 20424 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_219
timestamp 1649977179
transform 1 0 21252 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_237
timestamp 1649977179
transform 1 0 22908 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_249
timestamp 1649977179
transform 1 0 24012 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_256
timestamp 1649977179
transform 1 0 24656 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_268
timestamp 1649977179
transform 1 0 25760 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_280
timestamp 1649977179
transform 1 0 26864 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_286
timestamp 1649977179
transform 1 0 27416 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_299
timestamp 1649977179
transform 1 0 28612 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1649977179
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1649977179
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1649977179
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1649977179
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1649977179
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1649977179
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1649977179
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1649977179
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1649977179
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1649977179
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_401
timestamp 1649977179
transform 1 0 37996 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1649977179
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_17
timestamp 1649977179
transform 1 0 2668 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_29
timestamp 1649977179
transform 1 0 3772 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_41
timestamp 1649977179
transform 1 0 4876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_53
timestamp 1649977179
transform 1 0 5980 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_57
timestamp 1649977179
transform 1 0 6348 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_65
timestamp 1649977179
transform 1 0 7084 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_73
timestamp 1649977179
transform 1 0 7820 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_85
timestamp 1649977179
transform 1 0 8924 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_97
timestamp 1649977179
transform 1 0 10028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_109
timestamp 1649977179
transform 1 0 11132 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_113
timestamp 1649977179
transform 1 0 11500 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_127
timestamp 1649977179
transform 1 0 12788 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_139
timestamp 1649977179
transform 1 0 13892 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_151
timestamp 1649977179
transform 1 0 14996 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_43_162
timestamp 1649977179
transform 1 0 16008 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1649977179
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1649977179
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1649977179
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1649977179
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1649977179
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1649977179
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1649977179
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1649977179
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_249
timestamp 1649977179
transform 1 0 24012 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_264
timestamp 1649977179
transform 1 0 25392 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1649977179
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1649977179
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_283
timestamp 1649977179
transform 1 0 27140 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_298
timestamp 1649977179
transform 1 0 28520 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_310
timestamp 1649977179
transform 1 0 29624 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_322
timestamp 1649977179
transform 1 0 30728 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_334
timestamp 1649977179
transform 1 0 31832 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1649977179
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1649977179
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1649977179
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1649977179
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1649977179
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1649977179
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1649977179
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_405
timestamp 1649977179
transform 1 0 38364 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_7
timestamp 1649977179
transform 1 0 1748 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_11
timestamp 1649977179
transform 1 0 2116 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_15
timestamp 1649977179
transform 1 0 2484 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_24
timestamp 1649977179
transform 1 0 3312 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_31
timestamp 1649977179
transform 1 0 3956 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_43
timestamp 1649977179
transform 1 0 5060 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_55
timestamp 1649977179
transform 1 0 6164 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_67
timestamp 1649977179
transform 1 0 7268 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_80
timestamp 1649977179
transform 1 0 8464 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1649977179
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1649977179
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_109
timestamp 1649977179
transform 1 0 11132 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_117
timestamp 1649977179
transform 1 0 11868 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_123
timestamp 1649977179
transform 1 0 12420 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_135
timestamp 1649977179
transform 1 0 13524 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1649977179
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_141
timestamp 1649977179
transform 1 0 14076 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_149
timestamp 1649977179
transform 1 0 14812 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_155
timestamp 1649977179
transform 1 0 15364 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_171
timestamp 1649977179
transform 1 0 16836 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_183
timestamp 1649977179
transform 1 0 17940 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1649977179
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_202
timestamp 1649977179
transform 1 0 19688 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_214
timestamp 1649977179
transform 1 0 20792 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_226
timestamp 1649977179
transform 1 0 21896 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_238
timestamp 1649977179
transform 1 0 23000 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_250
timestamp 1649977179
transform 1 0 24104 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_253
timestamp 1649977179
transform 1 0 24380 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_257
timestamp 1649977179
transform 1 0 24748 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_261
timestamp 1649977179
transform 1 0 25116 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_273
timestamp 1649977179
transform 1 0 26220 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_285
timestamp 1649977179
transform 1 0 27324 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_297
timestamp 1649977179
transform 1 0 28428 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_305
timestamp 1649977179
transform 1 0 29164 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1649977179
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_321
timestamp 1649977179
transform 1 0 30636 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_329
timestamp 1649977179
transform 1 0 31372 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_335
timestamp 1649977179
transform 1 0 31924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_347
timestamp 1649977179
transform 1 0 33028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_359
timestamp 1649977179
transform 1 0 34132 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1649977179
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1649977179
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1649977179
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1649977179
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_401
timestamp 1649977179
transform 1 0 37996 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1649977179
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1649977179
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_39
timestamp 1649977179
transform 1 0 4692 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_47
timestamp 1649977179
transform 1 0 5428 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1649977179
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1649977179
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1649977179
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_69
timestamp 1649977179
transform 1 0 7452 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_74
timestamp 1649977179
transform 1 0 7912 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_86
timestamp 1649977179
transform 1 0 9016 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_98
timestamp 1649977179
transform 1 0 10120 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_110
timestamp 1649977179
transform 1 0 11224 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1649977179
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1649977179
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1649977179
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_149
timestamp 1649977179
transform 1 0 14812 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_45_157
timestamp 1649977179
transform 1 0 15548 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_165
timestamp 1649977179
transform 1 0 16284 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1649977179
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1649977179
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1649977179
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_205
timestamp 1649977179
transform 1 0 19964 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_209
timestamp 1649977179
transform 1 0 20332 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_212
timestamp 1649977179
transform 1 0 20608 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1649977179
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_237
timestamp 1649977179
transform 1 0 22908 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_245
timestamp 1649977179
transform 1 0 23644 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_251
timestamp 1649977179
transform 1 0 24196 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_263
timestamp 1649977179
transform 1 0 25300 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_275
timestamp 1649977179
transform 1 0 26404 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1649977179
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1649977179
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_293
timestamp 1649977179
transform 1 0 28060 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_297
timestamp 1649977179
transform 1 0 28428 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_301
timestamp 1649977179
transform 1 0 28796 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_313
timestamp 1649977179
transform 1 0 29900 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_325
timestamp 1649977179
transform 1 0 31004 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_332
timestamp 1649977179
transform 1 0 31648 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_350
timestamp 1649977179
transform 1 0 33304 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_362
timestamp 1649977179
transform 1 0 34408 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_374
timestamp 1649977179
transform 1 0 35512 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_388
timestamp 1649977179
transform 1 0 36800 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1649977179
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_405
timestamp 1649977179
transform 1 0 38364 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1649977179
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_15
timestamp 1649977179
transform 1 0 2484 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_20
timestamp 1649977179
transform 1 0 2944 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1649977179
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_41
timestamp 1649977179
transform 1 0 4876 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_55
timestamp 1649977179
transform 1 0 6164 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_64
timestamp 1649977179
transform 1 0 6992 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_76
timestamp 1649977179
transform 1 0 8096 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_90
timestamp 1649977179
transform 1 0 9384 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_96
timestamp 1649977179
transform 1 0 9936 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_108
timestamp 1649977179
transform 1 0 11040 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_120
timestamp 1649977179
transform 1 0 12144 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_132
timestamp 1649977179
transform 1 0 13248 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1649977179
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1649977179
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1649977179
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1649977179
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1649977179
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1649977179
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_197
timestamp 1649977179
transform 1 0 19228 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_201
timestamp 1649977179
transform 1 0 19596 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_210
timestamp 1649977179
transform 1 0 20424 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_217
timestamp 1649977179
transform 1 0 21068 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_229
timestamp 1649977179
transform 1 0 22172 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_241
timestamp 1649977179
transform 1 0 23276 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_249
timestamp 1649977179
transform 1 0 24012 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_253
timestamp 1649977179
transform 1 0 24380 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_261
timestamp 1649977179
transform 1 0 25116 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_273
timestamp 1649977179
transform 1 0 26220 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_285
timestamp 1649977179
transform 1 0 27324 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_302
timestamp 1649977179
transform 1 0 28888 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1649977179
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_321
timestamp 1649977179
transform 1 0 30636 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_329
timestamp 1649977179
transform 1 0 31372 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_334
timestamp 1649977179
transform 1 0 31832 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_346
timestamp 1649977179
transform 1 0 32936 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_358
timestamp 1649977179
transform 1 0 34040 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_46_365
timestamp 1649977179
transform 1 0 34684 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_371
timestamp 1649977179
transform 1 0 35236 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_388
timestamp 1649977179
transform 1 0 36800 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_400
timestamp 1649977179
transform 1 0 37904 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_406
timestamp 1649977179
transform 1 0 38456 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_7
timestamp 1649977179
transform 1 0 1748 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_13
timestamp 1649977179
transform 1 0 2300 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_25
timestamp 1649977179
transform 1 0 3404 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_37
timestamp 1649977179
transform 1 0 4508 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_49
timestamp 1649977179
transform 1 0 5612 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1649977179
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1649977179
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_69
timestamp 1649977179
transform 1 0 7452 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_75
timestamp 1649977179
transform 1 0 8004 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_88
timestamp 1649977179
transform 1 0 9200 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_100
timestamp 1649977179
transform 1 0 10304 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1649977179
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_125
timestamp 1649977179
transform 1 0 12604 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_129
timestamp 1649977179
transform 1 0 12972 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_135
timestamp 1649977179
transform 1 0 13524 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_147
timestamp 1649977179
transform 1 0 14628 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_159
timestamp 1649977179
transform 1 0 15732 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1649977179
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1649977179
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1649977179
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_193
timestamp 1649977179
transform 1 0 18860 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_196
timestamp 1649977179
transform 1 0 19136 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_204
timestamp 1649977179
transform 1 0 19872 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_220
timestamp 1649977179
transform 1 0 21344 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1649977179
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1649977179
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_251
timestamp 1649977179
transform 1 0 24196 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_260
timestamp 1649977179
transform 1 0 25024 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_272
timestamp 1649977179
transform 1 0 26128 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1649977179
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_293
timestamp 1649977179
transform 1 0 28060 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_306
timestamp 1649977179
transform 1 0 29256 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_318
timestamp 1649977179
transform 1 0 30360 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_330
timestamp 1649977179
transform 1 0 31464 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1649977179
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_349
timestamp 1649977179
transform 1 0 33212 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_357
timestamp 1649977179
transform 1 0 33948 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_364
timestamp 1649977179
transform 1 0 34592 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_373
timestamp 1649977179
transform 1 0 35420 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_380
timestamp 1649977179
transform 1 0 36064 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1649977179
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_405
timestamp 1649977179
transform 1 0 38364 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1649977179
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1649977179
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1649977179
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1649977179
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1649977179
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1649977179
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1649977179
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1649977179
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1649977179
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_88
timestamp 1649977179
transform 1 0 9200 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_100
timestamp 1649977179
transform 1 0 10304 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_112
timestamp 1649977179
transform 1 0 11408 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_125
timestamp 1649977179
transform 1 0 12604 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_132
timestamp 1649977179
transform 1 0 13248 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_151
timestamp 1649977179
transform 1 0 14996 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_157
timestamp 1649977179
transform 1 0 15548 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_172
timestamp 1649977179
transform 1 0 16928 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_184
timestamp 1649977179
transform 1 0 18032 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_197
timestamp 1649977179
transform 1 0 19228 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_205
timestamp 1649977179
transform 1 0 19964 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_209
timestamp 1649977179
transform 1 0 20332 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_223
timestamp 1649977179
transform 1 0 21620 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_229
timestamp 1649977179
transform 1 0 22172 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_241
timestamp 1649977179
transform 1 0 23276 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_249
timestamp 1649977179
transform 1 0 24012 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1649977179
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1649977179
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1649977179
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1649977179
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1649977179
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1649977179
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1649977179
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_321
timestamp 1649977179
transform 1 0 30636 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_329
timestamp 1649977179
transform 1 0 31372 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_333
timestamp 1649977179
transform 1 0 31740 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_48_341
timestamp 1649977179
transform 1 0 32476 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_353
timestamp 1649977179
transform 1 0 33580 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_361
timestamp 1649977179
transform 1 0 34316 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_48_365
timestamp 1649977179
transform 1 0 34684 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_368
timestamp 1649977179
transform 1 0 34960 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_380
timestamp 1649977179
transform 1 0 36064 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_392
timestamp 1649977179
transform 1 0 37168 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_404
timestamp 1649977179
transform 1 0 38272 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_7
timestamp 1649977179
transform 1 0 1748 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_13
timestamp 1649977179
transform 1 0 2300 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_49_21
timestamp 1649977179
transform 1 0 3036 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_33
timestamp 1649977179
transform 1 0 4140 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_45
timestamp 1649977179
transform 1 0 5244 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_53
timestamp 1649977179
transform 1 0 5980 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1649977179
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1649977179
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1649977179
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1649977179
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1649977179
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1649977179
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_123
timestamp 1649977179
transform 1 0 12420 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_130
timestamp 1649977179
transform 1 0 13064 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_136
timestamp 1649977179
transform 1 0 13616 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_148
timestamp 1649977179
transform 1 0 14720 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_156
timestamp 1649977179
transform 1 0 15456 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_163
timestamp 1649977179
transform 1 0 16100 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1649977179
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_169
timestamp 1649977179
transform 1 0 16652 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_49_187
timestamp 1649977179
transform 1 0 18308 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_199
timestamp 1649977179
transform 1 0 19412 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_211
timestamp 1649977179
transform 1 0 20516 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1649977179
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1649977179
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1649977179
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_249
timestamp 1649977179
transform 1 0 24012 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_260
timestamp 1649977179
transform 1 0 25024 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_272
timestamp 1649977179
transform 1 0 26128 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1649977179
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_293
timestamp 1649977179
transform 1 0 28060 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_299
timestamp 1649977179
transform 1 0 28612 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1649977179
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_317
timestamp 1649977179
transform 1 0 30268 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_325
timestamp 1649977179
transform 1 0 31004 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_331
timestamp 1649977179
transform 1 0 31556 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1649977179
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_337
timestamp 1649977179
transform 1 0 32108 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_345
timestamp 1649977179
transform 1 0 32844 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_357
timestamp 1649977179
transform 1 0 33948 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_369
timestamp 1649977179
transform 1 0 35052 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_381
timestamp 1649977179
transform 1 0 36156 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_389
timestamp 1649977179
transform 1 0 36892 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1649977179
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_405
timestamp 1649977179
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1649977179
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_15
timestamp 1649977179
transform 1 0 2484 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_19
timestamp 1649977179
transform 1 0 2852 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1649977179
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_31
timestamp 1649977179
transform 1 0 3956 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_43
timestamp 1649977179
transform 1 0 5060 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_55
timestamp 1649977179
transform 1 0 6164 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_67
timestamp 1649977179
transform 1 0 7268 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_79
timestamp 1649977179
transform 1 0 8372 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1649977179
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1649977179
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1649977179
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_109
timestamp 1649977179
transform 1 0 11132 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_115
timestamp 1649977179
transform 1 0 11684 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_128
timestamp 1649977179
transform 1 0 12880 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1649977179
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1649977179
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1649977179
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1649977179
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1649977179
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1649977179
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1649977179
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1649977179
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1649977179
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_233
timestamp 1649977179
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1649977179
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1649977179
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_253
timestamp 1649977179
transform 1 0 24380 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_262
timestamp 1649977179
transform 1 0 25208 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_268
timestamp 1649977179
transform 1 0 25760 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_280
timestamp 1649977179
transform 1 0 26864 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_292
timestamp 1649977179
transform 1 0 27968 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1649977179
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1649977179
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_311
timestamp 1649977179
transform 1 0 29716 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_323
timestamp 1649977179
transform 1 0 30820 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_335
timestamp 1649977179
transform 1 0 31924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_347
timestamp 1649977179
transform 1 0 33028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_359
timestamp 1649977179
transform 1 0 34132 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1649977179
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1649977179
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1649977179
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1649977179
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_401
timestamp 1649977179
transform 1 0 37996 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1649977179
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_15
timestamp 1649977179
transform 1 0 2484 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_28
timestamp 1649977179
transform 1 0 3680 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_35
timestamp 1649977179
transform 1 0 4324 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_47
timestamp 1649977179
transform 1 0 5428 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1649977179
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1649977179
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1649977179
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1649977179
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1649977179
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1649977179
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1649977179
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_118
timestamp 1649977179
transform 1 0 11960 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_124
timestamp 1649977179
transform 1 0 12512 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_136
timestamp 1649977179
transform 1 0 13616 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_148
timestamp 1649977179
transform 1 0 14720 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_160
timestamp 1649977179
transform 1 0 15824 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1649977179
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1649977179
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1649977179
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1649977179
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1649977179
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1649977179
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1649977179
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1649977179
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_249
timestamp 1649977179
transform 1 0 24012 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_253
timestamp 1649977179
transform 1 0 24380 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_266
timestamp 1649977179
transform 1 0 25576 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_278
timestamp 1649977179
transform 1 0 26680 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1649977179
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1649977179
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1649977179
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_317
timestamp 1649977179
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1649977179
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1649977179
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1649977179
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1649977179
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1649977179
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1649977179
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1649977179
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1649977179
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1649977179
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_405
timestamp 1649977179
transform 1 0 38364 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_7
timestamp 1649977179
transform 1 0 1748 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_19
timestamp 1649977179
transform 1 0 2852 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1649977179
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_29
timestamp 1649977179
transform 1 0 3772 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_43
timestamp 1649977179
transform 1 0 5060 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_55
timestamp 1649977179
transform 1 0 6164 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_67
timestamp 1649977179
transform 1 0 7268 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_79
timestamp 1649977179
transform 1 0 8372 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1649977179
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_90
timestamp 1649977179
transform 1 0 9384 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_96
timestamp 1649977179
transform 1 0 9936 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_108
timestamp 1649977179
transform 1 0 11040 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_120
timestamp 1649977179
transform 1 0 12144 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_132
timestamp 1649977179
transform 1 0 13248 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1649977179
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_153
timestamp 1649977179
transform 1 0 15180 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_158
timestamp 1649977179
transform 1 0 15640 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_170
timestamp 1649977179
transform 1 0 16744 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_182
timestamp 1649977179
transform 1 0 17848 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_194
timestamp 1649977179
transform 1 0 18952 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1649977179
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_209
timestamp 1649977179
transform 1 0 20332 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_215
timestamp 1649977179
transform 1 0 20884 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_221
timestamp 1649977179
transform 1 0 21436 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_227
timestamp 1649977179
transform 1 0 21988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_239
timestamp 1649977179
transform 1 0 23092 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1649977179
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_253
timestamp 1649977179
transform 1 0 24380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_258
timestamp 1649977179
transform 1 0 24840 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1649977179
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1649977179
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_289
timestamp 1649977179
transform 1 0 27692 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_297
timestamp 1649977179
transform 1 0 28428 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_302
timestamp 1649977179
transform 1 0 28888 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_312
timestamp 1649977179
transform 1 0 29808 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_324
timestamp 1649977179
transform 1 0 30912 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_336
timestamp 1649977179
transform 1 0 32016 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_348
timestamp 1649977179
transform 1 0 33120 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_360
timestamp 1649977179
transform 1 0 34224 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1649977179
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1649977179
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1649977179
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_401
timestamp 1649977179
transform 1 0 37996 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1649977179
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_15
timestamp 1649977179
transform 1 0 2484 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_22
timestamp 1649977179
transform 1 0 3128 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_28
timestamp 1649977179
transform 1 0 3680 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_40
timestamp 1649977179
transform 1 0 4784 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_52
timestamp 1649977179
transform 1 0 5888 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_62
timestamp 1649977179
transform 1 0 6808 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_74
timestamp 1649977179
transform 1 0 7912 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_87
timestamp 1649977179
transform 1 0 9108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_99
timestamp 1649977179
transform 1 0 10212 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1649977179
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_113
timestamp 1649977179
transform 1 0 11500 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_118
timestamp 1649977179
transform 1 0 11960 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_130
timestamp 1649977179
transform 1 0 13064 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_142
timestamp 1649977179
transform 1 0 14168 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_148
timestamp 1649977179
transform 1 0 14720 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_154
timestamp 1649977179
transform 1 0 15272 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_163
timestamp 1649977179
transform 1 0 16100 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1649977179
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_172
timestamp 1649977179
transform 1 0 16928 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_184
timestamp 1649977179
transform 1 0 18032 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_196
timestamp 1649977179
transform 1 0 19136 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_202
timestamp 1649977179
transform 1 0 19688 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_211
timestamp 1649977179
transform 1 0 20516 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1649977179
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_228
timestamp 1649977179
transform 1 0 22080 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_240
timestamp 1649977179
transform 1 0 23184 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_252
timestamp 1649977179
transform 1 0 24288 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_264
timestamp 1649977179
transform 1 0 25392 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_276
timestamp 1649977179
transform 1 0 26496 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1649977179
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_293
timestamp 1649977179
transform 1 0 28060 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_307
timestamp 1649977179
transform 1 0 29348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_319
timestamp 1649977179
transform 1 0 30452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_331
timestamp 1649977179
transform 1 0 31556 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1649977179
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1649977179
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1649977179
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1649977179
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1649977179
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1649977179
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1649977179
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1649977179
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_405
timestamp 1649977179
transform 1 0 38364 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_7
timestamp 1649977179
transform 1 0 1748 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_13
timestamp 1649977179
transform 1 0 2300 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_20
timestamp 1649977179
transform 1 0 2944 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1649977179
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1649977179
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_53
timestamp 1649977179
transform 1 0 5980 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_57
timestamp 1649977179
transform 1 0 6348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_61
timestamp 1649977179
transform 1 0 6716 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_73
timestamp 1649977179
transform 1 0 7820 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_81
timestamp 1649977179
transform 1 0 8556 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_88
timestamp 1649977179
transform 1 0 9200 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_100
timestamp 1649977179
transform 1 0 10304 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_112
timestamp 1649977179
transform 1 0 11408 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_125
timestamp 1649977179
transform 1 0 12604 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_137
timestamp 1649977179
transform 1 0 13708 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1649977179
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_153
timestamp 1649977179
transform 1 0 15180 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_161
timestamp 1649977179
transform 1 0 15916 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_54_167
timestamp 1649977179
transform 1 0 16468 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_175
timestamp 1649977179
transform 1 0 17204 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_188
timestamp 1649977179
transform 1 0 18400 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1649977179
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_209
timestamp 1649977179
transform 1 0 20332 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_216
timestamp 1649977179
transform 1 0 20976 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_232
timestamp 1649977179
transform 1 0 22448 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_248
timestamp 1649977179
transform 1 0 23920 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_253
timestamp 1649977179
transform 1 0 24380 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_259
timestamp 1649977179
transform 1 0 24932 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_272
timestamp 1649977179
transform 1 0 26128 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_284
timestamp 1649977179
transform 1 0 27232 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_304
timestamp 1649977179
transform 1 0 29072 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1649977179
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1649977179
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1649977179
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1649977179
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1649977179
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1649977179
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1649977179
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1649977179
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1649977179
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_401
timestamp 1649977179
transform 1 0 37996 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1649977179
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_15
timestamp 1649977179
transform 1 0 2484 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_28
timestamp 1649977179
transform 1 0 3680 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_40
timestamp 1649977179
transform 1 0 4784 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_52
timestamp 1649977179
transform 1 0 5888 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_57
timestamp 1649977179
transform 1 0 6348 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_70
timestamp 1649977179
transform 1 0 7544 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_82
timestamp 1649977179
transform 1 0 8648 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_94
timestamp 1649977179
transform 1 0 9752 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_108
timestamp 1649977179
transform 1 0 11040 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_130
timestamp 1649977179
transform 1 0 13064 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_142
timestamp 1649977179
transform 1 0 14168 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_154
timestamp 1649977179
transform 1 0 15272 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_166
timestamp 1649977179
transform 1 0 16376 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1649977179
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1649977179
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1649977179
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1649977179
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1649977179
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1649977179
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1649977179
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1649977179
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1649977179
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1649977179
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1649977179
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1649977179
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1649977179
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1649977179
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1649977179
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1649977179
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1649977179
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1649977179
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1649977179
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1649977179
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1649977179
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1649977179
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1649977179
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_393
timestamp 1649977179
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_405
timestamp 1649977179
transform 1 0 38364 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_7
timestamp 1649977179
transform 1 0 1748 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_13
timestamp 1649977179
transform 1 0 2300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_25
timestamp 1649977179
transform 1 0 3404 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1649977179
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1649977179
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1649977179
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1649977179
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1649977179
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1649977179
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_85
timestamp 1649977179
transform 1 0 8924 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_89
timestamp 1649977179
transform 1 0 9292 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_101
timestamp 1649977179
transform 1 0 10396 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_123
timestamp 1649977179
transform 1 0 12420 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_135
timestamp 1649977179
transform 1 0 13524 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1649977179
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1649977179
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1649977179
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1649977179
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1649977179
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1649977179
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1649977179
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1649977179
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1649977179
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1649977179
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1649977179
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1649977179
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1649977179
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1649977179
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1649977179
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1649977179
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1649977179
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1649977179
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1649977179
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1649977179
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1649977179
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1649977179
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1649977179
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1649977179
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1649977179
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1649977179
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1649977179
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1649977179
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_401
timestamp 1649977179
transform 1 0 37996 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_7
timestamp 1649977179
transform 1 0 1748 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_13
timestamp 1649977179
transform 1 0 2300 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_25
timestamp 1649977179
transform 1 0 3404 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_29
timestamp 1649977179
transform 1 0 3772 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_41
timestamp 1649977179
transform 1 0 4876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_53
timestamp 1649977179
transform 1 0 5980 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1649977179
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1649977179
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_81
timestamp 1649977179
transform 1 0 8556 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_85
timestamp 1649977179
transform 1 0 8924 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1649977179
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1649977179
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1649977179
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1649977179
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1649977179
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_137
timestamp 1649977179
transform 1 0 13708 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_141
timestamp 1649977179
transform 1 0 14076 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_153
timestamp 1649977179
transform 1 0 15180 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_165
timestamp 1649977179
transform 1 0 16284 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1649977179
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1649977179
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_193
timestamp 1649977179
transform 1 0 18860 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_57_197
timestamp 1649977179
transform 1 0 19228 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_205
timestamp 1649977179
transform 1 0 19964 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_209
timestamp 1649977179
transform 1 0 20332 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_221
timestamp 1649977179
transform 1 0 21436 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1649977179
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1649977179
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_249
timestamp 1649977179
transform 1 0 24012 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_253
timestamp 1649977179
transform 1 0 24380 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_265
timestamp 1649977179
transform 1 0 25484 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_57_271
timestamp 1649977179
transform 1 0 26036 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1649977179
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1649977179
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1649977179
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_305
timestamp 1649977179
transform 1 0 29164 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_309
timestamp 1649977179
transform 1 0 29532 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_321
timestamp 1649977179
transform 1 0 30636 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_333
timestamp 1649977179
transform 1 0 31740 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_340
timestamp 1649977179
transform 1 0 32384 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_352
timestamp 1649977179
transform 1 0 33488 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_365
timestamp 1649977179
transform 1 0 34684 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_377
timestamp 1649977179
transform 1 0 35788 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_389
timestamp 1649977179
transform 1 0 36892 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_57_396
timestamp 1649977179
transform 1 0 37536 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_404
timestamp 1649977179
transform 1 0 38272 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1649977179
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1649977179
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1649977179
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1649977179
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1649977179
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1649977179
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1649977179
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1649977179
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1649977179
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1649977179
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1649977179
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1649977179
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1649977179
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1649977179
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1649977179
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1649977179
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1649977179
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1649977179
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1649977179
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1649977179
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1649977179
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1649977179
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1649977179
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1649977179
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1649977179
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1649977179
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1649977179
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1649977179
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1649977179
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1649977179
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1649977179
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1649977179
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1649977179
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1649977179
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1649977179
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1649977179
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1649977179
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1649977179
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1649977179
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1649977179
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1649977179
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1649977179
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1649977179
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1649977179
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1649977179
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1649977179
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1649977179
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1649977179
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1649977179
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1649977179
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1649977179
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1649977179
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1649977179
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1649977179
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1649977179
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1649977179
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1649977179
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1649977179
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1649977179
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1649977179
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1649977179
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1649977179
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1649977179
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1649977179
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1649977179
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1649977179
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1649977179
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1649977179
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1649977179
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1649977179
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1649977179
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1649977179
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1649977179
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1649977179
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1649977179
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1649977179
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1649977179
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1649977179
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1649977179
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1649977179
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1649977179
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1649977179
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1649977179
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1649977179
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1649977179
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1649977179
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1649977179
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1649977179
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1649977179
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1649977179
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1649977179
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1649977179
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1649977179
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1649977179
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1649977179
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1649977179
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1649977179
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1649977179
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1649977179
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1649977179
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1649977179
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1649977179
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1649977179
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1649977179
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1649977179
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1649977179
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1649977179
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1649977179
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1649977179
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1649977179
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1649977179
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1649977179
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1649977179
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1649977179
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1649977179
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1649977179
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1649977179
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1649977179
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1649977179
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1649977179
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1649977179
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1649977179
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1649977179
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1649977179
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1649977179
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1649977179
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1649977179
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1649977179
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1649977179
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1649977179
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1649977179
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1649977179
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1649977179
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1649977179
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1649977179
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1649977179
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1649977179
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1649977179
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1649977179
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1649977179
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1649977179
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1649977179
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1649977179
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1649977179
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1649977179
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1649977179
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1649977179
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1649977179
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1649977179
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1649977179
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1649977179
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1649977179
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1649977179
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1649977179
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1649977179
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1649977179
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1649977179
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1649977179
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1649977179
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1649977179
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1649977179
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1649977179
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1649977179
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1649977179
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1649977179
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1649977179
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1649977179
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1649977179
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1649977179
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1649977179
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1649977179
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1649977179
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1649977179
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1649977179
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1649977179
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1649977179
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1649977179
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1649977179
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1649977179
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1649977179
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1649977179
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1649977179
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1649977179
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1649977179
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1649977179
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1649977179
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1649977179
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1649977179
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1649977179
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1649977179
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1649977179
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1649977179
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1649977179
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1649977179
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1649977179
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1649977179
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1649977179
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1649977179
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1649977179
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1649977179
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1649977179
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1649977179
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1649977179
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1649977179
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1649977179
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1649977179
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1649977179
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1649977179
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1649977179
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1649977179
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1649977179
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1649977179
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1649977179
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1649977179
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1649977179
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1649977179
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1649977179
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1649977179
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1649977179
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1649977179
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1649977179
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1649977179
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1649977179
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1649977179
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1649977179
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1649977179
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1649977179
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1649977179
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1649977179
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1649977179
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1649977179
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1649977179
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1649977179
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1649977179
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1649977179
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1649977179
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1649977179
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1649977179
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1649977179
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1649977179
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1649977179
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1649977179
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1649977179
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1649977179
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1649977179
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1649977179
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1649977179
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1649977179
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1649977179
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1649977179
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1649977179
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1649977179
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1649977179
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1649977179
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1649977179
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1649977179
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1649977179
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1649977179
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1649977179
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1649977179
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1649977179
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1649977179
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1649977179
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1649977179
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1649977179
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1649977179
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1649977179
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1649977179
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1649977179
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1649977179
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1649977179
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1649977179
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1649977179
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1649977179
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1649977179
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1649977179
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1649977179
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1649977179
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1649977179
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1649977179
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1649977179
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1649977179
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1649977179
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1649977179
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1649977179
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1649977179
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1649977179
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1649977179
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1649977179
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1649977179
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1649977179
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1649977179
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1649977179
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1649977179
transform 1 0 3680 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1649977179
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1649977179
transform 1 0 8832 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1649977179
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1649977179
transform 1 0 13984 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1649977179
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1649977179
transform 1 0 19136 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1649977179
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1649977179
transform 1 0 24288 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1649977179
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1649977179
transform 1 0 29440 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1649977179
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1649977179
transform 1 0 34592 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1649977179
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _293_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2944 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _294_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10120 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _295_
timestamp 1649977179
transform 1 0 17480 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _296_
timestamp 1649977179
transform 1 0 9660 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _297_
timestamp 1649977179
transform 1 0 16468 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _298_
timestamp 1649977179
transform -1 0 16100 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__and3b_1  _299_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 22908 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _300_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15824 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _301_
timestamp 1649977179
transform 1 0 19780 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _302_
timestamp 1649977179
transform 1 0 12052 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _303_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 18768 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _304_
timestamp 1649977179
transform 1 0 17848 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__and4b_1  _305_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 21804 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _306_
timestamp 1649977179
transform 1 0 15180 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__and4b_1  _307_
timestamp 1649977179
transform 1 0 21804 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nor4_1  _308_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 22632 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _309_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14720 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _310_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 14628 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _311_
timestamp 1649977179
transform 1 0 17572 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _312_
timestamp 1649977179
transform 1 0 17480 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _313_
timestamp 1649977179
transform -1 0 13616 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__a41o_1  _314_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _315_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13800 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _316_
timestamp 1649977179
transform -1 0 13248 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _317_
timestamp 1649977179
transform 1 0 6348 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _318_
timestamp 1649977179
transform 1 0 14444 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _319_
timestamp 1649977179
transform 1 0 16008 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__a21oi_1  _320_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 16468 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a311oi_1  _321_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 14720 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _322_
timestamp 1649977179
transform -1 0 3772 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _323_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 3864 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _324_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 18308 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _325_
timestamp 1649977179
transform 1 0 17756 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _326_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 18400 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _327_
timestamp 1649977179
transform 1 0 18860 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _328_
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _329_
timestamp 1649977179
transform 1 0 22908 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _330_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 28336 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _331_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 27692 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _332_
timestamp 1649977179
transform -1 0 22540 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _333_
timestamp 1649977179
transform 1 0 26680 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _334_
timestamp 1649977179
transform -1 0 22632 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _335_
timestamp 1649977179
transform -1 0 22080 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _336_
timestamp 1649977179
transform -1 0 18216 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _337_
timestamp 1649977179
transform 1 0 11500 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__nor3b_1  _338_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 10580 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _339_
timestamp 1649977179
transform -1 0 10120 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _340_
timestamp 1649977179
transform -1 0 7268 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _341_
timestamp 1649977179
transform -1 0 6808 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _342_
timestamp 1649977179
transform 1 0 26956 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _343_
timestamp 1649977179
transform 1 0 16836 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _344_
timestamp 1649977179
transform 1 0 24656 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__and4bb_1  _345_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9016 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__and4bb_1  _346_
timestamp 1649977179
transform -1 0 12420 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__nor4b_2  _347_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__or4_1  _348_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11868 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _349_
timestamp 1649977179
transform -1 0 19872 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _350_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 25852 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _351_
timestamp 1649977179
transform -1 0 6532 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _352_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _353_
timestamp 1649977179
transform -1 0 10120 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _354_
timestamp 1649977179
transform -1 0 11224 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _355_
timestamp 1649977179
transform 1 0 9936 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _356_
timestamp 1649977179
transform -1 0 22080 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _357_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 22724 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _358_
timestamp 1649977179
transform -1 0 24012 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _359_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 26312 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _360_
timestamp 1649977179
transform -1 0 19412 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _361_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 18584 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _362_
timestamp 1649977179
transform -1 0 19688 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _363_
timestamp 1649977179
transform 1 0 12972 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _364_
timestamp 1649977179
transform -1 0 27048 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _365_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 31096 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _366_
timestamp 1649977179
transform -1 0 33120 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _367_
timestamp 1649977179
transform -1 0 24932 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _368_
timestamp 1649977179
transform -1 0 25116 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _369_
timestamp 1649977179
transform 1 0 20884 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _370_
timestamp 1649977179
transform 1 0 26956 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _371_
timestamp 1649977179
transform 1 0 27232 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _372_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14720 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _373_
timestamp 1649977179
transform -1 0 22448 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _374_
timestamp 1649977179
transform 1 0 22540 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _375_
timestamp 1649977179
transform -1 0 23736 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _376_
timestamp 1649977179
transform -1 0 21712 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _377_
timestamp 1649977179
transform -1 0 16928 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nor4_1  _378_
timestamp 1649977179
transform -1 0 14628 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _379_
timestamp 1649977179
transform -1 0 37168 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _380_
timestamp 1649977179
transform 1 0 29808 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _381_
timestamp 1649977179
transform -1 0 32752 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _382_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 31280 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _383_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 18768 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _384_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2300 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _385_
timestamp 1649977179
transform 1 0 2668 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _386_
timestamp 1649977179
transform 1 0 22172 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _387_
timestamp 1649977179
transform 1 0 18032 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _388_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 18492 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _389_
timestamp 1649977179
transform 1 0 2668 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _390_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 31004 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_2  _391_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 20700 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _392_
timestamp 1649977179
transform -1 0 20424 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _393_
timestamp 1649977179
transform -1 0 15824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _394_
timestamp 1649977179
transform 1 0 20240 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _395_
timestamp 1649977179
transform -1 0 15180 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _396_
timestamp 1649977179
transform 1 0 14628 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _397_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13800 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _398_
timestamp 1649977179
transform 1 0 11960 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _399_
timestamp 1649977179
transform -1 0 27692 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _400_
timestamp 1649977179
transform 1 0 26956 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _401_
timestamp 1649977179
transform -1 0 19596 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _402_
timestamp 1649977179
transform -1 0 18768 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _403_
timestamp 1649977179
transform -1 0 9384 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _404_
timestamp 1649977179
transform 1 0 8924 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _405_
timestamp 1649977179
transform 1 0 8924 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _406_
timestamp 1649977179
transform -1 0 9384 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _407_
timestamp 1649977179
transform 1 0 8924 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _408_
timestamp 1649977179
transform -1 0 25300 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _409_
timestamp 1649977179
transform 1 0 24380 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _410_
timestamp 1649977179
transform -1 0 27048 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _411_
timestamp 1649977179
transform 1 0 20700 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _412_
timestamp 1649977179
transform 1 0 20056 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _413_
timestamp 1649977179
transform -1 0 20976 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _414_
timestamp 1649977179
transform -1 0 7360 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _415_
timestamp 1649977179
transform 1 0 4692 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _416_
timestamp 1649977179
transform -1 0 15088 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _417_
timestamp 1649977179
transform 1 0 14904 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _418_
timestamp 1649977179
transform -1 0 16008 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _419_
timestamp 1649977179
transform -1 0 20240 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _420_
timestamp 1649977179
transform 1 0 19872 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _421_
timestamp 1649977179
transform 1 0 20700 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _422_
timestamp 1649977179
transform -1 0 9384 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _423_
timestamp 1649977179
transform -1 0 32752 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _424_
timestamp 1649977179
transform 1 0 34684 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _425_
timestamp 1649977179
transform -1 0 36064 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _426_
timestamp 1649977179
transform 1 0 19504 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _427_
timestamp 1649977179
transform -1 0 4232 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _428_
timestamp 1649977179
transform -1 0 3312 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _429_
timestamp 1649977179
transform -1 0 4968 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _430_
timestamp 1649977179
transform 1 0 3220 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _431_
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _432_
timestamp 1649977179
transform 1 0 21068 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _433_
timestamp 1649977179
transform 1 0 21804 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _434_
timestamp 1649977179
transform 1 0 20792 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _435_
timestamp 1649977179
transform -1 0 22080 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _436_
timestamp 1649977179
transform -1 0 7360 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _437_
timestamp 1649977179
transform 1 0 6900 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _438_
timestamp 1649977179
transform 1 0 29532 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _439_
timestamp 1649977179
transform 1 0 29992 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _440_
timestamp 1649977179
transform 1 0 22080 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _441_
timestamp 1649977179
transform 1 0 30912 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _442_
timestamp 1649977179
transform 1 0 34592 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _443_
timestamp 1649977179
transform -1 0 35788 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _444_
timestamp 1649977179
transform 1 0 20792 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _445_
timestamp 1649977179
transform -1 0 30820 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _446_
timestamp 1649977179
transform 1 0 23552 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _447_
timestamp 1649977179
transform -1 0 27232 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _448_
timestamp 1649977179
transform 1 0 21068 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _449_
timestamp 1649977179
transform -1 0 24196 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _450_
timestamp 1649977179
transform 1 0 24564 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _451_
timestamp 1649977179
transform 1 0 24748 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _452_
timestamp 1649977179
transform 1 0 3220 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _453_
timestamp 1649977179
transform -1 0 4324 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _454_
timestamp 1649977179
transform 1 0 31464 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _455_
timestamp 1649977179
transform -1 0 33304 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _456_
timestamp 1649977179
transform 1 0 32476 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _457_
timestamp 1649977179
transform 1 0 20976 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _458_
timestamp 1649977179
transform -1 0 22080 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _459_
timestamp 1649977179
transform 1 0 2852 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _460_
timestamp 1649977179
transform -1 0 3312 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _461_
timestamp 1649977179
transform -1 0 17112 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _462_
timestamp 1649977179
transform 1 0 16652 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _463_
timestamp 1649977179
transform 1 0 34960 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _464_
timestamp 1649977179
transform -1 0 36064 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _465_
timestamp 1649977179
transform 1 0 31188 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _466_
timestamp 1649977179
transform -1 0 34960 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _467_
timestamp 1649977179
transform 1 0 24748 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _468_
timestamp 1649977179
transform -1 0 25484 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _469_
timestamp 1649977179
transform 1 0 34500 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _470_
timestamp 1649977179
transform -1 0 36248 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _471_
timestamp 1649977179
transform 1 0 13156 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _472_
timestamp 1649977179
transform -1 0 3128 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _473_
timestamp 1649977179
transform -1 0 2944 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _474_
timestamp 1649977179
transform -1 0 3312 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _475_
timestamp 1649977179
transform -1 0 2944 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _476_
timestamp 1649977179
transform -1 0 3404 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _477_
timestamp 1649977179
transform 1 0 2852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _478_
timestamp 1649977179
transform 1 0 32292 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _479_
timestamp 1649977179
transform -1 0 33948 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _480_
timestamp 1649977179
transform 1 0 15640 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _481_
timestamp 1649977179
transform -1 0 16928 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _482_
timestamp 1649977179
transform 1 0 2668 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _483_
timestamp 1649977179
transform -1 0 3956 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _484_
timestamp 1649977179
transform 1 0 14904 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _485_
timestamp 1649977179
transform -1 0 16008 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _486_
timestamp 1649977179
transform -1 0 31648 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _487_
timestamp 1649977179
transform -1 0 30636 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _488_
timestamp 1649977179
transform -1 0 29992 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _489_
timestamp 1649977179
transform 1 0 28428 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _490_
timestamp 1649977179
transform 1 0 29164 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _491_
timestamp 1649977179
transform 1 0 32568 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _492_
timestamp 1649977179
transform -1 0 33212 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _493_
timestamp 1649977179
transform 1 0 32108 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _494_
timestamp 1649977179
transform -1 0 34040 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _495_
timestamp 1649977179
transform 1 0 28428 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _496_
timestamp 1649977179
transform 1 0 28520 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _497_
timestamp 1649977179
transform 1 0 33120 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _498_
timestamp 1649977179
transform -1 0 34132 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _499_
timestamp 1649977179
transform 1 0 12604 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _500_
timestamp 1649977179
transform 1 0 6348 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _501_
timestamp 1649977179
transform -1 0 6716 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _502_
timestamp 1649977179
transform -1 0 6992 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _503_
timestamp 1649977179
transform 1 0 5520 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _504_
timestamp 1649977179
transform 1 0 5520 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _505_
timestamp 1649977179
transform -1 0 6072 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _506_
timestamp 1649977179
transform 1 0 31188 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _507_
timestamp 1649977179
transform -1 0 34868 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _508_
timestamp 1649977179
transform 1 0 14812 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _509_
timestamp 1649977179
transform -1 0 16468 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _510_
timestamp 1649977179
transform -1 0 20976 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _511_
timestamp 1649977179
transform -1 0 6624 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _512_
timestamp 1649977179
transform 1 0 5888 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _513_
timestamp 1649977179
transform -1 0 12696 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _514_
timestamp 1649977179
transform 1 0 12144 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _515_
timestamp 1649977179
transform 1 0 31004 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _516_
timestamp 1649977179
transform 1 0 29348 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _517_
timestamp 1649977179
transform 1 0 30360 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _518_
timestamp 1649977179
transform -1 0 28796 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _519_
timestamp 1649977179
transform 1 0 28244 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _520_
timestamp 1649977179
transform 1 0 34132 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _521_
timestamp 1649977179
transform -1 0 35236 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _522_
timestamp 1649977179
transform 1 0 30636 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _523_
timestamp 1649977179
transform -1 0 32292 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _524_
timestamp 1649977179
transform 1 0 28704 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _525_
timestamp 1649977179
transform 1 0 29532 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _526_
timestamp 1649977179
transform 1 0 34040 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _527_
timestamp 1649977179
transform -1 0 35328 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _528_
timestamp 1649977179
transform 1 0 14076 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _529_
timestamp 1649977179
transform 1 0 11500 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _530_
timestamp 1649977179
transform -1 0 11960 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _531_
timestamp 1649977179
transform 1 0 7360 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _532_
timestamp 1649977179
transform 1 0 7636 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _533_
timestamp 1649977179
transform -1 0 7268 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _534_
timestamp 1649977179
transform -1 0 7176 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _535_
timestamp 1649977179
transform 1 0 32108 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _536_
timestamp 1649977179
transform -1 0 33580 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _537_
timestamp 1649977179
transform 1 0 15640 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _538_
timestamp 1649977179
transform -1 0 16928 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _539_
timestamp 1649977179
transform -1 0 7268 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _540_
timestamp 1649977179
transform 1 0 6716 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _541_
timestamp 1649977179
transform 1 0 12420 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _542_
timestamp 1649977179
transform 1 0 13248 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _543_
timestamp 1649977179
transform 1 0 31188 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _544_
timestamp 1649977179
transform 1 0 26864 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _545_
timestamp 1649977179
transform -1 0 28336 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _546_
timestamp 1649977179
transform -1 0 26220 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _547_
timestamp 1649977179
transform -1 0 25116 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _548_
timestamp 1649977179
transform 1 0 31188 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _549_
timestamp 1649977179
transform -1 0 31924 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _550_
timestamp 1649977179
transform 1 0 31004 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _551_
timestamp 1649977179
transform -1 0 34960 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _552_
timestamp 1649977179
transform 1 0 28336 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _553_
timestamp 1649977179
transform 1 0 28612 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _554_
timestamp 1649977179
transform 1 0 33028 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _555_
timestamp 1649977179
transform -1 0 34224 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _556_
timestamp 1649977179
transform 1 0 12144 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _557_
timestamp 1649977179
transform 1 0 12788 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _558_
timestamp 1649977179
transform 1 0 9016 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _559_
timestamp 1649977179
transform 1 0 9844 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _560_
timestamp 1649977179
transform -1 0 4232 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _561_
timestamp 1649977179
transform -1 0 3036 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _562_
timestamp 1649977179
transform 1 0 26956 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _563_
timestamp 1649977179
transform 1 0 27140 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _564_
timestamp 1649977179
transform 1 0 19964 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _565_
timestamp 1649977179
transform -1 0 21068 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _566_
timestamp 1649977179
transform -1 0 8372 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _567_
timestamp 1649977179
transform 1 0 7544 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _568_
timestamp 1649977179
transform 1 0 16928 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _569_
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _570_
timestamp 1649977179
transform 1 0 17296 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _571_
timestamp 1649977179
transform 1 0 24380 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _572_
timestamp 1649977179
transform -1 0 25484 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _573_
timestamp 1649977179
transform 1 0 19412 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _574_
timestamp 1649977179
transform -1 0 20148 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _575_
timestamp 1649977179
transform 1 0 24932 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _576_
timestamp 1649977179
transform -1 0 25944 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _577_
timestamp 1649977179
transform 1 0 22448 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _578_
timestamp 1649977179
transform -1 0 24656 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _579_
timestamp 1649977179
transform 1 0 23276 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _580_
timestamp 1649977179
transform -1 0 23920 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _581_
timestamp 1649977179
transform 1 0 32108 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _582_
timestamp 1649977179
transform -1 0 33764 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _583_
timestamp 1649977179
transform -1 0 9476 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _584_
timestamp 1649977179
transform -1 0 13248 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _585_
timestamp 1649977179
transform 1 0 9844 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _586_
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _587_
timestamp 1649977179
transform -1 0 6624 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _588_
timestamp 1649977179
transform -1 0 10212 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _589_
timestamp 1649977179
transform -1 0 7912 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _590_
timestamp 1649977179
transform 1 0 10028 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_1  _591_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 21988 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_2  _592_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 26864 0 1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_1  _593_
timestamp 1649977179
transform 1 0 18032 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_2  _594_
timestamp 1649977179
transform 1 0 21804 0 -1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_1  _595_
timestamp 1649977179
transform 1 0 17480 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _596_
timestamp 1649977179
transform 1 0 27324 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_2  _597_
timestamp 1649977179
transform -1 0 24656 0 -1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_1  _598_
timestamp 1649977179
transform 1 0 10488 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _599_
timestamp 1649977179
transform -1 0 10580 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _600_
timestamp 1649977179
transform -1 0 26864 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_1  _601_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11776 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _602_
timestamp 1649977179
transform 1 0 9108 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _603_
timestamp 1649977179
transform 1 0 12696 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_2  _604_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11500 0 -1 32640
box -38 -48 1602 592
use sky130_fd_sc_hd__dlxtn_1  _605_
timestamp 1649977179
transform 1 0 36432 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _606_
timestamp 1649977179
transform 1 0 27600 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _607_
timestamp 1649977179
transform 1 0 21344 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _608_
timestamp 1649977179
transform 1 0 24472 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_2  _609_
timestamp 1649977179
transform 1 0 35604 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_1  _610_
timestamp 1649977179
transform -1 0 4232 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dfstp_1  _611_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _612_
timestamp 1649977179
transform -1 0 10856 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _613_
timestamp 1649977179
transform 1 0 5428 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _614_
timestamp 1649977179
transform 1 0 10580 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dlxtn_1  _615_
timestamp 1649977179
transform 1 0 3956 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _616_
timestamp 1649977179
transform 1 0 36616 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _617_
timestamp 1649977179
transform 1 0 34776 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _618_
timestamp 1649977179
transform -1 0 3956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _619_
timestamp 1649977179
transform 1 0 21804 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _620_
timestamp 1649977179
transform 1 0 16008 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _621_
timestamp 1649977179
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _622_
timestamp 1649977179
transform -1 0 23920 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _623_
timestamp 1649977179
transform 1 0 25024 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _624_
timestamp 1649977179
transform -1 0 3956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _625_
timestamp 1649977179
transform -1 0 21988 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_2  _626_
timestamp 1649977179
transform 1 0 35604 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_1  _627_
timestamp 1649977179
transform -1 0 3956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _628_
timestamp 1649977179
transform -1 0 9108 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _629_
timestamp 1649977179
transform 1 0 28428 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _630_
timestamp 1649977179
transform 1 0 8096 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _631_
timestamp 1649977179
transform -1 0 20976 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _632_
timestamp 1649977179
transform 1 0 15732 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _633_
timestamp 1649977179
transform 1 0 6348 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _634_
timestamp 1649977179
transform 1 0 29716 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _635_
timestamp 1649977179
transform -1 0 3680 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _636_
timestamp 1649977179
transform -1 0 35052 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _637_
timestamp 1649977179
transform 1 0 35512 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _638_
timestamp 1649977179
transform -1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _639_
timestamp 1649977179
transform 1 0 27692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _640_
timestamp 1649977179
transform 1 0 15548 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _641_
timestamp 1649977179
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _642_
timestamp 1649977179
transform 1 0 17296 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _643_
timestamp 1649977179
transform 1 0 28152 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _644_
timestamp 1649977179
transform -1 0 3312 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _645_
timestamp 1649977179
transform 1 0 29624 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_2  _646_
timestamp 1649977179
transform 1 0 32844 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_1  _647_
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _648_
timestamp 1649977179
transform 1 0 6440 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _649_
timestamp 1649977179
transform 1 0 35696 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _650_
timestamp 1649977179
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _651_
timestamp 1649977179
transform 1 0 5060 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _652_
timestamp 1649977179
transform 1 0 27508 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _653_
timestamp 1649977179
transform 1 0 11684 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _654_
timestamp 1649977179
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _655_
timestamp 1649977179
transform -1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _656_
timestamp 1649977179
transform 1 0 28244 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _657_
timestamp 1649977179
transform -1 0 6348 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _658_
timestamp 1649977179
transform 1 0 29624 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_2  _659_
timestamp 1649977179
transform 1 0 35604 0 1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_1  _660_
timestamp 1649977179
transform -1 0 5888 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _661_
timestamp 1649977179
transform -1 0 12604 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _662_
timestamp 1649977179
transform 1 0 35696 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _663_
timestamp 1649977179
transform 1 0 35328 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _664_
timestamp 1649977179
transform 1 0 7360 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _665_
timestamp 1649977179
transform -1 0 25392 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _666_
timestamp 1649977179
transform -1 0 13340 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _667_
timestamp 1649977179
transform 1 0 35696 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _668_
timestamp 1649977179
transform 1 0 17204 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _669_
timestamp 1649977179
transform 1 0 27968 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _670_
timestamp 1649977179
transform 1 0 6716 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _671_
timestamp 1649977179
transform 1 0 28796 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_2  _672_
timestamp 1649977179
transform -1 0 33304 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_1  _673_
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _674_
timestamp 1649977179
transform -1 0 12880 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _675_
timestamp 1649977179
transform 1 0 34500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _676_
timestamp 1649977179
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _677_
timestamp 1649977179
transform -1 0 9568 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _678_
timestamp 1649977179
transform 1 0 19964 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _679_
timestamp 1649977179
transform 1 0 15824 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _680_
timestamp 1649977179
transform -1 0 27508 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _681_
timestamp 1649977179
transform -1 0 21344 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _682_
timestamp 1649977179
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _683_
timestamp 1649977179
transform -1 0 3312 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _684_
timestamp 1649977179
transform 1 0 25208 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_2  _685_
timestamp 1649977179
transform 1 0 25944 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_1  _686_
timestamp 1649977179
transform 1 0 6440 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _692_
timestamp 1649977179
transform 1 0 7176 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _693_
timestamp 1649977179
transform 1 0 2208 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _694_
timestamp 1649977179
transform 1 0 7820 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _695_
timestamp 1649977179
transform 1 0 2576 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8280 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1649977179
transform 1 0 7820 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1649977179
transform 1 0 7820 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1649977179
transform -1 0 28704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1649977179
transform -1 0 29900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1649977179
transform -1 0 31096 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1649977179
transform -1 0 32384 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform 1 0 33212 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1649977179
transform 1 0 34684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1649977179
transform -1 0 35880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1649977179
transform 1 0 37260 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1649977179
transform 1 0 37904 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1649977179
transform 1 0 37904 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1649977179
transform -1 0 13156 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1649977179
transform -1 0 14352 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1649977179
transform -1 0 15548 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1649977179
transform 1 0 17664 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1649977179
transform -1 0 20332 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1649977179
transform 1 0 21804 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1649977179
transform 1 0 22448 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1649977179
transform 1 0 23644 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1649977179
transform -1 0 4048 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp 1649977179
transform 1 0 9292 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1649977179
transform -1 0 25208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1649977179
transform -1 0 27600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1649977179
transform -1 0 1748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1649977179
transform -1 0 1748 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1649977179
transform -1 0 1748 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1649977179
transform -1 0 1748 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1649977179
transform -1 0 1748 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1649977179
transform -1 0 1748 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1649977179
transform -1 0 1748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1649977179
transform -1 0 1748 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1649977179
transform -1 0 1748 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1649977179
transform -1 0 1748 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1649977179
transform -1 0 1748 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 1649977179
transform -1 0 1748 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 1649977179
transform -1 0 1748 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 1649977179
transform -1 0 1748 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp 1649977179
transform -1 0 1748 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp 1649977179
transform -1 0 1748 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 1649977179
transform -1 0 9660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1649977179
transform -1 0 12052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 1649977179
transform -1 0 2484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp 1649977179
transform -1 0 4876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp 1649977179
transform -1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp 1649977179
transform -1 0 7268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp 1649977179
transform -1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 1649977179
transform -1 0 1748 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1649977179
transform -1 0 1748 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 1649977179
transform -1 0 1748 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1649977179
transform -1 0 1748 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 1649977179
transform -1 0 1748 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1649977179
transform -1 0 1748 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1649977179
transform -1 0 1748 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1649977179
transform -1 0 1748 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  pixel_82 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 1656 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_83
timestamp 1649977179
transform -1 0 20332 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_84
timestamp 1649977179
transform -1 0 26036 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_85
timestamp 1649977179
transform -1 0 32384 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_86
timestamp 1649977179
transform -1 0 37536 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater56
timestamp 1649977179
transform -1 0 24840 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater57
timestamp 1649977179
transform 1 0 11500 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  repeater58
timestamp 1649977179
transform -1 0 8096 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater59
timestamp 1649977179
transform -1 0 27968 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater60
timestamp 1649977179
transform 1 0 20056 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater61
timestamp 1649977179
transform -1 0 35972 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater62
timestamp 1649977179
transform 1 0 24380 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater63
timestamp 1649977179
transform 1 0 15364 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater64
timestamp 1649977179
transform -1 0 11868 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater65
timestamp 1649977179
transform -1 0 33856 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater66
timestamp 1649977179
transform -1 0 6440 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  repeater67
timestamp 1649977179
transform 1 0 30912 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  repeater68
timestamp 1649977179
transform -1 0 19320 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater69
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  repeater70
timestamp 1649977179
transform 1 0 19504 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  repeater71 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 28060 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  repeater72
timestamp 1649977179
transform 1 0 31188 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  repeater73
timestamp 1649977179
transform -1 0 32200 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  repeater74
timestamp 1649977179
transform 1 0 24748 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  repeater75
timestamp 1649977179
transform -1 0 6716 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  repeater76
timestamp 1649977179
transform 1 0 6900 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  repeater77
timestamp 1649977179
transform -1 0 25576 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater78
timestamp 1649977179
transform -1 0 26220 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  repeater79
timestamp 1649977179
transform -1 0 20332 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater80
timestamp 1649977179
transform 1 0 19320 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater81
timestamp 1649977179
transform -1 0 11776 0 1 15232
box -38 -48 406 592
<< labels >>
flabel metal2 s 28354 0 28410 800 0 FreeSans 224 90 0 0 adj_max_clk[0]
port 0 nsew signal input
flabel metal2 s 29550 0 29606 800 0 FreeSans 224 90 0 0 adj_max_clk[1]
port 1 nsew signal input
flabel metal2 s 30746 0 30802 800 0 FreeSans 224 90 0 0 adj_max_clk[2]
port 2 nsew signal input
flabel metal2 s 31942 0 31998 800 0 FreeSans 224 90 0 0 adj_max_clk[3]
port 3 nsew signal input
flabel metal2 s 33138 0 33194 800 0 FreeSans 224 90 0 0 adj_max_clk[4]
port 4 nsew signal input
flabel metal2 s 34334 0 34390 800 0 FreeSans 224 90 0 0 adj_max_clk[5]
port 5 nsew signal input
flabel metal2 s 35530 0 35586 800 0 FreeSans 224 90 0 0 adj_max_clk[6]
port 6 nsew signal input
flabel metal2 s 36726 0 36782 800 0 FreeSans 224 90 0 0 adj_max_clk[7]
port 7 nsew signal input
flabel metal2 s 37922 0 37978 800 0 FreeSans 224 90 0 0 adj_max_clk[8]
port 8 nsew signal input
flabel metal2 s 39118 0 39174 800 0 FreeSans 224 90 0 0 adj_max_clk[9]
port 9 nsew signal input
flabel metal2 s 24766 0 24822 800 0 FreeSans 224 90 0 0 adj_timer_en
port 10 nsew signal tristate
flabel metal2 s 25962 0 26018 800 0 FreeSans 224 90 0 0 adj_timer_m_i
port 11 nsew signal input
flabel metal2 s 27158 0 27214 800 0 FreeSans 224 90 0 0 adj_timer_max
port 12 nsew signal tristate
flabel metal2 s 2870 35200 2926 36000 0 FreeSans 224 90 0 0 clk
port 13 nsew signal input
flabel metal2 s 14278 35200 14334 36000 0 FreeSans 224 90 0 0 data_in
port 14 nsew signal input
flabel metal3 s 0 1640 800 1760 0 FreeSans 480 0 0 0 data_out[0]
port 15 nsew signal tristate
flabel metal3 s 0 15240 800 15360 0 FreeSans 480 0 0 0 data_out[10]
port 16 nsew signal tristate
flabel metal3 s 0 16600 800 16720 0 FreeSans 480 0 0 0 data_out[11]
port 17 nsew signal tristate
flabel metal3 s 0 17960 800 18080 0 FreeSans 480 0 0 0 data_out[12]
port 18 nsew signal tristate
flabel metal3 s 0 19320 800 19440 0 FreeSans 480 0 0 0 data_out[13]
port 19 nsew signal tristate
flabel metal3 s 0 20680 800 20800 0 FreeSans 480 0 0 0 data_out[14]
port 20 nsew signal tristate
flabel metal3 s 0 22040 800 22160 0 FreeSans 480 0 0 0 data_out[15]
port 21 nsew signal tristate
flabel metal3 s 0 3000 800 3120 0 FreeSans 480 0 0 0 data_out[1]
port 22 nsew signal tristate
flabel metal3 s 0 4360 800 4480 0 FreeSans 480 0 0 0 data_out[2]
port 23 nsew signal tristate
flabel metal3 s 0 5720 800 5840 0 FreeSans 480 0 0 0 data_out[3]
port 24 nsew signal tristate
flabel metal3 s 0 7080 800 7200 0 FreeSans 480 0 0 0 data_out[4]
port 25 nsew signal tristate
flabel metal3 s 0 8440 800 8560 0 FreeSans 480 0 0 0 data_out[5]
port 26 nsew signal tristate
flabel metal3 s 0 9800 800 9920 0 FreeSans 480 0 0 0 data_out[6]
port 27 nsew signal tristate
flabel metal3 s 0 11160 800 11280 0 FreeSans 480 0 0 0 data_out[7]
port 28 nsew signal tristate
flabel metal3 s 0 12520 800 12640 0 FreeSans 480 0 0 0 data_out[8]
port 29 nsew signal tristate
flabel metal3 s 0 13880 800 14000 0 FreeSans 480 0 0 0 data_out[9]
port 30 nsew signal tristate
flabel metal2 s 19982 35200 20038 36000 0 FreeSans 224 90 0 0 data_sel[0]
port 31 nsew signal tristate
flabel metal2 s 25686 35200 25742 36000 0 FreeSans 224 90 0 0 data_sel[1]
port 32 nsew signal tristate
flabel metal2 s 31390 35200 31446 36000 0 FreeSans 224 90 0 0 data_sel[2]
port 33 nsew signal tristate
flabel metal2 s 37094 35200 37150 36000 0 FreeSans 224 90 0 0 data_sel[3]
port 34 nsew signal tristate
flabel metal3 s 0 34280 800 34400 0 FreeSans 480 0 0 0 kernel_done_o
port 35 nsew signal tristate
flabel metal2 s 12806 0 12862 800 0 FreeSans 224 90 0 0 loc_max_clk[0]
port 36 nsew signal input
flabel metal2 s 14002 0 14058 800 0 FreeSans 224 90 0 0 loc_max_clk[1]
port 37 nsew signal input
flabel metal2 s 15198 0 15254 800 0 FreeSans 224 90 0 0 loc_max_clk[2]
port 38 nsew signal input
flabel metal2 s 16394 0 16450 800 0 FreeSans 224 90 0 0 loc_max_clk[3]
port 39 nsew signal input
flabel metal2 s 17590 0 17646 800 0 FreeSans 224 90 0 0 loc_max_clk[4]
port 40 nsew signal input
flabel metal2 s 18786 0 18842 800 0 FreeSans 224 90 0 0 loc_max_clk[5]
port 41 nsew signal input
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 loc_max_clk[6]
port 42 nsew signal input
flabel metal2 s 21178 0 21234 800 0 FreeSans 224 90 0 0 loc_max_clk[7]
port 43 nsew signal input
flabel metal2 s 22374 0 22430 800 0 FreeSans 224 90 0 0 loc_max_clk[8]
port 44 nsew signal input
flabel metal2 s 23570 0 23626 800 0 FreeSans 224 90 0 0 loc_max_clk[9]
port 45 nsew signal input
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 loc_timer_en
port 46 nsew signal tristate
flabel metal2 s 10414 0 10470 800 0 FreeSans 224 90 0 0 loc_timer_m_i
port 47 nsew signal input
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 loc_timer_max
port 48 nsew signal tristate
flabel metal2 s 846 0 902 800 0 FreeSans 224 90 0 0 pxl_done_i
port 49 nsew signal input
flabel metal2 s 2042 0 2098 800 0 FreeSans 224 90 0 0 pxl_done_o
port 50 nsew signal tristate
flabel metal2 s 4434 0 4490 800 0 FreeSans 224 90 0 0 pxl_q[0]
port 51 nsew signal tristate
flabel metal2 s 5630 0 5686 800 0 FreeSans 224 90 0 0 pxl_q[1]
port 52 nsew signal tristate
flabel metal2 s 6826 0 6882 800 0 FreeSans 224 90 0 0 pxl_q[2]
port 53 nsew signal tristate
flabel metal2 s 8022 0 8078 800 0 FreeSans 224 90 0 0 pxl_q[3]
port 54 nsew signal tristate
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 pxl_start_i
port 55 nsew signal input
flabel metal2 s 8574 35200 8630 36000 0 FreeSans 224 90 0 0 reset
port 56 nsew signal input
flabel metal3 s 0 23400 800 23520 0 FreeSans 480 0 0 0 s1
port 57 nsew signal tristate
flabel metal3 s 0 24760 800 24880 0 FreeSans 480 0 0 0 s1_inv
port 58 nsew signal tristate
flabel metal3 s 0 26120 800 26240 0 FreeSans 480 0 0 0 s2
port 59 nsew signal tristate
flabel metal3 s 0 27480 800 27600 0 FreeSans 480 0 0 0 s2_inv
port 60 nsew signal tristate
flabel metal3 s 0 28840 800 28960 0 FreeSans 480 0 0 0 s_p1
port 61 nsew signal tristate
flabel metal3 s 0 30200 800 30320 0 FreeSans 480 0 0 0 s_p2
port 62 nsew signal tristate
flabel metal3 s 0 31560 800 31680 0 FreeSans 480 0 0 0 v_b0
port 63 nsew signal tristate
flabel metal3 s 0 32920 800 33040 0 FreeSans 480 0 0 0 v_b1
port 64 nsew signal tristate
flabel metal4 s 5668 2128 5988 33776 0 FreeSans 1920 90 0 0 vccd1
port 65 nsew power bidirectional
flabel metal4 s 15116 2128 15436 33776 0 FreeSans 1920 90 0 0 vccd1
port 65 nsew power bidirectional
flabel metal4 s 24564 2128 24884 33776 0 FreeSans 1920 90 0 0 vccd1
port 65 nsew power bidirectional
flabel metal4 s 34012 2128 34332 33776 0 FreeSans 1920 90 0 0 vccd1
port 65 nsew power bidirectional
flabel metal4 s 10392 2128 10712 33776 0 FreeSans 1920 90 0 0 vssd1
port 66 nsew ground bidirectional
flabel metal4 s 19840 2128 20160 33776 0 FreeSans 1920 90 0 0 vssd1
port 66 nsew ground bidirectional
flabel metal4 s 29288 2128 29608 33776 0 FreeSans 1920 90 0 0 vssd1
port 66 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 40000 36000
<< end >>
