** sch_path: /home/icarosix/asic/analog/MixPix/analog/xschem/Diode_Dtemp_tb.sch
**.subckt Diode_Dtemp_tb
.model 1N914 D(level=3 Is=252f N=1.752 Rs=.568 ISR=0 NR=1 JSW =0 IKR = 0 IK = 0 Cjo=4p M=.4 tt=20n )
V2 net1 GND 0
V1 net2 GND 0
V3 net3 GND 0
D1 net1 net3 1N914 area=1 dtemp=10
D2 net1 net2 1N914 area=1
**** begin user architecture code
.control
set hcopydevtype = svg
set nolegend
set color0=white
set color1=black
set color2=blue
set color3=red
save all
dc V2 -10 0 100u
plot I(V1) I(V3)
hardcopy Inverse.svg I(V1) I(V3)
.endc
*.lib /home/icarosix/asic/pdks/sky130A/libs.tech/ngspice/models/sky130.lib.spice tt
*.lib /home/icarosix/asic/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.option wnflag=1
**** end user architecture code
**.ends
.GLOBAL GND
**** begin user architecture code
?
**** end user architecture code
.end
