magic
tech sky130B
magscale 1 2
timestamp 1667007431
<< obsli1 >>
rect 121104 82159 188816 257681
<< obsm1 >>
rect 14 2864 582714 703044
<< metal2 >>
rect 634 703520 746 704960
rect 4498 703520 4610 704960
rect 8362 703520 8474 704960
rect 12226 703520 12338 704960
rect 16090 703520 16202 704960
rect 19954 703520 20066 704960
rect 23818 703520 23930 704960
rect 27682 703520 27794 704960
rect 31546 703520 31658 704960
rect 34766 703520 34878 704960
rect 38630 703520 38742 704960
rect 42494 703520 42606 704960
rect 46358 703520 46470 704960
rect 50222 703520 50334 704960
rect 54086 703520 54198 704960
rect 57950 703520 58062 704960
rect 61814 703520 61926 704960
rect 65678 703520 65790 704960
rect 68898 703520 69010 704960
rect 72762 703520 72874 704960
rect 76626 703520 76738 704960
rect 80490 703520 80602 704960
rect 84354 703520 84466 704960
rect 88218 703520 88330 704960
rect 92082 703520 92194 704960
rect 95946 703520 96058 704960
rect 99810 703520 99922 704960
rect 103674 703520 103786 704960
rect 106894 703520 107006 704960
rect 110758 703520 110870 704960
rect 114622 703520 114734 704960
rect 118486 703520 118598 704960
rect 122350 703520 122462 704960
rect 126214 703520 126326 704960
rect 130078 703520 130190 704960
rect 133942 703520 134054 704960
rect 137806 703520 137918 704960
rect 141670 703520 141782 704960
rect 144890 703520 145002 704960
rect 148754 703520 148866 704960
rect 152618 703520 152730 704960
rect 156482 703520 156594 704960
rect 160346 703520 160458 704960
rect 164210 703520 164322 704960
rect 168074 703520 168186 704960
rect 171938 703520 172050 704960
rect 175802 703520 175914 704960
rect 179022 703520 179134 704960
rect 182886 703520 182998 704960
rect 186750 703520 186862 704960
rect 190614 703520 190726 704960
rect 194478 703520 194590 704960
rect 198342 703520 198454 704960
rect 202206 703520 202318 704960
rect 206070 703520 206182 704960
rect 209934 703520 210046 704960
rect 213798 703520 213910 704960
rect 217018 703520 217130 704960
rect 220882 703520 220994 704960
rect 224746 703520 224858 704960
rect 228610 703520 228722 704960
rect 232474 703520 232586 704960
rect 236338 703520 236450 704960
rect 240202 703520 240314 704960
rect 244066 703520 244178 704960
rect 247930 703520 248042 704960
rect 251794 703520 251906 704960
rect 255014 703520 255126 704960
rect 258878 703520 258990 704960
rect 262742 703520 262854 704960
rect 266606 703520 266718 704960
rect 270470 703520 270582 704960
rect 274334 703520 274446 704960
rect 278198 703520 278310 704960
rect 282062 703520 282174 704960
rect 285926 703520 286038 704960
rect 289146 703520 289258 704960
rect 293010 703520 293122 704960
rect 296874 703520 296986 704960
rect 300738 703520 300850 704960
rect 304602 703520 304714 704960
rect 308466 703520 308578 704960
rect 312330 703520 312442 704960
rect 316194 703520 316306 704960
rect 320058 703520 320170 704960
rect 323922 703520 324034 704960
rect 327142 703520 327254 704960
rect 331006 703520 331118 704960
rect 334870 703520 334982 704960
rect 338734 703520 338846 704960
rect 342598 703520 342710 704960
rect 346462 703520 346574 704960
rect 350326 703520 350438 704960
rect 354190 703520 354302 704960
rect 358054 703520 358166 704960
rect 361918 703520 362030 704960
rect 365138 703520 365250 704960
rect 369002 703520 369114 704960
rect 372866 703520 372978 704960
rect 376730 703520 376842 704960
rect 380594 703520 380706 704960
rect 384458 703520 384570 704960
rect 388322 703520 388434 704960
rect 392186 703520 392298 704960
rect 396050 703520 396162 704960
rect 399914 703520 400026 704960
rect 403134 703520 403246 704960
rect 406998 703520 407110 704960
rect 410862 703520 410974 704960
rect 414726 703520 414838 704960
rect 418590 703520 418702 704960
rect 422454 703520 422566 704960
rect 426318 703520 426430 704960
rect 430182 703520 430294 704960
rect 434046 703520 434158 704960
rect 437266 703520 437378 704960
rect 441130 703520 441242 704960
rect 444994 703520 445106 704960
rect 448858 703520 448970 704960
rect 452722 703520 452834 704960
rect 456586 703520 456698 704960
rect 460450 703520 460562 704960
rect 464314 703520 464426 704960
rect 468178 703520 468290 704960
rect 472042 703520 472154 704960
rect 475262 703520 475374 704960
rect 479126 703520 479238 704960
rect 482990 703520 483102 704960
rect 486854 703520 486966 704960
rect 490718 703520 490830 704960
rect 494582 703520 494694 704960
rect 498446 703520 498558 704960
rect 502310 703520 502422 704960
rect 506174 703520 506286 704960
rect 510038 703520 510150 704960
rect 513258 703520 513370 704960
rect 517122 703520 517234 704960
rect 520986 703520 521098 704960
rect 524850 703520 524962 704960
rect 528714 703520 528826 704960
rect 532578 703520 532690 704960
rect 536442 703520 536554 704960
rect 540306 703520 540418 704960
rect 544170 703520 544282 704960
rect 547390 703520 547502 704960
rect 551254 703520 551366 704960
rect 555118 703520 555230 704960
rect 558982 703520 559094 704960
rect 562846 703520 562958 704960
rect 566710 703520 566822 704960
rect 570574 703520 570686 704960
rect 574438 703520 574550 704960
rect 578302 703520 578414 704960
rect 582166 703520 582278 704960
rect -10 -960 102 480
rect 3210 -960 3322 480
rect 7074 -960 7186 480
rect 10938 -960 11050 480
rect 14802 -960 14914 480
rect 18666 -960 18778 480
rect 22530 -960 22642 480
rect 26394 -960 26506 480
rect 30258 -960 30370 480
rect 34122 -960 34234 480
rect 37342 -960 37454 480
rect 41206 -960 41318 480
rect 45070 -960 45182 480
rect 48934 -960 49046 480
rect 52798 -960 52910 480
rect 56662 -960 56774 480
rect 60526 -960 60638 480
rect 64390 -960 64502 480
rect 68254 -960 68366 480
rect 72118 -960 72230 480
rect 75338 -960 75450 480
rect 79202 -960 79314 480
rect 83066 -960 83178 480
rect 86930 -960 87042 480
rect 90794 -960 90906 480
rect 94658 -960 94770 480
rect 98522 -960 98634 480
rect 102386 -960 102498 480
rect 106250 -960 106362 480
rect 110114 -960 110226 480
rect 113334 -960 113446 480
rect 117198 -960 117310 480
rect 121062 -960 121174 480
rect 124926 -960 125038 480
rect 128790 -960 128902 480
rect 132654 -960 132766 480
rect 136518 -960 136630 480
rect 140382 -960 140494 480
rect 144246 -960 144358 480
rect 147466 -960 147578 480
rect 151330 -960 151442 480
rect 155194 -960 155306 480
rect 159058 -960 159170 480
rect 162922 -960 163034 480
rect 166786 -960 166898 480
rect 170650 -960 170762 480
rect 174514 -960 174626 480
rect 178378 -960 178490 480
rect 182242 -960 182354 480
rect 185462 -960 185574 480
rect 189326 -960 189438 480
rect 193190 -960 193302 480
rect 197054 -960 197166 480
rect 200918 -960 201030 480
rect 204782 -960 204894 480
rect 208646 -960 208758 480
rect 212510 -960 212622 480
rect 216374 -960 216486 480
rect 220238 -960 220350 480
rect 223458 -960 223570 480
rect 227322 -960 227434 480
rect 231186 -960 231298 480
rect 235050 -960 235162 480
rect 238914 -960 239026 480
rect 242778 -960 242890 480
rect 246642 -960 246754 480
rect 250506 -960 250618 480
rect 254370 -960 254482 480
rect 257590 -960 257702 480
rect 261454 -960 261566 480
rect 265318 -960 265430 480
rect 269182 -960 269294 480
rect 273046 -960 273158 480
rect 276910 -960 277022 480
rect 280774 -960 280886 480
rect 284638 -960 284750 480
rect 288502 -960 288614 480
rect 292366 -960 292478 480
rect 295586 -960 295698 480
rect 299450 -960 299562 480
rect 303314 -960 303426 480
rect 307178 -960 307290 480
rect 311042 -960 311154 480
rect 314906 -960 315018 480
rect 318770 -960 318882 480
rect 322634 -960 322746 480
rect 326498 -960 326610 480
rect 330362 -960 330474 480
rect 333582 -960 333694 480
rect 337446 -960 337558 480
rect 341310 -960 341422 480
rect 345174 -960 345286 480
rect 349038 -960 349150 480
rect 352902 -960 353014 480
rect 356766 -960 356878 480
rect 360630 -960 360742 480
rect 364494 -960 364606 480
rect 367714 -960 367826 480
rect 371578 -960 371690 480
rect 375442 -960 375554 480
rect 379306 -960 379418 480
rect 383170 -960 383282 480
rect 387034 -960 387146 480
rect 390898 -960 391010 480
rect 394762 -960 394874 480
rect 398626 -960 398738 480
rect 402490 -960 402602 480
rect 405710 -960 405822 480
rect 409574 -960 409686 480
rect 413438 -960 413550 480
rect 417302 -960 417414 480
rect 421166 -960 421278 480
rect 425030 -960 425142 480
rect 428894 -960 429006 480
rect 432758 -960 432870 480
rect 436622 -960 436734 480
rect 440486 -960 440598 480
rect 443706 -960 443818 480
rect 447570 -960 447682 480
rect 451434 -960 451546 480
rect 455298 -960 455410 480
rect 459162 -960 459274 480
rect 463026 -960 463138 480
rect 466890 -960 467002 480
rect 470754 -960 470866 480
rect 474618 -960 474730 480
rect 477838 -960 477950 480
rect 481702 -960 481814 480
rect 485566 -960 485678 480
rect 489430 -960 489542 480
rect 493294 -960 493406 480
rect 497158 -960 497270 480
rect 501022 -960 501134 480
rect 504886 -960 504998 480
rect 508750 -960 508862 480
rect 512614 -960 512726 480
rect 515834 -960 515946 480
rect 519698 -960 519810 480
rect 523562 -960 523674 480
rect 527426 -960 527538 480
rect 531290 -960 531402 480
rect 535154 -960 535266 480
rect 539018 -960 539130 480
rect 542882 -960 542994 480
rect 546746 -960 546858 480
rect 550610 -960 550722 480
rect 553830 -960 553942 480
rect 557694 -960 557806 480
rect 561558 -960 561670 480
rect 565422 -960 565534 480
rect 569286 -960 569398 480
rect 573150 -960 573262 480
rect 577014 -960 577126 480
rect 580878 -960 580990 480
<< obsm2 >>
rect 20 703464 578 703610
rect 802 703464 4442 703610
rect 4666 703464 8306 703610
rect 8530 703464 12170 703610
rect 12394 703464 16034 703610
rect 16258 703464 19898 703610
rect 20122 703464 23762 703610
rect 23986 703464 27626 703610
rect 27850 703464 31490 703610
rect 31714 703464 34710 703610
rect 34934 703464 38574 703610
rect 38798 703464 42438 703610
rect 42662 703464 46302 703610
rect 46526 703464 50166 703610
rect 50390 703464 54030 703610
rect 54254 703464 57894 703610
rect 58118 703464 61758 703610
rect 61982 703464 65622 703610
rect 65846 703464 68842 703610
rect 69066 703464 72706 703610
rect 72930 703464 76570 703610
rect 76794 703464 80434 703610
rect 80658 703464 84298 703610
rect 84522 703464 88162 703610
rect 88386 703464 92026 703610
rect 92250 703464 95890 703610
rect 96114 703464 99754 703610
rect 99978 703464 103618 703610
rect 103842 703464 106838 703610
rect 107062 703464 110702 703610
rect 110926 703464 114566 703610
rect 114790 703464 118430 703610
rect 118654 703464 122294 703610
rect 122518 703464 126158 703610
rect 126382 703464 130022 703610
rect 130246 703464 133886 703610
rect 134110 703464 137750 703610
rect 137974 703464 141614 703610
rect 141838 703464 144834 703610
rect 145058 703464 148698 703610
rect 148922 703464 152562 703610
rect 152786 703464 156426 703610
rect 156650 703464 160290 703610
rect 160514 703464 164154 703610
rect 164378 703464 168018 703610
rect 168242 703464 171882 703610
rect 172106 703464 175746 703610
rect 175970 703464 178966 703610
rect 179190 703464 182830 703610
rect 183054 703464 186694 703610
rect 186918 703464 190558 703610
rect 190782 703464 194422 703610
rect 194646 703464 198286 703610
rect 198510 703464 202150 703610
rect 202374 703464 206014 703610
rect 206238 703464 209878 703610
rect 210102 703464 213742 703610
rect 213966 703464 216962 703610
rect 217186 703464 220826 703610
rect 221050 703464 224690 703610
rect 224914 703464 228554 703610
rect 228778 703464 232418 703610
rect 232642 703464 236282 703610
rect 236506 703464 240146 703610
rect 240370 703464 244010 703610
rect 244234 703464 247874 703610
rect 248098 703464 251738 703610
rect 251962 703464 254958 703610
rect 255182 703464 258822 703610
rect 259046 703464 262686 703610
rect 262910 703464 266550 703610
rect 266774 703464 270414 703610
rect 270638 703464 274278 703610
rect 274502 703464 278142 703610
rect 278366 703464 282006 703610
rect 282230 703464 285870 703610
rect 286094 703464 289090 703610
rect 289314 703464 292954 703610
rect 293178 703464 296818 703610
rect 297042 703464 300682 703610
rect 300906 703464 304546 703610
rect 304770 703464 308410 703610
rect 308634 703464 312274 703610
rect 312498 703464 316138 703610
rect 316362 703464 320002 703610
rect 320226 703464 323866 703610
rect 324090 703464 327086 703610
rect 327310 703464 330950 703610
rect 331174 703464 334814 703610
rect 335038 703464 338678 703610
rect 338902 703464 342542 703610
rect 342766 703464 346406 703610
rect 346630 703464 350270 703610
rect 350494 703464 354134 703610
rect 354358 703464 357998 703610
rect 358222 703464 361862 703610
rect 362086 703464 365082 703610
rect 365306 703464 368946 703610
rect 369170 703464 372810 703610
rect 373034 703464 376674 703610
rect 376898 703464 380538 703610
rect 380762 703464 384402 703610
rect 384626 703464 388266 703610
rect 388490 703464 392130 703610
rect 392354 703464 395994 703610
rect 396218 703464 399858 703610
rect 400082 703464 403078 703610
rect 403302 703464 406942 703610
rect 407166 703464 410806 703610
rect 411030 703464 414670 703610
rect 414894 703464 418534 703610
rect 418758 703464 422398 703610
rect 422622 703464 426262 703610
rect 426486 703464 430126 703610
rect 430350 703464 433990 703610
rect 434214 703464 437210 703610
rect 437434 703464 441074 703610
rect 441298 703464 444938 703610
rect 445162 703464 448802 703610
rect 449026 703464 452666 703610
rect 452890 703464 456530 703610
rect 456754 703464 460394 703610
rect 460618 703464 464258 703610
rect 464482 703464 468122 703610
rect 468346 703464 471986 703610
rect 472210 703464 475206 703610
rect 475430 703464 479070 703610
rect 479294 703464 482934 703610
rect 483158 703464 486798 703610
rect 487022 703464 490662 703610
rect 490886 703464 494526 703610
rect 494750 703464 498390 703610
rect 498614 703464 502254 703610
rect 502478 703464 506118 703610
rect 506342 703464 509982 703610
rect 510206 703464 513202 703610
rect 513426 703464 517066 703610
rect 517290 703464 520930 703610
rect 521154 703464 524794 703610
rect 525018 703464 528658 703610
rect 528882 703464 532522 703610
rect 532746 703464 536386 703610
rect 536610 703464 540250 703610
rect 540474 703464 544114 703610
rect 544338 703464 547334 703610
rect 547558 703464 551198 703610
rect 551422 703464 555062 703610
rect 555286 703464 558926 703610
rect 559150 703464 562790 703610
rect 563014 703464 566654 703610
rect 566878 703464 570518 703610
rect 570742 703464 574382 703610
rect 574606 703464 578246 703610
rect 578470 703464 582110 703610
rect 582334 703464 582894 703610
rect 20 536 582894 703464
rect 158 326 3154 536
rect 3378 326 7018 536
rect 7242 326 10882 536
rect 11106 326 14746 536
rect 14970 326 18610 536
rect 18834 326 22474 536
rect 22698 326 26338 536
rect 26562 326 30202 536
rect 30426 326 34066 536
rect 34290 326 37286 536
rect 37510 326 41150 536
rect 41374 326 45014 536
rect 45238 326 48878 536
rect 49102 326 52742 536
rect 52966 326 56606 536
rect 56830 326 60470 536
rect 60694 326 64334 536
rect 64558 326 68198 536
rect 68422 326 72062 536
rect 72286 326 75282 536
rect 75506 326 79146 536
rect 79370 326 83010 536
rect 83234 326 86874 536
rect 87098 326 90738 536
rect 90962 326 94602 536
rect 94826 326 98466 536
rect 98690 326 102330 536
rect 102554 326 106194 536
rect 106418 326 110058 536
rect 110282 326 113278 536
rect 113502 326 117142 536
rect 117366 326 121006 536
rect 121230 326 124870 536
rect 125094 326 128734 536
rect 128958 326 132598 536
rect 132822 326 136462 536
rect 136686 326 140326 536
rect 140550 326 144190 536
rect 144414 326 147410 536
rect 147634 326 151274 536
rect 151498 326 155138 536
rect 155362 326 159002 536
rect 159226 326 162866 536
rect 163090 326 166730 536
rect 166954 326 170594 536
rect 170818 326 174458 536
rect 174682 326 178322 536
rect 178546 326 182186 536
rect 182410 326 185406 536
rect 185630 326 189270 536
rect 189494 326 193134 536
rect 193358 326 196998 536
rect 197222 326 200862 536
rect 201086 326 204726 536
rect 204950 326 208590 536
rect 208814 326 212454 536
rect 212678 326 216318 536
rect 216542 326 220182 536
rect 220406 326 223402 536
rect 223626 326 227266 536
rect 227490 326 231130 536
rect 231354 326 234994 536
rect 235218 326 238858 536
rect 239082 326 242722 536
rect 242946 326 246586 536
rect 246810 326 250450 536
rect 250674 326 254314 536
rect 254538 326 257534 536
rect 257758 326 261398 536
rect 261622 326 265262 536
rect 265486 326 269126 536
rect 269350 326 272990 536
rect 273214 326 276854 536
rect 277078 326 280718 536
rect 280942 326 284582 536
rect 284806 326 288446 536
rect 288670 326 292310 536
rect 292534 326 295530 536
rect 295754 326 299394 536
rect 299618 326 303258 536
rect 303482 326 307122 536
rect 307346 326 310986 536
rect 311210 326 314850 536
rect 315074 326 318714 536
rect 318938 326 322578 536
rect 322802 326 326442 536
rect 326666 326 330306 536
rect 330530 326 333526 536
rect 333750 326 337390 536
rect 337614 326 341254 536
rect 341478 326 345118 536
rect 345342 326 348982 536
rect 349206 326 352846 536
rect 353070 326 356710 536
rect 356934 326 360574 536
rect 360798 326 364438 536
rect 364662 326 367658 536
rect 367882 326 371522 536
rect 371746 326 375386 536
rect 375610 326 379250 536
rect 379474 326 383114 536
rect 383338 326 386978 536
rect 387202 326 390842 536
rect 391066 326 394706 536
rect 394930 326 398570 536
rect 398794 326 402434 536
rect 402658 326 405654 536
rect 405878 326 409518 536
rect 409742 326 413382 536
rect 413606 326 417246 536
rect 417470 326 421110 536
rect 421334 326 424974 536
rect 425198 326 428838 536
rect 429062 326 432702 536
rect 432926 326 436566 536
rect 436790 326 440430 536
rect 440654 326 443650 536
rect 443874 326 447514 536
rect 447738 326 451378 536
rect 451602 326 455242 536
rect 455466 326 459106 536
rect 459330 326 462970 536
rect 463194 326 466834 536
rect 467058 326 470698 536
rect 470922 326 474562 536
rect 474786 326 477782 536
rect 478006 326 481646 536
rect 481870 326 485510 536
rect 485734 326 489374 536
rect 489598 326 493238 536
rect 493462 326 497102 536
rect 497326 326 500966 536
rect 501190 326 504830 536
rect 505054 326 508694 536
rect 508918 326 512558 536
rect 512782 326 515778 536
rect 516002 326 519642 536
rect 519866 326 523506 536
rect 523730 326 527370 536
rect 527594 326 531234 536
rect 531458 326 535098 536
rect 535322 326 538962 536
rect 539186 326 542826 536
rect 543050 326 546690 536
rect 546914 326 550554 536
rect 550778 326 553774 536
rect 553998 326 557638 536
rect 557862 326 561502 536
rect 561726 326 565366 536
rect 565590 326 569230 536
rect 569454 326 573094 536
rect 573318 326 576958 536
rect 577182 326 580822 536
rect 581046 326 582894 536
<< metal3 >>
rect 583520 702388 584960 702628
rect -960 701028 480 701268
rect 583520 698308 584960 698548
rect -960 697628 480 697868
rect 583520 694228 584960 694468
rect -960 693548 480 693788
rect 583520 690148 584960 690388
rect -960 689468 480 689708
rect 583520 686068 584960 686308
rect -960 685388 480 685628
rect 583520 681988 584960 682228
rect -960 681308 480 681548
rect 583520 677908 584960 678148
rect -960 677228 480 677468
rect 583520 673828 584960 674068
rect -960 673148 480 673388
rect 583520 669748 584960 669988
rect -960 669068 480 669308
rect 583520 665668 584960 665908
rect -960 664988 480 665228
rect 583520 662268 584960 662508
rect -960 660908 480 661148
rect 583520 658188 584960 658428
rect -960 657508 480 657748
rect 583520 654108 584960 654348
rect -960 653428 480 653668
rect 583520 650028 584960 650268
rect -960 649348 480 649588
rect 583520 645948 584960 646188
rect -960 645268 480 645508
rect 583520 641868 584960 642108
rect -960 641188 480 641428
rect 583520 637788 584960 638028
rect -960 637108 480 637348
rect 583520 633708 584960 633948
rect -960 633028 480 633268
rect 583520 629628 584960 629868
rect -960 628948 480 629188
rect 583520 626228 584960 626468
rect -960 624868 480 625108
rect 583520 622148 584960 622388
rect -960 621468 480 621708
rect 583520 618068 584960 618308
rect -960 617388 480 617628
rect 583520 613988 584960 614228
rect -960 613308 480 613548
rect 583520 609908 584960 610148
rect -960 609228 480 609468
rect 583520 605828 584960 606068
rect -960 605148 480 605388
rect 583520 601748 584960 601988
rect -960 601068 480 601308
rect 583520 597668 584960 597908
rect -960 596988 480 597228
rect 583520 593588 584960 593828
rect -960 592908 480 593148
rect 583520 589508 584960 589748
rect -960 588828 480 589068
rect 583520 586108 584960 586348
rect -960 584748 480 584988
rect 583520 582028 584960 582268
rect -960 581348 480 581588
rect 583520 577948 584960 578188
rect -960 577268 480 577508
rect 583520 573868 584960 574108
rect -960 573188 480 573428
rect 583520 569788 584960 570028
rect -960 569108 480 569348
rect 583520 565708 584960 565948
rect -960 565028 480 565268
rect 583520 561628 584960 561868
rect -960 560948 480 561188
rect 583520 557548 584960 557788
rect -960 556868 480 557108
rect 583520 553468 584960 553708
rect -960 552788 480 553028
rect 583520 549388 584960 549628
rect -960 548708 480 548948
rect 583520 545988 584960 546228
rect -960 544628 480 544868
rect 583520 541908 584960 542148
rect -960 541228 480 541468
rect 583520 537828 584960 538068
rect -960 537148 480 537388
rect 583520 533748 584960 533988
rect -960 533068 480 533308
rect 583520 529668 584960 529908
rect -960 528988 480 529228
rect 583520 525588 584960 525828
rect -960 524908 480 525148
rect 583520 521508 584960 521748
rect -960 520828 480 521068
rect 583520 517428 584960 517668
rect -960 516748 480 516988
rect 583520 513348 584960 513588
rect -960 512668 480 512908
rect 583520 509948 584960 510188
rect -960 508588 480 508828
rect 583520 505868 584960 506108
rect -960 504508 480 504748
rect 583520 501788 584960 502028
rect -960 501108 480 501348
rect 583520 497708 584960 497948
rect -960 497028 480 497268
rect 583520 493628 584960 493868
rect -960 492948 480 493188
rect 583520 489548 584960 489788
rect -960 488868 480 489108
rect 583520 485468 584960 485708
rect -960 484788 480 485028
rect 583520 481388 584960 481628
rect -960 480708 480 480948
rect 583520 477308 584960 477548
rect -960 476628 480 476868
rect 583520 473228 584960 473468
rect -960 472548 480 472788
rect 583520 469828 584960 470068
rect -960 468468 480 468708
rect 583520 465748 584960 465988
rect -960 465068 480 465308
rect 583520 461668 584960 461908
rect -960 460988 480 461228
rect 583520 457588 584960 457828
rect -960 456908 480 457148
rect 583520 453508 584960 453748
rect -960 452828 480 453068
rect 583520 449428 584960 449668
rect -960 448748 480 448988
rect 583520 445348 584960 445588
rect -960 444668 480 444908
rect 583520 441268 584960 441508
rect -960 440588 480 440828
rect 583520 437188 584960 437428
rect -960 436508 480 436748
rect 583520 433108 584960 433348
rect -960 432428 480 432668
rect 583520 429708 584960 429948
rect -960 428348 480 428588
rect 583520 425628 584960 425868
rect -960 424948 480 425188
rect 583520 421548 584960 421788
rect -960 420868 480 421108
rect 583520 417468 584960 417708
rect -960 416788 480 417028
rect 583520 413388 584960 413628
rect -960 412708 480 412948
rect 583520 409308 584960 409548
rect -960 408628 480 408868
rect 583520 405228 584960 405468
rect -960 404548 480 404788
rect 583520 401148 584960 401388
rect -960 400468 480 400708
rect 583520 397068 584960 397308
rect -960 396388 480 396628
rect 583520 392988 584960 393228
rect -960 392308 480 392548
rect 583520 389588 584960 389828
rect -960 388228 480 388468
rect 583520 385508 584960 385748
rect -960 384828 480 385068
rect 583520 381428 584960 381668
rect -960 380748 480 380988
rect 583520 377348 584960 377588
rect -960 376668 480 376908
rect 583520 373268 584960 373508
rect -960 372588 480 372828
rect 583520 369188 584960 369428
rect -960 368508 480 368748
rect 583520 365108 584960 365348
rect -960 364428 480 364668
rect 583520 361028 584960 361268
rect -960 360348 480 360588
rect 583520 356948 584960 357188
rect -960 356268 480 356508
rect 583520 353548 584960 353788
rect -960 352188 480 352428
rect 583520 349468 584960 349708
rect -960 348788 480 349028
rect 583520 345388 584960 345628
rect -960 344708 480 344948
rect 583520 341308 584960 341548
rect -960 340628 480 340868
rect 583520 337228 584960 337468
rect -960 336548 480 336788
rect 583520 333148 584960 333388
rect -960 332468 480 332708
rect 583520 329068 584960 329308
rect -960 328388 480 328628
rect 583520 324988 584960 325228
rect -960 324308 480 324548
rect 583520 320908 584960 321148
rect -960 320228 480 320468
rect 583520 316828 584960 317068
rect -960 316148 480 316388
rect 583520 313428 584960 313668
rect -960 312068 480 312308
rect 583520 309348 584960 309588
rect -960 308668 480 308908
rect 583520 305268 584960 305508
rect -960 304588 480 304828
rect 583520 301188 584960 301428
rect -960 300508 480 300748
rect 583520 297108 584960 297348
rect -960 296428 480 296668
rect 583520 293028 584960 293268
rect -960 292348 480 292588
rect 583520 288948 584960 289188
rect -960 288268 480 288508
rect 583520 284868 584960 285108
rect -960 284188 480 284428
rect 583520 280788 584960 281028
rect -960 280108 480 280348
rect 583520 276708 584960 276948
rect -960 276028 480 276268
rect 583520 273308 584960 273548
rect -960 271948 480 272188
rect 583520 269228 584960 269468
rect -960 268548 480 268788
rect 583520 265148 584960 265388
rect -960 264468 480 264708
rect 583520 261068 584960 261308
rect -960 260388 480 260628
rect 583520 256988 584960 257228
rect -960 256308 480 256548
rect 583520 252908 584960 253148
rect -960 252228 480 252468
rect 583520 248828 584960 249068
rect -960 248148 480 248388
rect 583520 244748 584960 244988
rect -960 244068 480 244308
rect 583520 240668 584960 240908
rect -960 239988 480 240228
rect 583520 237268 584960 237508
rect -960 235908 480 236148
rect 583520 233188 584960 233428
rect -960 232508 480 232748
rect 583520 229108 584960 229348
rect -960 228428 480 228668
rect 583520 225028 584960 225268
rect -960 224348 480 224588
rect 583520 220948 584960 221188
rect -960 220268 480 220508
rect 583520 216868 584960 217108
rect -960 216188 480 216428
rect 583520 212788 584960 213028
rect -960 212108 480 212348
rect 583520 208708 584960 208948
rect -960 208028 480 208268
rect 583520 204628 584960 204868
rect -960 203948 480 204188
rect 583520 200548 584960 200788
rect -960 199868 480 200108
rect 583520 197148 584960 197388
rect -960 195788 480 196028
rect 583520 193068 584960 193308
rect -960 192388 480 192628
rect 583520 188988 584960 189228
rect -960 188308 480 188548
rect 583520 184908 584960 185148
rect -960 184228 480 184468
rect 583520 180828 584960 181068
rect -960 180148 480 180388
rect 583520 176748 584960 176988
rect -960 176068 480 176308
rect 583520 172668 584960 172908
rect -960 171988 480 172228
rect 583520 168588 584960 168828
rect -960 167908 480 168148
rect 583520 164508 584960 164748
rect -960 163828 480 164068
rect 583520 160428 584960 160668
rect -960 159748 480 159988
rect 583520 157028 584960 157268
rect -960 155668 480 155908
rect 583520 152948 584960 153188
rect -960 152268 480 152508
rect 583520 148868 584960 149108
rect -960 148188 480 148428
rect 583520 144788 584960 145028
rect -960 144108 480 144348
rect 583520 140708 584960 140948
rect -960 140028 480 140268
rect 583520 136628 584960 136868
rect -960 135948 480 136188
rect 583520 132548 584960 132788
rect -960 131868 480 132108
rect 583520 128468 584960 128708
rect -960 127788 480 128028
rect 583520 124388 584960 124628
rect -960 123708 480 123948
rect 583520 120988 584960 121228
rect -960 119628 480 119868
rect 583520 116908 584960 117148
rect -960 116228 480 116468
rect 583520 112828 584960 113068
rect -960 112148 480 112388
rect 583520 108748 584960 108988
rect -960 108068 480 108308
rect 583520 104668 584960 104908
rect -960 103988 480 104228
rect 583520 100588 584960 100828
rect -960 99908 480 100148
rect 583520 96508 584960 96748
rect -960 95828 480 96068
rect 583520 92428 584960 92668
rect -960 91748 480 91988
rect 583520 88348 584960 88588
rect -960 87668 480 87908
rect 583520 84268 584960 84508
rect -960 83588 480 83828
rect 583520 80868 584960 81108
rect -960 79508 480 79748
rect 583520 76788 584960 77028
rect -960 76108 480 76348
rect 583520 72708 584960 72948
rect -960 72028 480 72268
rect 583520 68628 584960 68868
rect -960 67948 480 68188
rect 583520 64548 584960 64788
rect -960 63868 480 64108
rect 583520 60468 584960 60708
rect -960 59788 480 60028
rect 583520 56388 584960 56628
rect -960 55708 480 55948
rect 583520 52308 584960 52548
rect -960 51628 480 51868
rect 583520 48228 584960 48468
rect -960 47548 480 47788
rect 583520 44148 584960 44388
rect -960 43468 480 43708
rect 583520 40748 584960 40988
rect -960 39388 480 39628
rect 583520 36668 584960 36908
rect -960 35988 480 36228
rect 583520 32588 584960 32828
rect -960 31908 480 32148
rect 583520 28508 584960 28748
rect -960 27828 480 28068
rect 583520 24428 584960 24668
rect -960 23748 480 23988
rect 583520 20348 584960 20588
rect -960 19668 480 19908
rect 583520 16268 584960 16508
rect -960 15588 480 15828
rect 583520 12188 584960 12428
rect -960 11508 480 11748
rect 583520 8108 584960 8348
rect -960 7428 480 7668
rect 583520 4708 584960 4948
rect -960 3348 480 3588
rect 583520 628 584960 868
<< obsm3 >>
rect 246 702308 583440 702541
rect 246 701348 583586 702308
rect 560 700948 583586 701348
rect 246 698628 583586 700948
rect 246 698228 583440 698628
rect 246 697948 583586 698228
rect 560 697548 583586 697948
rect 246 694548 583586 697548
rect 246 694148 583440 694548
rect 246 693868 583586 694148
rect 560 693468 583586 693868
rect 246 690468 583586 693468
rect 246 690068 583440 690468
rect 246 689788 583586 690068
rect 560 689388 583586 689788
rect 246 686388 583586 689388
rect 246 685988 583440 686388
rect 246 685708 583586 685988
rect 560 685308 583586 685708
rect 246 682308 583586 685308
rect 246 681908 583440 682308
rect 246 681628 583586 681908
rect 560 681228 583586 681628
rect 246 678228 583586 681228
rect 246 677828 583440 678228
rect 246 677548 583586 677828
rect 560 677148 583586 677548
rect 246 674148 583586 677148
rect 246 673748 583440 674148
rect 246 673468 583586 673748
rect 560 673068 583586 673468
rect 246 670068 583586 673068
rect 246 669668 583440 670068
rect 246 669388 583586 669668
rect 560 668988 583586 669388
rect 246 665988 583586 668988
rect 246 665588 583440 665988
rect 246 665308 583586 665588
rect 560 664908 583586 665308
rect 246 662588 583586 664908
rect 246 662188 583440 662588
rect 246 661228 583586 662188
rect 560 660828 583586 661228
rect 246 658508 583586 660828
rect 246 658108 583440 658508
rect 246 657828 583586 658108
rect 560 657428 583586 657828
rect 246 654428 583586 657428
rect 246 654028 583440 654428
rect 246 653748 583586 654028
rect 560 653348 583586 653748
rect 246 650348 583586 653348
rect 246 649948 583440 650348
rect 246 649668 583586 649948
rect 560 649268 583586 649668
rect 246 646268 583586 649268
rect 246 645868 583440 646268
rect 246 645588 583586 645868
rect 560 645188 583586 645588
rect 246 642188 583586 645188
rect 246 641788 583440 642188
rect 246 641508 583586 641788
rect 560 641108 583586 641508
rect 246 638108 583586 641108
rect 246 637708 583440 638108
rect 246 637428 583586 637708
rect 560 637028 583586 637428
rect 246 634028 583586 637028
rect 246 633628 583440 634028
rect 246 633348 583586 633628
rect 560 632948 583586 633348
rect 246 629948 583586 632948
rect 246 629548 583440 629948
rect 246 629268 583586 629548
rect 560 628868 583586 629268
rect 246 626548 583586 628868
rect 246 626148 583440 626548
rect 246 625188 583586 626148
rect 560 624788 583586 625188
rect 246 622468 583586 624788
rect 246 622068 583440 622468
rect 246 621788 583586 622068
rect 560 621388 583586 621788
rect 246 618388 583586 621388
rect 246 617988 583440 618388
rect 246 617708 583586 617988
rect 560 617308 583586 617708
rect 246 614308 583586 617308
rect 246 613908 583440 614308
rect 246 613628 583586 613908
rect 560 613228 583586 613628
rect 246 610228 583586 613228
rect 246 609828 583440 610228
rect 246 609548 583586 609828
rect 560 609148 583586 609548
rect 246 606148 583586 609148
rect 246 605748 583440 606148
rect 246 605468 583586 605748
rect 560 605068 583586 605468
rect 246 602068 583586 605068
rect 246 601668 583440 602068
rect 246 601388 583586 601668
rect 560 600988 583586 601388
rect 246 597988 583586 600988
rect 246 597588 583440 597988
rect 246 597308 583586 597588
rect 560 596908 583586 597308
rect 246 593908 583586 596908
rect 246 593508 583440 593908
rect 246 593228 583586 593508
rect 560 592828 583586 593228
rect 246 589828 583586 592828
rect 246 589428 583440 589828
rect 246 589148 583586 589428
rect 560 588748 583586 589148
rect 246 586428 583586 588748
rect 246 586028 583440 586428
rect 246 585068 583586 586028
rect 560 584668 583586 585068
rect 246 582348 583586 584668
rect 246 581948 583440 582348
rect 246 581668 583586 581948
rect 560 581268 583586 581668
rect 246 578268 583586 581268
rect 246 577868 583440 578268
rect 246 577588 583586 577868
rect 560 577188 583586 577588
rect 246 574188 583586 577188
rect 246 573788 583440 574188
rect 246 573508 583586 573788
rect 560 573108 583586 573508
rect 246 570108 583586 573108
rect 246 569708 583440 570108
rect 246 569428 583586 569708
rect 560 569028 583586 569428
rect 246 566028 583586 569028
rect 246 565628 583440 566028
rect 246 565348 583586 565628
rect 560 564948 583586 565348
rect 246 561948 583586 564948
rect 246 561548 583440 561948
rect 246 561268 583586 561548
rect 560 560868 583586 561268
rect 246 557868 583586 560868
rect 246 557468 583440 557868
rect 246 557188 583586 557468
rect 560 556788 583586 557188
rect 246 553788 583586 556788
rect 246 553388 583440 553788
rect 246 553108 583586 553388
rect 560 552708 583586 553108
rect 246 549708 583586 552708
rect 246 549308 583440 549708
rect 246 549028 583586 549308
rect 560 548628 583586 549028
rect 246 546308 583586 548628
rect 246 545908 583440 546308
rect 246 544948 583586 545908
rect 560 544548 583586 544948
rect 246 542228 583586 544548
rect 246 541828 583440 542228
rect 246 541548 583586 541828
rect 560 541148 583586 541548
rect 246 538148 583586 541148
rect 246 537748 583440 538148
rect 246 537468 583586 537748
rect 560 537068 583586 537468
rect 246 534068 583586 537068
rect 246 533668 583440 534068
rect 246 533388 583586 533668
rect 560 532988 583586 533388
rect 246 529988 583586 532988
rect 246 529588 583440 529988
rect 246 529308 583586 529588
rect 560 528908 583586 529308
rect 246 525908 583586 528908
rect 246 525508 583440 525908
rect 246 525228 583586 525508
rect 560 524828 583586 525228
rect 246 521828 583586 524828
rect 246 521428 583440 521828
rect 246 521148 583586 521428
rect 560 520748 583586 521148
rect 246 517748 583586 520748
rect 246 517348 583440 517748
rect 246 517068 583586 517348
rect 560 516668 583586 517068
rect 246 513668 583586 516668
rect 246 513268 583440 513668
rect 246 512988 583586 513268
rect 560 512588 583586 512988
rect 246 510268 583586 512588
rect 246 509868 583440 510268
rect 246 508908 583586 509868
rect 560 508508 583586 508908
rect 246 506188 583586 508508
rect 246 505788 583440 506188
rect 246 504828 583586 505788
rect 560 504428 583586 504828
rect 246 502108 583586 504428
rect 246 501708 583440 502108
rect 246 501428 583586 501708
rect 560 501028 583586 501428
rect 246 498028 583586 501028
rect 246 497628 583440 498028
rect 246 497348 583586 497628
rect 560 496948 583586 497348
rect 246 493948 583586 496948
rect 246 493548 583440 493948
rect 246 493268 583586 493548
rect 560 492868 583586 493268
rect 246 489868 583586 492868
rect 246 489468 583440 489868
rect 246 489188 583586 489468
rect 560 488788 583586 489188
rect 246 485788 583586 488788
rect 246 485388 583440 485788
rect 246 485108 583586 485388
rect 560 484708 583586 485108
rect 246 481708 583586 484708
rect 246 481308 583440 481708
rect 246 481028 583586 481308
rect 560 480628 583586 481028
rect 246 477628 583586 480628
rect 246 477228 583440 477628
rect 246 476948 583586 477228
rect 560 476548 583586 476948
rect 246 473548 583586 476548
rect 246 473148 583440 473548
rect 246 472868 583586 473148
rect 560 472468 583586 472868
rect 246 470148 583586 472468
rect 246 469748 583440 470148
rect 246 468788 583586 469748
rect 560 468388 583586 468788
rect 246 466068 583586 468388
rect 246 465668 583440 466068
rect 246 465388 583586 465668
rect 560 464988 583586 465388
rect 246 461988 583586 464988
rect 246 461588 583440 461988
rect 246 461308 583586 461588
rect 560 460908 583586 461308
rect 246 457908 583586 460908
rect 246 457508 583440 457908
rect 246 457228 583586 457508
rect 560 456828 583586 457228
rect 246 453828 583586 456828
rect 246 453428 583440 453828
rect 246 453148 583586 453428
rect 560 452748 583586 453148
rect 246 449748 583586 452748
rect 246 449348 583440 449748
rect 246 449068 583586 449348
rect 560 448668 583586 449068
rect 246 445668 583586 448668
rect 246 445268 583440 445668
rect 246 444988 583586 445268
rect 560 444588 583586 444988
rect 246 441588 583586 444588
rect 246 441188 583440 441588
rect 246 440908 583586 441188
rect 560 440508 583586 440908
rect 246 437508 583586 440508
rect 246 437108 583440 437508
rect 246 436828 583586 437108
rect 560 436428 583586 436828
rect 246 433428 583586 436428
rect 246 433028 583440 433428
rect 246 432748 583586 433028
rect 560 432348 583586 432748
rect 246 430028 583586 432348
rect 246 429628 583440 430028
rect 246 428668 583586 429628
rect 560 428268 583586 428668
rect 246 425948 583586 428268
rect 246 425548 583440 425948
rect 246 425268 583586 425548
rect 560 424868 583586 425268
rect 246 421868 583586 424868
rect 246 421468 583440 421868
rect 246 421188 583586 421468
rect 560 420788 583586 421188
rect 246 417788 583586 420788
rect 246 417388 583440 417788
rect 246 417108 583586 417388
rect 560 416708 583586 417108
rect 246 413708 583586 416708
rect 246 413308 583440 413708
rect 246 413028 583586 413308
rect 560 412628 583586 413028
rect 246 409628 583586 412628
rect 246 409228 583440 409628
rect 246 408948 583586 409228
rect 560 408548 583586 408948
rect 246 405548 583586 408548
rect 246 405148 583440 405548
rect 246 404868 583586 405148
rect 560 404468 583586 404868
rect 246 401468 583586 404468
rect 246 401068 583440 401468
rect 246 400788 583586 401068
rect 560 400388 583586 400788
rect 246 397388 583586 400388
rect 246 396988 583440 397388
rect 246 396708 583586 396988
rect 560 396308 583586 396708
rect 246 393308 583586 396308
rect 246 392908 583440 393308
rect 246 392628 583586 392908
rect 560 392228 583586 392628
rect 246 389908 583586 392228
rect 246 389508 583440 389908
rect 246 388548 583586 389508
rect 560 388148 583586 388548
rect 246 385828 583586 388148
rect 246 385428 583440 385828
rect 246 385148 583586 385428
rect 560 384748 583586 385148
rect 246 381748 583586 384748
rect 246 381348 583440 381748
rect 246 381068 583586 381348
rect 560 380668 583586 381068
rect 246 377668 583586 380668
rect 246 377268 583440 377668
rect 246 376988 583586 377268
rect 560 376588 583586 376988
rect 246 373588 583586 376588
rect 246 373188 583440 373588
rect 246 372908 583586 373188
rect 560 372508 583586 372908
rect 246 369508 583586 372508
rect 246 369108 583440 369508
rect 246 368828 583586 369108
rect 560 368428 583586 368828
rect 246 365428 583586 368428
rect 246 365028 583440 365428
rect 246 364748 583586 365028
rect 560 364348 583586 364748
rect 246 361348 583586 364348
rect 246 360948 583440 361348
rect 246 360668 583586 360948
rect 560 360268 583586 360668
rect 246 357268 583586 360268
rect 246 356868 583440 357268
rect 246 356588 583586 356868
rect 560 356188 583586 356588
rect 246 353868 583586 356188
rect 246 353468 583440 353868
rect 246 352508 583586 353468
rect 560 352108 583586 352508
rect 246 349788 583586 352108
rect 246 349388 583440 349788
rect 246 349108 583586 349388
rect 560 348708 583586 349108
rect 246 345708 583586 348708
rect 246 345308 583440 345708
rect 246 345028 583586 345308
rect 560 344628 583586 345028
rect 246 341628 583586 344628
rect 246 341228 583440 341628
rect 246 340948 583586 341228
rect 560 340548 583586 340948
rect 246 337548 583586 340548
rect 246 337148 583440 337548
rect 246 336868 583586 337148
rect 560 336468 583586 336868
rect 246 333468 583586 336468
rect 246 333068 583440 333468
rect 246 332788 583586 333068
rect 560 332388 583586 332788
rect 246 329388 583586 332388
rect 246 328988 583440 329388
rect 246 328708 583586 328988
rect 560 328308 583586 328708
rect 246 325308 583586 328308
rect 246 324908 583440 325308
rect 246 324628 583586 324908
rect 560 324228 583586 324628
rect 246 321228 583586 324228
rect 246 320828 583440 321228
rect 246 320548 583586 320828
rect 560 320148 583586 320548
rect 246 317148 583586 320148
rect 246 316748 583440 317148
rect 246 316468 583586 316748
rect 560 316068 583586 316468
rect 246 313748 583586 316068
rect 246 313348 583440 313748
rect 246 312388 583586 313348
rect 560 311988 583586 312388
rect 246 309668 583586 311988
rect 246 309268 583440 309668
rect 246 308988 583586 309268
rect 560 308588 583586 308988
rect 246 305588 583586 308588
rect 246 305188 583440 305588
rect 246 304908 583586 305188
rect 560 304508 583586 304908
rect 246 301508 583586 304508
rect 246 301108 583440 301508
rect 246 300828 583586 301108
rect 560 300428 583586 300828
rect 246 297428 583586 300428
rect 246 297028 583440 297428
rect 246 296748 583586 297028
rect 560 296348 583586 296748
rect 246 293348 583586 296348
rect 246 292948 583440 293348
rect 246 292668 583586 292948
rect 560 292268 583586 292668
rect 246 289268 583586 292268
rect 246 288868 583440 289268
rect 246 288588 583586 288868
rect 560 288188 583586 288588
rect 246 285188 583586 288188
rect 246 284788 583440 285188
rect 246 284508 583586 284788
rect 560 284108 583586 284508
rect 246 281108 583586 284108
rect 246 280708 583440 281108
rect 246 280428 583586 280708
rect 560 280028 583586 280428
rect 246 277028 583586 280028
rect 246 276628 583440 277028
rect 246 276348 583586 276628
rect 560 275948 583586 276348
rect 246 273628 583586 275948
rect 246 273228 583440 273628
rect 246 272268 583586 273228
rect 560 271868 583586 272268
rect 246 269548 583586 271868
rect 246 269148 583440 269548
rect 246 268868 583586 269148
rect 560 268468 583586 268868
rect 246 265468 583586 268468
rect 246 265068 583440 265468
rect 246 264788 583586 265068
rect 560 264388 583586 264788
rect 246 261388 583586 264388
rect 246 260988 583440 261388
rect 246 260708 583586 260988
rect 560 260308 583586 260708
rect 246 257308 583586 260308
rect 246 256908 583440 257308
rect 246 256628 583586 256908
rect 560 256228 583586 256628
rect 246 253228 583586 256228
rect 246 252828 583440 253228
rect 246 252548 583586 252828
rect 560 252148 583586 252548
rect 246 249148 583586 252148
rect 246 248748 583440 249148
rect 246 248468 583586 248748
rect 560 248068 583586 248468
rect 246 245068 583586 248068
rect 246 244668 583440 245068
rect 246 244388 583586 244668
rect 560 243988 583586 244388
rect 246 240988 583586 243988
rect 246 240588 583440 240988
rect 246 240308 583586 240588
rect 560 239908 583586 240308
rect 246 237588 583586 239908
rect 246 237188 583440 237588
rect 246 236228 583586 237188
rect 560 235828 583586 236228
rect 246 233508 583586 235828
rect 246 233108 583440 233508
rect 246 232828 583586 233108
rect 560 232428 583586 232828
rect 246 229428 583586 232428
rect 246 229028 583440 229428
rect 246 228748 583586 229028
rect 560 228348 583586 228748
rect 246 225348 583586 228348
rect 246 224948 583440 225348
rect 246 224668 583586 224948
rect 560 224268 583586 224668
rect 246 221268 583586 224268
rect 246 220868 583440 221268
rect 246 220588 583586 220868
rect 560 220188 583586 220588
rect 246 217188 583586 220188
rect 246 216788 583440 217188
rect 246 216508 583586 216788
rect 560 216108 583586 216508
rect 246 213108 583586 216108
rect 246 212708 583440 213108
rect 246 212428 583586 212708
rect 560 212028 583586 212428
rect 246 209028 583586 212028
rect 246 208628 583440 209028
rect 246 208348 583586 208628
rect 560 207948 583586 208348
rect 246 204948 583586 207948
rect 246 204548 583440 204948
rect 246 204268 583586 204548
rect 560 203868 583586 204268
rect 246 200868 583586 203868
rect 246 200468 583440 200868
rect 246 200188 583586 200468
rect 560 199788 583586 200188
rect 246 197468 583586 199788
rect 246 197068 583440 197468
rect 246 196108 583586 197068
rect 560 195708 583586 196108
rect 246 193388 583586 195708
rect 246 192988 583440 193388
rect 246 192708 583586 192988
rect 560 192308 583586 192708
rect 246 189308 583586 192308
rect 246 188908 583440 189308
rect 246 188628 583586 188908
rect 560 188228 583586 188628
rect 246 185228 583586 188228
rect 246 184828 583440 185228
rect 246 184548 583586 184828
rect 560 184148 583586 184548
rect 246 181148 583586 184148
rect 246 180748 583440 181148
rect 246 180468 583586 180748
rect 560 180068 583586 180468
rect 246 177068 583586 180068
rect 246 176668 583440 177068
rect 246 176388 583586 176668
rect 560 175988 583586 176388
rect 246 172988 583586 175988
rect 246 172588 583440 172988
rect 246 172308 583586 172588
rect 560 171908 583586 172308
rect 246 168908 583586 171908
rect 246 168508 583440 168908
rect 246 168228 583586 168508
rect 560 167828 583586 168228
rect 246 164828 583586 167828
rect 246 164428 583440 164828
rect 246 164148 583586 164428
rect 560 163748 583586 164148
rect 246 160748 583586 163748
rect 246 160348 583440 160748
rect 246 160068 583586 160348
rect 560 159668 583586 160068
rect 246 157348 583586 159668
rect 246 156948 583440 157348
rect 246 155988 583586 156948
rect 560 155588 583586 155988
rect 246 153268 583586 155588
rect 246 152868 583440 153268
rect 246 152588 583586 152868
rect 560 152188 583586 152588
rect 246 149188 583586 152188
rect 246 148788 583440 149188
rect 246 148508 583586 148788
rect 560 148108 583586 148508
rect 246 145108 583586 148108
rect 246 144708 583440 145108
rect 246 144428 583586 144708
rect 560 144028 583586 144428
rect 246 141028 583586 144028
rect 246 140628 583440 141028
rect 246 140348 583586 140628
rect 560 139948 583586 140348
rect 246 136948 583586 139948
rect 246 136548 583440 136948
rect 246 136268 583586 136548
rect 560 135868 583586 136268
rect 246 132868 583586 135868
rect 246 132468 583440 132868
rect 246 132188 583586 132468
rect 560 131788 583586 132188
rect 246 128788 583586 131788
rect 246 128388 583440 128788
rect 246 128108 583586 128388
rect 560 127708 583586 128108
rect 246 124708 583586 127708
rect 246 124308 583440 124708
rect 246 124028 583586 124308
rect 560 123628 583586 124028
rect 246 121308 583586 123628
rect 246 120908 583440 121308
rect 246 119948 583586 120908
rect 560 119548 583586 119948
rect 246 117228 583586 119548
rect 246 116828 583440 117228
rect 246 116548 583586 116828
rect 560 116148 583586 116548
rect 246 113148 583586 116148
rect 246 112748 583440 113148
rect 246 112468 583586 112748
rect 560 112068 583586 112468
rect 246 109068 583586 112068
rect 246 108668 583440 109068
rect 246 108388 583586 108668
rect 560 107988 583586 108388
rect 246 104988 583586 107988
rect 246 104588 583440 104988
rect 246 104308 583586 104588
rect 560 103908 583586 104308
rect 246 100908 583586 103908
rect 246 100508 583440 100908
rect 246 100228 583586 100508
rect 560 99828 583586 100228
rect 246 96828 583586 99828
rect 246 96428 583440 96828
rect 246 96148 583586 96428
rect 560 95748 583586 96148
rect 246 92748 583586 95748
rect 246 92348 583440 92748
rect 246 92068 583586 92348
rect 560 91668 583586 92068
rect 246 88668 583586 91668
rect 246 88268 583440 88668
rect 246 87988 583586 88268
rect 560 87588 583586 87988
rect 246 84588 583586 87588
rect 246 84188 583440 84588
rect 246 83908 583586 84188
rect 560 83508 583586 83908
rect 246 81188 583586 83508
rect 246 80788 583440 81188
rect 246 79828 583586 80788
rect 560 79428 583586 79828
rect 246 77108 583586 79428
rect 246 76708 583440 77108
rect 246 76428 583586 76708
rect 560 76028 583586 76428
rect 246 73028 583586 76028
rect 246 72628 583440 73028
rect 246 72348 583586 72628
rect 560 71948 583586 72348
rect 246 68948 583586 71948
rect 246 68548 583440 68948
rect 246 68268 583586 68548
rect 560 67868 583586 68268
rect 246 64868 583586 67868
rect 246 64468 583440 64868
rect 246 64188 583586 64468
rect 560 63788 583586 64188
rect 246 60788 583586 63788
rect 246 60388 583440 60788
rect 246 60108 583586 60388
rect 560 59708 583586 60108
rect 246 56708 583586 59708
rect 246 56308 583440 56708
rect 246 56028 583586 56308
rect 560 55628 583586 56028
rect 246 52628 583586 55628
rect 246 52228 583440 52628
rect 246 51948 583586 52228
rect 560 51548 583586 51948
rect 246 48548 583586 51548
rect 246 48148 583440 48548
rect 246 47868 583586 48148
rect 560 47468 583586 47868
rect 246 44468 583586 47468
rect 246 44068 583440 44468
rect 246 43788 583586 44068
rect 560 43388 583586 43788
rect 246 41068 583586 43388
rect 246 40668 583440 41068
rect 246 39708 583586 40668
rect 560 39308 583586 39708
rect 246 36988 583586 39308
rect 246 36588 583440 36988
rect 246 36308 583586 36588
rect 560 35908 583586 36308
rect 246 32908 583586 35908
rect 246 32508 583440 32908
rect 246 32228 583586 32508
rect 560 31828 583586 32228
rect 246 28828 583586 31828
rect 246 28428 583440 28828
rect 246 28148 583586 28428
rect 560 27748 583586 28148
rect 246 24748 583586 27748
rect 246 24348 583440 24748
rect 246 24068 583586 24348
rect 560 23668 583586 24068
rect 246 20668 583586 23668
rect 246 20268 583440 20668
rect 246 19988 583586 20268
rect 560 19588 583586 19988
rect 246 16588 583586 19588
rect 246 16188 583440 16588
rect 246 15908 583586 16188
rect 560 15508 583586 15908
rect 246 12508 583586 15508
rect 246 12108 583440 12508
rect 246 11828 583586 12108
rect 560 11428 583586 11828
rect 246 8428 583586 11428
rect 246 8028 583440 8428
rect 246 7748 583586 8028
rect 560 7348 583586 7748
rect 246 5028 583586 7348
rect 246 4628 583440 5028
rect 246 3668 583586 4628
rect 560 3268 583586 3668
rect 246 948 583586 3268
rect 246 715 583440 948
<< metal4 >>
rect -8726 -7654 -8106 711590
rect -7766 -6694 -7146 710630
rect -6806 -5734 -6186 709670
rect -5846 -4774 -5226 708710
rect -4886 -3814 -4266 707750
rect -3926 -2854 -3306 706790
rect -2966 -1894 -2346 705830
rect -2006 -934 -1386 704870
rect 1794 -7654 2414 711590
rect 6294 -7654 6914 711590
rect 10794 -7654 11414 711590
rect 15294 -7654 15914 711590
rect 19794 -7654 20414 711590
rect 24294 -7654 24914 711590
rect 28794 -7654 29414 711590
rect 33294 -7654 33914 711590
rect 37794 -7654 38414 711590
rect 42294 -7654 42914 711590
rect 46794 -7654 47414 711590
rect 51294 -7654 51914 711590
rect 55794 -7654 56414 711590
rect 60294 -7654 60914 711590
rect 64794 -7654 65414 711590
rect 69294 -7654 69914 711590
rect 73794 -7654 74414 711590
rect 78294 -7654 78914 711590
rect 82794 -7654 83414 711590
rect 87294 -7654 87914 711590
rect 91794 -7654 92414 711590
rect 96294 -7654 96914 711590
rect 100794 -7654 101414 711590
rect 105294 -7654 105914 711590
rect 109794 -7654 110414 711590
rect 114294 -7654 114914 711590
rect 118794 262000 119414 711590
rect 123294 262000 123914 711590
rect 127794 262000 128414 711590
rect 132294 262000 132914 711590
rect 136794 262000 137414 711590
rect 141294 262000 141914 711590
rect 145794 262000 146414 711590
rect 150294 262000 150914 711590
rect 154794 262000 155414 711590
rect 159294 262000 159914 711590
rect 163794 262000 164414 711590
rect 168294 262000 168914 711590
rect 172794 262000 173414 711590
rect 177294 262000 177914 711590
rect 181794 262000 182414 711590
rect 186294 262000 186914 711590
rect 190794 262000 191414 711590
rect 118794 142000 119414 198000
rect 123294 142000 123914 198000
rect 141294 142000 141914 198000
rect 145794 142000 146414 198000
rect 150294 142000 150914 198000
rect 154794 142000 155414 198000
rect 159294 142000 159914 198000
rect 177294 142000 177914 198000
rect 181794 142000 182414 198000
rect 186294 142000 186914 198000
rect 190794 142000 191414 198000
rect 118794 -7654 119414 78000
rect 123294 -7654 123914 78000
rect 127794 -7654 128414 78000
rect 132294 -7654 132914 78000
rect 136794 -7654 137414 78000
rect 141294 -7654 141914 78000
rect 145794 -7654 146414 78000
rect 150294 -7654 150914 78000
rect 154794 -7654 155414 78000
rect 159294 -7654 159914 78000
rect 163794 -7654 164414 78000
rect 168294 -7654 168914 78000
rect 172794 -7654 173414 78000
rect 177294 -7654 177914 78000
rect 181794 -7654 182414 78000
rect 186294 -7654 186914 78000
rect 190794 -7654 191414 78000
rect 195294 -7654 195914 711590
rect 199794 -7654 200414 711590
rect 204294 -7654 204914 711590
rect 208794 -7654 209414 711590
rect 213294 -7654 213914 711590
rect 217794 -7654 218414 711590
rect 222294 -7654 222914 711590
rect 226794 -7654 227414 711590
rect 231294 -7654 231914 711590
rect 235794 -7654 236414 711590
rect 240294 -7654 240914 711590
rect 244794 -7654 245414 711590
rect 249294 -7654 249914 711590
rect 253794 -7654 254414 711590
rect 258294 -7654 258914 711590
rect 262794 -7654 263414 711590
rect 267294 -7654 267914 711590
rect 271794 -7654 272414 711590
rect 276294 -7654 276914 711590
rect 280794 -7654 281414 711590
rect 285294 -7654 285914 711590
rect 289794 -7654 290414 711590
rect 294294 -7654 294914 711590
rect 298794 -7654 299414 711590
rect 303294 -7654 303914 711590
rect 307794 -7654 308414 711590
rect 312294 -7654 312914 711590
rect 316794 -7654 317414 711590
rect 321294 -7654 321914 711590
rect 325794 -7654 326414 711590
rect 330294 -7654 330914 711590
rect 334794 -7654 335414 711590
rect 339294 -7654 339914 711590
rect 343794 -7654 344414 711590
rect 348294 -7654 348914 711590
rect 352794 -7654 353414 711590
rect 357294 -7654 357914 711590
rect 361794 -7654 362414 711590
rect 366294 -7654 366914 711590
rect 370794 -7654 371414 711590
rect 375294 -7654 375914 711590
rect 379794 -7654 380414 711590
rect 384294 -7654 384914 711590
rect 388794 -7654 389414 711590
rect 393294 -7654 393914 711590
rect 397794 -7654 398414 711590
rect 402294 -7654 402914 711590
rect 406794 -7654 407414 711590
rect 411294 -7654 411914 711590
rect 415794 -7654 416414 711590
rect 420294 -7654 420914 711590
rect 424794 -7654 425414 711590
rect 429294 -7654 429914 711590
rect 433794 -7654 434414 711590
rect 438294 -7654 438914 711590
rect 442794 -7654 443414 711590
rect 447294 -7654 447914 711590
rect 451794 -7654 452414 711590
rect 456294 -7654 456914 711590
rect 460794 -7654 461414 711590
rect 465294 -7654 465914 711590
rect 469794 -7654 470414 711590
rect 474294 -7654 474914 711590
rect 478794 -7654 479414 711590
rect 483294 -7654 483914 711590
rect 487794 -7654 488414 711590
rect 492294 -7654 492914 711590
rect 496794 -7654 497414 711590
rect 501294 -7654 501914 711590
rect 505794 -7654 506414 711590
rect 510294 -7654 510914 711590
rect 514794 -7654 515414 711590
rect 519294 -7654 519914 711590
rect 523794 -7654 524414 711590
rect 528294 -7654 528914 711590
rect 532794 -7654 533414 711590
rect 537294 -7654 537914 711590
rect 541794 -7654 542414 711590
rect 546294 -7654 546914 711590
rect 550794 -7654 551414 711590
rect 555294 -7654 555914 711590
rect 559794 -7654 560414 711590
rect 564294 -7654 564914 711590
rect 568794 -7654 569414 711590
rect 573294 -7654 573914 711590
rect 577794 -7654 578414 711590
rect 582294 -7654 582914 711590
rect 585310 -934 585930 704870
rect 586270 -1894 586890 705830
rect 587230 -2854 587850 706790
rect 588190 -3814 588810 707750
rect 589150 -4774 589770 708710
rect 590110 -5734 590730 709670
rect 591070 -6694 591690 710630
rect 592030 -7654 592650 711590
<< obsm4 >>
rect 95739 34443 96214 656981
rect 96994 34443 100714 656981
rect 101494 34443 105214 656981
rect 105994 34443 109714 656981
rect 110494 34443 114214 656981
rect 114994 261920 118714 656981
rect 119494 261920 123214 656981
rect 123994 261920 127714 656981
rect 128494 261920 132214 656981
rect 132994 261920 136714 656981
rect 137494 261920 141214 656981
rect 141994 261920 145714 656981
rect 146494 261920 150214 656981
rect 150994 261920 154714 656981
rect 155494 261920 159214 656981
rect 159994 261920 163714 656981
rect 164494 261920 168214 656981
rect 168994 261920 172714 656981
rect 173494 261920 177214 656981
rect 177994 261920 181714 656981
rect 182494 261920 186214 656981
rect 186994 261920 190714 656981
rect 191494 261920 195214 656981
rect 114994 198080 195214 261920
rect 114994 141920 118714 198080
rect 119494 141920 123214 198080
rect 123994 141920 141214 198080
rect 141994 141920 145714 198080
rect 146494 141920 150214 198080
rect 150994 141920 154714 198080
rect 155494 141920 159214 198080
rect 159994 141920 177214 198080
rect 177994 141920 181714 198080
rect 182494 141920 186214 198080
rect 186994 141920 190714 198080
rect 191494 141920 195214 198080
rect 114994 78080 195214 141920
rect 114994 34443 118714 78080
rect 119494 34443 123214 78080
rect 123994 34443 127714 78080
rect 128494 34443 132214 78080
rect 132994 34443 136714 78080
rect 137494 34443 141214 78080
rect 141994 34443 145714 78080
rect 146494 34443 150214 78080
rect 150994 34443 154714 78080
rect 155494 34443 159214 78080
rect 159994 34443 163714 78080
rect 164494 34443 168214 78080
rect 168994 34443 172714 78080
rect 173494 34443 177214 78080
rect 177994 34443 181714 78080
rect 182494 34443 186214 78080
rect 186994 34443 190714 78080
rect 191494 34443 195214 78080
rect 195994 34443 199714 656981
rect 200494 34443 204214 656981
rect 204994 34443 208714 656981
rect 209494 34443 211173 656981
<< metal5 >>
rect -8726 710970 592650 711590
rect -7766 710010 591690 710630
rect -6806 709050 590730 709670
rect -5846 708090 589770 708710
rect -4886 707130 588810 707750
rect -3926 706170 587850 706790
rect -2966 705210 586890 705830
rect -2006 704250 585930 704870
rect -8726 700366 592650 700986
rect -8726 695866 592650 696486
rect -8726 691366 592650 691986
rect -8726 686866 592650 687486
rect -8726 682366 592650 682986
rect -8726 677866 592650 678486
rect -8726 673366 592650 673986
rect -8726 668866 592650 669486
rect -8726 664366 592650 664986
rect -8726 659866 592650 660486
rect -8726 655366 592650 655986
rect -8726 650866 592650 651486
rect -8726 646366 592650 646986
rect -8726 641866 592650 642486
rect -8726 637366 592650 637986
rect -8726 632866 592650 633486
rect -8726 628366 592650 628986
rect -8726 623866 592650 624486
rect -8726 619366 592650 619986
rect -8726 614866 592650 615486
rect -8726 610366 592650 610986
rect -8726 605866 592650 606486
rect -8726 601366 592650 601986
rect -8726 596866 592650 597486
rect -8726 592366 592650 592986
rect -8726 587866 592650 588486
rect -8726 583366 592650 583986
rect -8726 578866 592650 579486
rect -8726 574366 592650 574986
rect -8726 569866 592650 570486
rect -8726 565366 592650 565986
rect -8726 560866 592650 561486
rect -8726 556366 592650 556986
rect -8726 551866 592650 552486
rect -8726 547366 592650 547986
rect -8726 542866 592650 543486
rect -8726 538366 592650 538986
rect -8726 533866 592650 534486
rect -8726 529366 592650 529986
rect -8726 524866 592650 525486
rect -8726 520366 592650 520986
rect -8726 515866 592650 516486
rect -8726 511366 592650 511986
rect -8726 506866 592650 507486
rect -8726 502366 592650 502986
rect -8726 497866 592650 498486
rect -8726 493366 592650 493986
rect -8726 488866 592650 489486
rect -8726 484366 592650 484986
rect -8726 479866 592650 480486
rect -8726 475366 592650 475986
rect -8726 470866 592650 471486
rect -8726 466366 592650 466986
rect -8726 461866 592650 462486
rect -8726 457366 592650 457986
rect -8726 452866 592650 453486
rect -8726 448366 592650 448986
rect -8726 443866 592650 444486
rect -8726 439366 592650 439986
rect -8726 434866 592650 435486
rect -8726 430366 592650 430986
rect -8726 425866 592650 426486
rect -8726 421366 592650 421986
rect -8726 416866 592650 417486
rect -8726 412366 592650 412986
rect -8726 407866 592650 408486
rect -8726 403366 592650 403986
rect -8726 398866 592650 399486
rect -8726 394366 592650 394986
rect -8726 389866 592650 390486
rect -8726 385366 592650 385986
rect -8726 380866 592650 381486
rect -8726 376366 592650 376986
rect -8726 371866 592650 372486
rect -8726 367366 592650 367986
rect -8726 362866 592650 363486
rect -8726 358366 592650 358986
rect -8726 353866 592650 354486
rect -8726 349366 592650 349986
rect -8726 344866 592650 345486
rect -8726 340366 592650 340986
rect -8726 335866 592650 336486
rect -8726 331366 592650 331986
rect -8726 326866 592650 327486
rect -8726 322366 592650 322986
rect -8726 317866 592650 318486
rect -8726 313366 592650 313986
rect -8726 308866 592650 309486
rect -8726 304366 592650 304986
rect -8726 299866 592650 300486
rect -8726 295366 592650 295986
rect -8726 290866 592650 291486
rect -8726 286366 592650 286986
rect -8726 281866 592650 282486
rect -8726 277366 592650 277986
rect -8726 272866 592650 273486
rect -8726 268366 592650 268986
rect -8726 263866 592650 264486
rect -8726 259366 592650 259986
rect -8726 254866 592650 255486
rect -8726 250366 592650 250986
rect -8726 245866 592650 246486
rect -8726 241366 592650 241986
rect -8726 236866 592650 237486
rect -8726 232366 592650 232986
rect -8726 227866 592650 228486
rect -8726 223366 592650 223986
rect -8726 218866 592650 219486
rect -8726 214366 592650 214986
rect -8726 209866 592650 210486
rect -8726 205366 592650 205986
rect -8726 200866 592650 201486
rect -8726 196366 592650 196986
rect -8726 191866 592650 192486
rect -8726 187366 592650 187986
rect -8726 182866 592650 183486
rect -8726 178366 592650 178986
rect -8726 173866 592650 174486
rect -8726 169366 592650 169986
rect -8726 164866 592650 165486
rect -8726 160366 592650 160986
rect -8726 155866 592650 156486
rect -8726 151366 592650 151986
rect -8726 146866 592650 147486
rect -8726 142366 592650 142986
rect -8726 137866 592650 138486
rect -8726 133366 592650 133986
rect -8726 128866 592650 129486
rect -8726 124366 592650 124986
rect -8726 119866 592650 120486
rect -8726 115366 592650 115986
rect -8726 110866 592650 111486
rect -8726 106366 592650 106986
rect -8726 101866 592650 102486
rect -8726 97366 592650 97986
rect -8726 92866 592650 93486
rect -8726 88366 592650 88986
rect -8726 83866 592650 84486
rect -8726 79366 592650 79986
rect -8726 74866 592650 75486
rect -8726 70366 592650 70986
rect -8726 65866 592650 66486
rect -8726 61366 592650 61986
rect -8726 56866 592650 57486
rect -8726 52366 592650 52986
rect -8726 47866 592650 48486
rect -8726 43366 592650 43986
rect -8726 38866 592650 39486
rect -8726 34366 592650 34986
rect -8726 29866 592650 30486
rect -8726 25366 592650 25986
rect -8726 20866 592650 21486
rect -8726 16366 592650 16986
rect -8726 11866 592650 12486
rect -8726 7366 592650 7986
rect -8726 2866 592650 3486
rect -2006 -934 585930 -314
rect -2966 -1894 586890 -1274
rect -3926 -2854 587850 -2234
rect -4886 -3814 588810 -3194
rect -5846 -4774 589770 -4154
rect -6806 -5734 590730 -5114
rect -7766 -6694 591690 -6074
rect -8726 -7654 592650 -7034
<< labels >>
rlabel metal2 s 506174 703520 506286 704960 6 gpio_analog[0]
port 1 nsew signal bidirectional
rlabel metal2 s 159058 -960 159170 480 8 gpio_analog[10]
port 2 nsew signal bidirectional
rlabel metal3 s 583520 417468 584960 417708 6 gpio_analog[11]
port 3 nsew signal bidirectional
rlabel metal3 s -960 573188 480 573428 4 gpio_analog[12]
port 4 nsew signal bidirectional
rlabel metal3 s 583520 593588 584960 593828 6 gpio_analog[13]
port 5 nsew signal bidirectional
rlabel metal2 s 56662 -960 56774 480 8 gpio_analog[14]
port 6 nsew signal bidirectional
rlabel metal2 s 160346 703520 160458 704960 6 gpio_analog[15]
port 7 nsew signal bidirectional
rlabel metal3 s 583520 212788 584960 213028 6 gpio_analog[16]
port 8 nsew signal bidirectional
rlabel metal3 s -960 501108 480 501348 4 gpio_analog[17]
port 9 nsew signal bidirectional
rlabel metal2 s 223458 -960 223570 480 8 gpio_analog[1]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 229108 584960 229348 6 gpio_analog[2]
port 11 nsew signal bidirectional
rlabel metal3 s -960 268548 480 268788 4 gpio_analog[3]
port 12 nsew signal bidirectional
rlabel metal2 s 428894 -960 429006 480 8 gpio_analog[4]
port 13 nsew signal bidirectional
rlabel metal3 s 583520 124388 584960 124628 6 gpio_analog[5]
port 14 nsew signal bidirectional
rlabel metal3 s 583520 513348 584960 513588 6 gpio_analog[6]
port 15 nsew signal bidirectional
rlabel metal2 s 270470 703520 270582 704960 6 gpio_analog[7]
port 16 nsew signal bidirectional
rlabel metal3 s 583520 329068 584960 329308 6 gpio_analog[8]
port 17 nsew signal bidirectional
rlabel metal2 s 405710 -960 405822 480 8 gpio_analog[9]
port 18 nsew signal bidirectional
rlabel metal2 s 37342 -960 37454 480 8 gpio_noesd[0]
port 19 nsew signal bidirectional
rlabel metal3 s 583520 136628 584960 136868 6 gpio_noesd[10]
port 20 nsew signal bidirectional
rlabel metal2 s 337446 -960 337558 480 8 gpio_noesd[11]
port 21 nsew signal bidirectional
rlabel metal2 s 440486 -960 440598 480 8 gpio_noesd[12]
port 22 nsew signal bidirectional
rlabel metal3 s -960 276028 480 276268 4 gpio_noesd[13]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 409308 584960 409548 6 gpio_noesd[14]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 120988 584960 121228 6 gpio_noesd[15]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 665668 584960 665908 6 gpio_noesd[16]
port 26 nsew signal bidirectional
rlabel metal2 s 367714 -960 367826 480 8 gpio_noesd[17]
port 27 nsew signal bidirectional
rlabel metal2 s 292366 -960 292478 480 8 gpio_noesd[1]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 324988 584960 325228 6 gpio_noesd[2]
port 29 nsew signal bidirectional
rlabel metal3 s 583520 421548 584960 421788 6 gpio_noesd[3]
port 30 nsew signal bidirectional
rlabel metal2 s 569286 -960 569398 480 8 gpio_noesd[4]
port 31 nsew signal bidirectional
rlabel metal2 s 224746 703520 224858 704960 6 gpio_noesd[5]
port 32 nsew signal bidirectional
rlabel metal3 s -960 669068 480 669308 4 gpio_noesd[6]
port 33 nsew signal bidirectional
rlabel metal2 s 372866 703520 372978 704960 6 gpio_noesd[7]
port 34 nsew signal bidirectional
rlabel metal2 s 413438 -960 413550 480 8 gpio_noesd[8]
port 35 nsew signal bidirectional
rlabel metal3 s 583520 633708 584960 633948 6 gpio_noesd[9]
port 36 nsew signal bidirectional
rlabel metal3 s -960 148188 480 148428 4 io_analog[0]
port 37 nsew signal bidirectional
rlabel metal2 s 238914 -960 239026 480 8 io_analog[10]
port 38 nsew signal bidirectional
rlabel metal2 s 130078 703520 130190 704960 6 io_analog[1]
port 39 nsew signal bidirectional
rlabel metal3 s -960 31908 480 32148 4 io_analog[2]
port 40 nsew signal bidirectional
rlabel metal3 s -960 203948 480 204188 4 io_analog[3]
port 41 nsew signal bidirectional
rlabel metal2 s 60526 -960 60638 480 8 io_analog[4]
port 42 nsew signal bidirectional
rlabel metal2 s 296874 703520 296986 704960 6 io_analog[5]
port 43 nsew signal bidirectional
rlabel metal3 s -960 693548 480 693788 4 io_analog[6]
port 44 nsew signal bidirectional
rlabel metal3 s 583520 561628 584960 561868 6 io_analog[7]
port 45 nsew signal bidirectional
rlabel metal3 s -960 673148 480 673388 4 io_analog[8]
port 46 nsew signal bidirectional
rlabel metal2 s 388322 703520 388434 704960 6 io_analog[9]
port 47 nsew signal bidirectional
rlabel metal2 s 186750 703520 186862 704960 6 io_clamp_high[0]
port 48 nsew signal bidirectional
rlabel metal3 s -960 424948 480 425188 4 io_clamp_high[1]
port 49 nsew signal bidirectional
rlabel metal2 s 22530 -960 22642 480 8 io_clamp_high[2]
port 50 nsew signal bidirectional
rlabel metal3 s 583520 618068 584960 618308 6 io_clamp_low[0]
port 51 nsew signal bidirectional
rlabel metal3 s 583520 160428 584960 160668 6 io_clamp_low[1]
port 52 nsew signal bidirectional
rlabel metal3 s -960 55708 480 55948 4 io_clamp_low[2]
port 53 nsew signal bidirectional
rlabel metal3 s 583520 537828 584960 538068 6 io_in[0]
port 54 nsew signal input
rlabel metal3 s 583520 356948 584960 357188 6 io_in[10]
port 55 nsew signal input
rlabel metal3 s 583520 92428 584960 92668 6 io_in[11]
port 56 nsew signal input
rlabel metal2 s 113334 -960 113446 480 8 io_in[12]
port 57 nsew signal input
rlabel metal2 s 34766 703520 34878 704960 6 io_in[13]
port 58 nsew signal input
rlabel metal2 s 441130 703520 441242 704960 6 io_in[14]
port 59 nsew signal input
rlabel metal3 s 583520 216868 584960 217108 6 io_in[15]
port 60 nsew signal input
rlabel metal2 s 493294 -960 493406 480 8 io_in[16]
port 61 nsew signal input
rlabel metal3 s 583520 381428 584960 381668 6 io_in[17]
port 62 nsew signal input
rlabel metal2 s 147466 -960 147578 480 8 io_in[18]
port 63 nsew signal input
rlabel metal3 s -960 533068 480 533308 4 io_in[19]
port 64 nsew signal input
rlabel metal2 s 95946 703520 96058 704960 6 io_in[1]
port 65 nsew signal input
rlabel metal2 s 361918 703520 362030 704960 6 io_in[20]
port 66 nsew signal input
rlabel metal2 s 68898 703520 69010 704960 6 io_in[21]
port 67 nsew signal input
rlabel metal2 s 417302 -960 417414 480 8 io_in[22]
port 68 nsew signal input
rlabel metal2 s 136518 -960 136630 480 8 io_in[23]
port 69 nsew signal input
rlabel metal3 s -960 239988 480 240228 4 io_in[24]
port 70 nsew signal input
rlabel metal2 s 133942 703520 134054 704960 6 io_in[25]
port 71 nsew signal input
rlabel metal3 s 583520 485468 584960 485708 6 io_in[26]
port 72 nsew signal input
rlabel metal2 s 98522 -960 98634 480 8 io_in[2]
port 73 nsew signal input
rlabel metal2 s 83066 -960 83178 480 8 io_in[3]
port 74 nsew signal input
rlabel metal3 s 583520 565708 584960 565948 6 io_in[4]
port 75 nsew signal input
rlabel metal2 s 288502 -960 288614 480 8 io_in[5]
port 76 nsew signal input
rlabel metal3 s -960 617388 480 617628 4 io_in[6]
port 77 nsew signal input
rlabel metal3 s -960 340628 480 340868 4 io_in[7]
port 78 nsew signal input
rlabel metal3 s 583520 68628 584960 68868 6 io_in[8]
port 79 nsew signal input
rlabel metal3 s -960 192388 480 192628 4 io_in[9]
port 80 nsew signal input
rlabel metal2 s 338734 703520 338846 704960 6 io_in_3v3[0]
port 81 nsew signal input
rlabel metal3 s -960 392308 480 392548 4 io_in_3v3[10]
port 82 nsew signal input
rlabel metal2 s 86930 -960 87042 480 8 io_in_3v3[11]
port 83 nsew signal input
rlabel metal2 s 258878 703520 258990 704960 6 io_in_3v3[12]
port 84 nsew signal input
rlabel metal2 s 122350 703520 122462 704960 6 io_in_3v3[13]
port 85 nsew signal input
rlabel metal3 s -960 312068 480 312308 4 io_in_3v3[14]
port 86 nsew signal input
rlabel metal3 s 583520 148868 584960 149108 6 io_in_3v3[15]
port 87 nsew signal input
rlabel metal3 s -960 176068 480 176308 4 io_in_3v3[16]
port 88 nsew signal input
rlabel metal2 s 10938 -960 11050 480 8 io_in_3v3[17]
port 89 nsew signal input
rlabel metal3 s -960 649348 480 649588 4 io_in_3v3[18]
port 90 nsew signal input
rlabel metal2 s 414726 703520 414838 704960 6 io_in_3v3[19]
port 91 nsew signal input
rlabel metal3 s 583520 577948 584960 578188 6 io_in_3v3[1]
port 92 nsew signal input
rlabel metal3 s -960 420868 480 421108 4 io_in_3v3[20]
port 93 nsew signal input
rlabel metal2 s 217018 703520 217130 704960 6 io_in_3v3[21]
port 94 nsew signal input
rlabel metal2 s 451434 -960 451546 480 8 io_in_3v3[22]
port 95 nsew signal input
rlabel metal3 s 583520 64548 584960 64788 6 io_in_3v3[23]
port 96 nsew signal input
rlabel metal3 s -960 628948 480 629188 4 io_in_3v3[24]
port 97 nsew signal input
rlabel metal3 s 583520 397068 584960 397308 6 io_in_3v3[25]
port 98 nsew signal input
rlabel metal2 s 213798 703520 213910 704960 6 io_in_3v3[26]
port 99 nsew signal input
rlabel metal3 s 583520 650028 584960 650268 6 io_in_3v3[2]
port 100 nsew signal input
rlabel metal3 s -960 565028 480 565268 4 io_in_3v3[3]
port 101 nsew signal input
rlabel metal2 s 126214 703520 126326 704960 6 io_in_3v3[4]
port 102 nsew signal input
rlabel metal2 s 273046 -960 273158 480 8 io_in_3v3[5]
port 103 nsew signal input
rlabel metal3 s 583520 582028 584960 582268 6 io_in_3v3[6]
port 104 nsew signal input
rlabel metal2 s 346462 703520 346574 704960 6 io_in_3v3[7]
port 105 nsew signal input
rlabel metal3 s -960 63868 480 64108 4 io_in_3v3[8]
port 106 nsew signal input
rlabel metal2 s 523562 -960 523674 480 8 io_in_3v3[9]
port 107 nsew signal input
rlabel metal3 s 583520 605828 584960 606068 6 io_oeb[0]
port 108 nsew signal output
rlabel metal3 s 583520 297108 584960 297348 6 io_oeb[10]
port 109 nsew signal output
rlabel metal2 s 289146 703520 289258 704960 6 io_oeb[11]
port 110 nsew signal output
rlabel metal2 s 212510 -960 212622 480 8 io_oeb[12]
port 111 nsew signal output
rlabel metal3 s 583520 204628 584960 204868 6 io_oeb[13]
port 112 nsew signal output
rlabel metal3 s -960 396388 480 396628 4 io_oeb[14]
port 113 nsew signal output
rlabel metal3 s 583520 172668 584960 172908 6 io_oeb[15]
port 114 nsew signal output
rlabel metal3 s 583520 168588 584960 168828 6 io_oeb[16]
port 115 nsew signal output
rlabel metal3 s -960 119628 480 119868 4 io_oeb[17]
port 116 nsew signal output
rlabel metal3 s -960 364428 480 364668 4 io_oeb[18]
port 117 nsew signal output
rlabel metal3 s 583520 84268 584960 84508 6 io_oeb[19]
port 118 nsew signal output
rlabel metal2 s 396050 703520 396162 704960 6 io_oeb[1]
port 119 nsew signal output
rlabel metal3 s -960 271948 480 272188 4 io_oeb[20]
port 120 nsew signal output
rlabel metal3 s -960 87668 480 87908 4 io_oeb[21]
port 121 nsew signal output
rlabel metal3 s 583520 252908 584960 253148 6 io_oeb[22]
port 122 nsew signal output
rlabel metal2 s 166786 -960 166898 480 8 io_oeb[23]
port 123 nsew signal output
rlabel metal3 s -960 588828 480 589068 4 io_oeb[24]
port 124 nsew signal output
rlabel metal2 s 330362 -960 330474 480 8 io_oeb[25]
port 125 nsew signal output
rlabel metal3 s -960 400468 480 400708 4 io_oeb[26]
port 126 nsew signal output
rlabel metal3 s -960 320228 480 320468 4 io_oeb[2]
port 127 nsew signal output
rlabel metal2 s 148754 703520 148866 704960 6 io_oeb[3]
port 128 nsew signal output
rlabel metal2 s 327142 703520 327254 704960 6 io_oeb[4]
port 129 nsew signal output
rlabel metal3 s 583520 76788 584960 77028 6 io_oeb[5]
port 130 nsew signal output
rlabel metal3 s -960 116228 480 116468 4 io_oeb[6]
port 131 nsew signal output
rlabel metal2 s 144890 703520 145002 704960 6 io_oeb[7]
port 132 nsew signal output
rlabel metal2 s 547390 703520 547502 704960 6 io_oeb[8]
port 133 nsew signal output
rlabel metal2 s 128790 -960 128902 480 8 io_oeb[9]
port 134 nsew signal output
rlabel metal3 s -960 23748 480 23988 4 io_out[0]
port 135 nsew signal output
rlabel metal3 s -960 416788 480 417028 4 io_out[10]
port 136 nsew signal output
rlabel metal2 s 512614 -960 512726 480 8 io_out[11]
port 137 nsew signal output
rlabel metal3 s 583520 698308 584960 698548 6 io_out[12]
port 138 nsew signal output
rlabel metal2 s 482990 703520 483102 704960 6 io_out[13]
port 139 nsew signal output
rlabel metal2 s 182886 703520 182998 704960 6 io_out[14]
port 140 nsew signal output
rlabel metal3 s 583520 673828 584960 674068 6 io_out[15]
port 141 nsew signal output
rlabel metal3 s -960 296428 480 296668 4 io_out[16]
port 142 nsew signal output
rlabel metal2 s 38630 703520 38742 704960 6 io_out[17]
port 143 nsew signal output
rlabel metal2 s 570574 703520 570686 704960 6 io_out[18]
port 144 nsew signal output
rlabel metal2 s 468178 703520 468290 704960 6 io_out[19]
port 145 nsew signal output
rlabel metal3 s 583520 658188 584960 658428 6 io_out[1]
port 146 nsew signal output
rlabel metal2 s 285926 703520 286038 704960 6 io_out[20]
port 147 nsew signal output
rlabel metal3 s -960 637108 480 637348 4 io_out[21]
port 148 nsew signal output
rlabel metal2 s 444994 703520 445106 704960 6 io_out[22]
port 149 nsew signal output
rlabel metal3 s 583520 645948 584960 646188 6 io_out[23]
port 150 nsew signal output
rlabel metal3 s -960 3348 480 3588 4 io_out[24]
port 151 nsew signal output
rlabel metal3 s -960 436508 480 436748 4 io_out[25]
port 152 nsew signal output
rlabel metal3 s 583520 60468 584960 60708 6 io_out[26]
port 153 nsew signal output
rlabel metal3 s -960 504508 480 504748 4 io_out[2]
port 154 nsew signal output
rlabel metal3 s 583520 337228 584960 337468 6 io_out[3]
port 155 nsew signal output
rlabel metal3 s -960 701028 480 701268 4 io_out[4]
port 156 nsew signal output
rlabel metal3 s -960 689468 480 689708 4 io_out[5]
port 157 nsew signal output
rlabel metal3 s -960 452828 480 453068 4 io_out[6]
port 158 nsew signal output
rlabel metal2 s 174514 -960 174626 480 8 io_out[7]
port 159 nsew signal output
rlabel metal2 s 45070 -960 45182 480 8 io_out[8]
port 160 nsew signal output
rlabel metal2 s 519698 -960 519810 480 8 io_out[9]
port 161 nsew signal output
rlabel metal2 s 23818 703520 23930 704960 6 la_data_in[0]
port 162 nsew signal input
rlabel metal3 s 583520 597668 584960 597908 6 la_data_in[100]
port 163 nsew signal input
rlabel metal3 s -960 560948 480 561188 4 la_data_in[101]
port 164 nsew signal input
rlabel metal3 s -960 380748 480 380988 4 la_data_in[102]
port 165 nsew signal input
rlabel metal2 s 376730 703520 376842 704960 6 la_data_in[103]
port 166 nsew signal input
rlabel metal2 s 269182 -960 269294 480 8 la_data_in[104]
port 167 nsew signal input
rlabel metal3 s 583520 225028 584960 225268 6 la_data_in[105]
port 168 nsew signal input
rlabel metal3 s 583520 8108 584960 8348 6 la_data_in[106]
port 169 nsew signal input
rlabel metal3 s -960 624868 480 625108 4 la_data_in[107]
port 170 nsew signal input
rlabel metal3 s -960 520828 480 521068 4 la_data_in[108]
port 171 nsew signal input
rlabel metal2 s 485566 -960 485678 480 8 la_data_in[109]
port 172 nsew signal input
rlabel metal3 s -960 47548 480 47788 4 la_data_in[10]
port 173 nsew signal input
rlabel metal3 s 583520 529668 584960 529908 6 la_data_in[110]
port 174 nsew signal input
rlabel metal3 s 583520 24428 584960 24668 6 la_data_in[111]
port 175 nsew signal input
rlabel metal3 s -960 681308 480 681548 4 la_data_in[112]
port 176 nsew signal input
rlabel metal3 s -960 184228 480 184468 4 la_data_in[113]
port 177 nsew signal input
rlabel metal2 s 314906 -960 315018 480 8 la_data_in[114]
port 178 nsew signal input
rlabel metal3 s 583520 389588 584960 389828 6 la_data_in[115]
port 179 nsew signal input
rlabel metal3 s -960 180148 480 180388 4 la_data_in[116]
port 180 nsew signal input
rlabel metal2 s 121062 -960 121174 480 8 la_data_in[117]
port 181 nsew signal input
rlabel metal3 s -960 512668 480 512908 4 la_data_in[118]
port 182 nsew signal input
rlabel metal2 s 447570 -960 447682 480 8 la_data_in[119]
port 183 nsew signal input
rlabel metal2 s 535154 -960 535266 480 8 la_data_in[11]
port 184 nsew signal input
rlabel metal3 s 583520 301188 584960 301428 6 la_data_in[120]
port 185 nsew signal input
rlabel metal2 s 342598 703520 342710 704960 6 la_data_in[121]
port 186 nsew signal input
rlabel metal3 s -960 484788 480 485028 4 la_data_in[122]
port 187 nsew signal input
rlabel metal3 s 583520 493628 584960 493868 6 la_data_in[123]
port 188 nsew signal input
rlabel metal2 s 244066 703520 244178 704960 6 la_data_in[124]
port 189 nsew signal input
rlabel metal2 s 162922 -960 163034 480 8 la_data_in[125]
port 190 nsew signal input
rlabel metal3 s -960 621468 480 621708 4 la_data_in[126]
port 191 nsew signal input
rlabel metal3 s 583520 269228 584960 269468 6 la_data_in[127]
port 192 nsew signal input
rlabel metal3 s -960 444668 480 444908 4 la_data_in[12]
port 193 nsew signal input
rlabel metal2 s 489430 -960 489542 480 8 la_data_in[13]
port 194 nsew signal input
rlabel metal3 s 583520 589508 584960 589748 6 la_data_in[14]
port 195 nsew signal input
rlabel metal3 s 583520 626228 584960 626468 6 la_data_in[15]
port 196 nsew signal input
rlabel metal3 s 583520 425628 584960 425868 6 la_data_in[16]
port 197 nsew signal input
rlabel metal2 s 261454 -960 261566 480 8 la_data_in[17]
port 198 nsew signal input
rlabel metal3 s 583520 553468 584960 553708 6 la_data_in[18]
port 199 nsew signal input
rlabel metal3 s -960 544628 480 544868 4 la_data_in[19]
port 200 nsew signal input
rlabel metal2 s 477838 -960 477950 480 8 la_data_in[1]
port 201 nsew signal input
rlabel metal3 s -960 163828 480 164068 4 la_data_in[20]
port 202 nsew signal input
rlabel metal3 s 583520 108748 584960 108988 6 la_data_in[21]
port 203 nsew signal input
rlabel metal3 s -960 344708 480 344948 4 la_data_in[22]
port 204 nsew signal input
rlabel metal2 s 303314 -960 303426 480 8 la_data_in[23]
port 205 nsew signal input
rlabel metal2 s 517122 703520 517234 704960 6 la_data_in[24]
port 206 nsew signal input
rlabel metal3 s 583520 188988 584960 189228 6 la_data_in[25]
port 207 nsew signal input
rlabel metal2 s 463026 -960 463138 480 8 la_data_in[26]
port 208 nsew signal input
rlabel metal3 s -960 697628 480 697868 4 la_data_in[27]
port 209 nsew signal input
rlabel metal2 s 528714 703520 528826 704960 6 la_data_in[28]
port 210 nsew signal input
rlabel metal3 s -960 605148 480 605388 4 la_data_in[29]
port 211 nsew signal input
rlabel metal3 s -960 304588 480 304828 4 la_data_in[2]
port 212 nsew signal input
rlabel metal2 s 295586 -960 295698 480 8 la_data_in[30]
port 213 nsew signal input
rlabel metal3 s -960 456908 480 457148 4 la_data_in[31]
port 214 nsew signal input
rlabel metal2 s 75338 -960 75450 480 8 la_data_in[32]
port 215 nsew signal input
rlabel metal2 s 175802 703520 175914 704960 6 la_data_in[33]
port 216 nsew signal input
rlabel metal2 s 304602 703520 304714 704960 6 la_data_in[34]
port 217 nsew signal input
rlabel metal3 s -960 332468 480 332708 4 la_data_in[35]
port 218 nsew signal input
rlabel metal3 s -960 657508 480 657748 4 la_data_in[36]
port 219 nsew signal input
rlabel metal3 s 583520 521508 584960 521748 6 la_data_in[37]
port 220 nsew signal input
rlabel metal3 s 583520 453508 584960 453748 6 la_data_in[38]
port 221 nsew signal input
rlabel metal3 s -960 159748 480 159988 4 la_data_in[39]
port 222 nsew signal input
rlabel metal2 s 546746 -960 546858 480 8 la_data_in[3]
port 223 nsew signal input
rlabel metal2 s 540306 703520 540418 704960 6 la_data_in[40]
port 224 nsew signal input
rlabel metal3 s 583520 52308 584960 52548 6 la_data_in[41]
port 225 nsew signal input
rlabel metal3 s 583520 365108 584960 365348 6 la_data_in[42]
port 226 nsew signal input
rlabel metal3 s -960 76108 480 76348 4 la_data_in[43]
port 227 nsew signal input
rlabel metal3 s -960 7428 480 7668 4 la_data_in[44]
port 228 nsew signal input
rlabel metal2 s 204782 -960 204894 480 8 la_data_in[45]
port 229 nsew signal input
rlabel metal3 s -960 144108 480 144348 4 la_data_in[46]
port 230 nsew signal input
rlabel metal3 s 583520 40748 584960 40988 6 la_data_in[47]
port 231 nsew signal input
rlabel metal2 s 151330 -960 151442 480 8 la_data_in[48]
port 232 nsew signal input
rlabel metal2 s 197054 -960 197166 480 8 la_data_in[49]
port 233 nsew signal input
rlabel metal3 s 583520 313428 584960 313668 6 la_data_in[4]
port 234 nsew signal input
rlabel metal2 s 580878 -960 580990 480 8 la_data_in[50]
port 235 nsew signal input
rlabel metal2 s 266606 703520 266718 704960 6 la_data_in[51]
port 236 nsew signal input
rlabel metal3 s -960 428348 480 428588 4 la_data_in[52]
port 237 nsew signal input
rlabel metal3 s -960 123708 480 123948 4 la_data_in[53]
port 238 nsew signal input
rlabel metal2 s 262742 703520 262854 704960 6 la_data_in[54]
port 239 nsew signal input
rlabel metal3 s 583520 509948 584960 510188 6 la_data_in[55]
port 240 nsew signal input
rlabel metal3 s -960 548708 480 548948 4 la_data_in[56]
port 241 nsew signal input
rlabel metal2 s 257590 -960 257702 480 8 la_data_in[57]
port 242 nsew signal input
rlabel metal2 s 3210 -960 3322 480 8 la_data_in[58]
port 243 nsew signal input
rlabel metal3 s 583520 441268 584960 441508 6 la_data_in[59]
port 244 nsew signal input
rlabel metal3 s 583520 32588 584960 32828 6 la_data_in[5]
port 245 nsew signal input
rlabel metal2 s 57950 703520 58062 704960 6 la_data_in[60]
port 246 nsew signal input
rlabel metal3 s 583520 501788 584960 502028 6 la_data_in[61]
port 247 nsew signal input
rlabel metal3 s -960 95828 480 96068 4 la_data_in[62]
port 248 nsew signal input
rlabel metal3 s -960 488868 480 489108 4 la_data_in[63]
port 249 nsew signal input
rlabel metal3 s -960 528988 480 529228 4 la_data_in[64]
port 250 nsew signal input
rlabel metal3 s -960 677228 480 677468 4 la_data_in[65]
port 251 nsew signal input
rlabel metal3 s 583520 56388 584960 56628 6 la_data_in[66]
port 252 nsew signal input
rlabel metal2 s 448858 703520 448970 704960 6 la_data_in[67]
port 253 nsew signal input
rlabel metal3 s 583520 180828 584960 181068 6 la_data_in[68]
port 254 nsew signal input
rlabel metal3 s 583520 586108 584960 586348 6 la_data_in[69]
port 255 nsew signal input
rlabel metal3 s 583520 341308 584960 341548 6 la_data_in[6]
port 256 nsew signal input
rlabel metal2 s 79202 -960 79314 480 8 la_data_in[70]
port 257 nsew signal input
rlabel metal3 s 583520 573868 584960 574108 6 la_data_in[71]
port 258 nsew signal input
rlabel metal3 s -960 308668 480 308908 4 la_data_in[72]
port 259 nsew signal input
rlabel metal2 s 118486 703520 118598 704960 6 la_data_in[73]
port 260 nsew signal input
rlabel metal3 s 583520 549388 584960 549628 6 la_data_in[74]
port 261 nsew signal input
rlabel metal2 s 392186 703520 392298 704960 6 la_data_in[75]
port 262 nsew signal input
rlabel metal2 s 520986 703520 521098 704960 6 la_data_in[76]
port 263 nsew signal input
rlabel metal3 s -960 288268 480 288508 4 la_data_in[77]
port 264 nsew signal input
rlabel metal3 s 583520 333148 584960 333388 6 la_data_in[78]
port 265 nsew signal input
rlabel metal3 s 583520 677908 584960 678148 6 la_data_in[79]
port 266 nsew signal input
rlabel metal2 s 194478 703520 194590 704960 6 la_data_in[7]
port 267 nsew signal input
rlabel metal2 s 494582 703520 494694 704960 6 la_data_in[80]
port 268 nsew signal input
rlabel metal2 s 232474 703520 232586 704960 6 la_data_in[81]
port 269 nsew signal input
rlabel metal3 s -960 480708 480 480948 4 la_data_in[82]
port 270 nsew signal input
rlabel metal3 s -960 72028 480 72268 4 la_data_in[83]
port 271 nsew signal input
rlabel metal2 s 490718 703520 490830 704960 6 la_data_in[84]
port 272 nsew signal input
rlabel metal3 s -960 328388 480 328628 4 la_data_in[85]
port 273 nsew signal input
rlabel metal3 s 583520 349468 584960 349708 6 la_data_in[86]
port 274 nsew signal input
rlabel metal3 s -960 91748 480 91988 4 la_data_in[87]
port 275 nsew signal input
rlabel metal3 s 583520 628 584960 868 6 la_data_in[88]
port 276 nsew signal input
rlabel metal3 s -960 284188 480 284428 4 la_data_in[89]
port 277 nsew signal input
rlabel metal3 s -960 103988 480 104228 4 la_data_in[8]
port 278 nsew signal input
rlabel metal2 s 94658 -960 94770 480 8 la_data_in[90]
port 279 nsew signal input
rlabel metal3 s -960 195788 480 196028 4 la_data_in[91]
port 280 nsew signal input
rlabel metal2 s 254370 -960 254482 480 8 la_data_in[92]
port 281 nsew signal input
rlabel metal2 s 276910 -960 277022 480 8 la_data_in[93]
port 282 nsew signal input
rlabel metal2 s 50222 703520 50334 704960 6 la_data_in[94]
port 283 nsew signal input
rlabel metal2 s 553830 -960 553942 480 8 la_data_in[95]
port 284 nsew signal input
rlabel metal2 s 555118 703520 555230 704960 6 la_data_in[96]
port 285 nsew signal input
rlabel metal3 s -960 232508 480 232748 4 la_data_in[97]
port 286 nsew signal input
rlabel metal3 s 583520 320908 584960 321148 6 la_data_in[98]
port 287 nsew signal input
rlabel metal2 s 189326 -960 189438 480 8 la_data_in[99]
port 288 nsew signal input
rlabel metal3 s -960 508588 480 508828 4 la_data_in[9]
port 289 nsew signal input
rlabel metal3 s -960 609228 480 609468 4 la_data_out[0]
port 290 nsew signal output
rlabel metal2 s 284638 -960 284750 480 8 la_data_out[100]
port 291 nsew signal output
rlabel metal3 s 583520 197148 584960 197388 6 la_data_out[101]
port 292 nsew signal output
rlabel metal3 s 583520 413388 584960 413628 6 la_data_out[102]
port 293 nsew signal output
rlabel metal3 s -960 685388 480 685628 4 la_data_out[103]
port 294 nsew signal output
rlabel metal3 s -960 645268 480 645508 4 la_data_out[104]
port 295 nsew signal output
rlabel metal2 s 231186 -960 231298 480 8 la_data_out[105]
port 296 nsew signal output
rlabel metal2 s 164210 703520 164322 704960 6 la_data_out[106]
port 297 nsew signal output
rlabel metal3 s 583520 261068 584960 261308 6 la_data_out[107]
port 298 nsew signal output
rlabel metal2 s 156482 703520 156594 704960 6 la_data_out[108]
port 299 nsew signal output
rlabel metal2 s 84354 703520 84466 704960 6 la_data_out[109]
port 300 nsew signal output
rlabel metal2 s 155194 -960 155306 480 8 la_data_out[10]
port 301 nsew signal output
rlabel metal3 s 583520 392988 584960 393228 6 la_data_out[110]
port 302 nsew signal output
rlabel metal3 s -960 465068 480 465308 4 la_data_out[111]
port 303 nsew signal output
rlabel metal2 s 502310 703520 502422 704960 6 la_data_out[112]
port 304 nsew signal output
rlabel metal3 s -960 384828 480 385068 4 la_data_out[113]
port 305 nsew signal output
rlabel metal3 s -960 212108 480 212348 4 la_data_out[114]
port 306 nsew signal output
rlabel metal2 s 566710 703520 566822 704960 6 la_data_out[115]
port 307 nsew signal output
rlabel metal3 s -960 497028 480 497268 4 la_data_out[116]
port 308 nsew signal output
rlabel metal2 s 200918 -960 201030 480 8 la_data_out[117]
port 309 nsew signal output
rlabel metal2 s 562846 703520 562958 704960 6 la_data_out[118]
port 310 nsew signal output
rlabel metal3 s -960 67948 480 68188 4 la_data_out[119]
port 311 nsew signal output
rlabel metal2 s 409574 -960 409686 480 8 la_data_out[11]
port 312 nsew signal output
rlabel metal3 s 583520 654108 584960 654348 6 la_data_out[120]
port 313 nsew signal output
rlabel metal3 s 583520 401148 584960 401388 6 la_data_out[121]
port 314 nsew signal output
rlabel metal3 s 583520 28508 584960 28748 6 la_data_out[122]
port 315 nsew signal output
rlabel metal3 s -960 188308 480 188548 4 la_data_out[123]
port 316 nsew signal output
rlabel metal2 s 18666 -960 18778 480 8 la_data_out[124]
port 317 nsew signal output
rlabel metal2 s 179022 703520 179134 704960 6 la_data_out[125]
port 318 nsew signal output
rlabel metal2 s 106894 703520 107006 704960 6 la_data_out[126]
port 319 nsew signal output
rlabel metal2 s 475262 703520 475374 704960 6 la_data_out[127]
port 320 nsew signal output
rlabel metal3 s 583520 140708 584960 140948 6 la_data_out[12]
port 321 nsew signal output
rlabel metal3 s 583520 489548 584960 489788 6 la_data_out[13]
port 322 nsew signal output
rlabel metal3 s -960 27828 480 28068 4 la_data_out[14]
port 323 nsew signal output
rlabel metal3 s 583520 284868 584960 285108 6 la_data_out[15]
port 324 nsew signal output
rlabel metal2 s 227322 -960 227434 480 8 la_data_out[16]
port 325 nsew signal output
rlabel metal3 s 583520 44148 584960 44388 6 la_data_out[17]
port 326 nsew signal output
rlabel metal2 s 394762 -960 394874 480 8 la_data_out[18]
port 327 nsew signal output
rlabel metal2 s 88218 703520 88330 704960 6 la_data_out[19]
port 328 nsew signal output
rlabel metal2 s 334870 703520 334982 704960 6 la_data_out[1]
port 329 nsew signal output
rlabel metal2 s 168074 703520 168186 704960 6 la_data_out[20]
port 330 nsew signal output
rlabel metal2 s 110114 -960 110226 480 8 la_data_out[21]
port 331 nsew signal output
rlabel metal3 s 583520 469828 584960 470068 6 la_data_out[22]
port 332 nsew signal output
rlabel metal3 s -960 448748 480 448988 4 la_data_out[23]
port 333 nsew signal output
rlabel metal2 s 504886 -960 504998 480 8 la_data_out[24]
port 334 nsew signal output
rlabel metal3 s 583520 233188 584960 233428 6 la_data_out[25]
port 335 nsew signal output
rlabel metal2 s 582166 703520 582278 704960 6 la_data_out[26]
port 336 nsew signal output
rlabel metal3 s -960 440588 480 440828 4 la_data_out[27]
port 337 nsew signal output
rlabel metal3 s 583520 16268 584960 16508 6 la_data_out[28]
port 338 nsew signal output
rlabel metal2 s 472042 703520 472154 704960 6 la_data_out[29]
port 339 nsew signal output
rlabel metal3 s 583520 477308 584960 477548 6 la_data_out[2]
port 340 nsew signal output
rlabel metal3 s 583520 377348 584960 377588 6 la_data_out[30]
port 341 nsew signal output
rlabel metal2 s 311042 -960 311154 480 8 la_data_out[31]
port 342 nsew signal output
rlabel metal2 s 307178 -960 307290 480 8 la_data_out[32]
port 343 nsew signal output
rlabel metal3 s -960 412708 480 412948 4 la_data_out[33]
port 344 nsew signal output
rlabel metal3 s 583520 433108 584960 433348 6 la_data_out[34]
port 345 nsew signal output
rlabel metal3 s -960 235908 480 236148 4 la_data_out[35]
port 346 nsew signal output
rlabel metal3 s 583520 316828 584960 317068 6 la_data_out[36]
port 347 nsew signal output
rlabel metal3 s 583520 208708 584960 208948 6 la_data_out[37]
port 348 nsew signal output
rlabel metal3 s -960 127788 480 128028 4 la_data_out[38]
port 349 nsew signal output
rlabel metal3 s 583520 157028 584960 157268 6 la_data_out[39]
port 350 nsew signal output
rlabel metal2 s 524850 703520 524962 704960 6 la_data_out[3]
port 351 nsew signal output
rlabel metal3 s 583520 12188 584960 12428 6 la_data_out[40]
port 352 nsew signal output
rlabel metal3 s 583520 72708 584960 72948 6 la_data_out[41]
port 353 nsew signal output
rlabel metal3 s 583520 132548 584960 132788 6 la_data_out[42]
port 354 nsew signal output
rlabel metal2 s 251794 703520 251906 704960 6 la_data_out[43]
port 355 nsew signal output
rlabel metal3 s 583520 353548 584960 353788 6 la_data_out[44]
port 356 nsew signal output
rlabel metal2 s 322634 -960 322746 480 8 la_data_out[45]
port 357 nsew signal output
rlabel metal2 s 240202 703520 240314 704960 6 la_data_out[46]
port 358 nsew signal output
rlabel metal3 s -960 633028 480 633268 4 la_data_out[47]
port 359 nsew signal output
rlabel metal2 s 470754 -960 470866 480 8 la_data_out[48]
port 360 nsew signal output
rlabel metal2 s 379306 -960 379418 480 8 la_data_out[49]
port 361 nsew signal output
rlabel metal2 s 80490 703520 80602 704960 6 la_data_out[4]
port 362 nsew signal output
rlabel metal2 s 61814 703520 61926 704960 6 la_data_out[50]
port 363 nsew signal output
rlabel metal3 s -960 516748 480 516988 4 la_data_out[51]
port 364 nsew signal output
rlabel metal2 s 141670 703520 141782 704960 6 la_data_out[52]
port 365 nsew signal output
rlabel metal3 s -960 228428 480 228668 4 la_data_out[53]
port 366 nsew signal output
rlabel metal3 s -960 352188 480 352428 4 la_data_out[54]
port 367 nsew signal output
rlabel metal2 s 371578 -960 371690 480 8 la_data_out[55]
port 368 nsew signal output
rlabel metal3 s -960 83588 480 83828 4 la_data_out[56]
port 369 nsew signal output
rlabel metal2 s 434046 703520 434158 704960 6 la_data_out[57]
port 370 nsew signal output
rlabel metal2 s 398626 -960 398738 480 8 la_data_out[58]
port 371 nsew signal output
rlabel metal3 s -960 199868 480 200108 4 la_data_out[59]
port 372 nsew signal output
rlabel metal2 s 274334 703520 274446 704960 6 la_data_out[5]
port 373 nsew signal output
rlabel metal3 s 583520 449428 584960 449668 6 la_data_out[60]
port 374 nsew signal output
rlabel metal3 s 583520 128468 584960 128708 6 la_data_out[61]
port 375 nsew signal output
rlabel metal3 s 583520 429708 584960 429948 6 la_data_out[62]
port 376 nsew signal output
rlabel metal2 s 356766 -960 356878 480 8 la_data_out[63]
port 377 nsew signal output
rlabel metal3 s -960 641188 480 641428 4 la_data_out[64]
port 378 nsew signal output
rlabel metal2 s 452722 703520 452834 704960 6 la_data_out[65]
port 379 nsew signal output
rlabel metal2 s 364494 -960 364606 480 8 la_data_out[66]
port 380 nsew signal output
rlabel metal2 s 430182 703520 430294 704960 6 la_data_out[67]
port 381 nsew signal output
rlabel metal3 s -960 468468 480 468708 4 la_data_out[68]
port 382 nsew signal output
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[69]
port 383 nsew signal output
rlabel metal3 s -960 537148 480 537388 4 la_data_out[6]
port 384 nsew signal output
rlabel metal2 s 190614 703520 190726 704960 6 la_data_out[70]
port 385 nsew signal output
rlabel metal3 s 583520 244748 584960 244988 6 la_data_out[71]
port 386 nsew signal output
rlabel metal3 s 583520 184908 584960 185148 6 la_data_out[72]
port 387 nsew signal output
rlabel metal2 s 318770 -960 318882 480 8 la_data_out[73]
port 388 nsew signal output
rlabel metal2 s 474618 -960 474730 480 8 la_data_out[74]
port 389 nsew signal output
rlabel metal2 s 246642 -960 246754 480 8 la_data_out[75]
port 390 nsew signal output
rlabel metal2 s 437266 703520 437378 704960 6 la_data_out[76]
port 391 nsew signal output
rlabel metal2 s 360630 -960 360742 480 8 la_data_out[77]
port 392 nsew signal output
rlabel metal2 s 634 703520 746 704960 6 la_data_out[78]
port 393 nsew signal output
rlabel metal3 s -960 460988 480 461228 4 la_data_out[79]
port 394 nsew signal output
rlabel metal3 s -960 664988 480 665228 4 la_data_out[7]
port 395 nsew signal output
rlabel metal3 s 583520 481388 584960 481628 6 la_data_out[80]
port 396 nsew signal output
rlabel metal2 s 333582 -960 333694 480 8 la_data_out[81]
port 397 nsew signal output
rlabel metal3 s 583520 152948 584960 153188 6 la_data_out[82]
port 398 nsew signal output
rlabel metal3 s 583520 48228 584960 48468 6 la_data_out[83]
port 399 nsew signal output
rlabel metal3 s 583520 237268 584960 237508 6 la_data_out[84]
port 400 nsew signal output
rlabel metal3 s -960 569108 480 569348 4 la_data_out[85]
port 401 nsew signal output
rlabel metal2 s 250506 -960 250618 480 8 la_data_out[86]
port 402 nsew signal output
rlabel metal3 s -960 59788 480 60028 4 la_data_out[87]
port 403 nsew signal output
rlabel metal2 s 466890 -960 467002 480 8 la_data_out[88]
port 404 nsew signal output
rlabel metal2 s 513258 703520 513370 704960 6 la_data_out[89]
port 405 nsew signal output
rlabel metal2 s 110758 703520 110870 704960 6 la_data_out[8]
port 406 nsew signal output
rlabel metal3 s -960 280108 480 280348 4 la_data_out[90]
port 407 nsew signal output
rlabel metal3 s -960 112148 480 112388 4 la_data_out[91]
port 408 nsew signal output
rlabel metal3 s 583520 80868 584960 81108 6 la_data_out[92]
port 409 nsew signal output
rlabel metal2 s 42494 703520 42606 704960 6 la_data_out[93]
port 410 nsew signal output
rlabel metal2 s 220882 703520 220994 704960 6 la_data_out[94]
port 411 nsew signal output
rlabel metal2 s 425030 -960 425142 480 8 la_data_out[95]
port 412 nsew signal output
rlabel metal3 s -960 368508 480 368748 4 la_data_out[96]
port 413 nsew signal output
rlabel metal3 s -960 208028 480 208268 4 la_data_out[97]
port 414 nsew signal output
rlabel metal2 s 497158 -960 497270 480 8 la_data_out[98]
port 415 nsew signal output
rlabel metal2 s 561558 -960 561670 480 8 la_data_out[99]
port 416 nsew signal output
rlabel metal2 s 4498 703520 4610 704960 6 la_data_out[9]
port 417 nsew signal output
rlabel metal2 s 76626 703520 76738 704960 6 la_oenb[0]
port 418 nsew signal input
rlabel metal2 s 551254 703520 551366 704960 6 la_oenb[100]
port 419 nsew signal input
rlabel metal2 s 515834 -960 515946 480 8 la_oenb[101]
port 420 nsew signal input
rlabel metal2 s 12226 703520 12338 704960 6 la_oenb[102]
port 421 nsew signal input
rlabel metal2 s 422454 703520 422566 704960 6 la_oenb[103]
port 422 nsew signal input
rlabel metal2 s 403134 703520 403246 704960 6 la_oenb[104]
port 423 nsew signal input
rlabel metal3 s -960 476628 480 476868 4 la_oenb[105]
port 424 nsew signal input
rlabel metal2 s 299450 -960 299562 480 8 la_oenb[106]
port 425 nsew signal input
rlabel metal2 s 352902 -960 353014 480 8 la_oenb[107]
port 426 nsew signal input
rlabel metal2 s 532578 703520 532690 704960 6 la_oenb[108]
port 427 nsew signal input
rlabel metal3 s 583520 164508 584960 164748 6 la_oenb[109]
port 428 nsew signal input
rlabel metal2 s 418590 703520 418702 704960 6 la_oenb[10]
port 429 nsew signal input
rlabel metal2 s 170650 -960 170762 480 8 la_oenb[110]
port 430 nsew signal input
rlabel metal3 s 583520 473228 584960 473468 6 la_oenb[111]
port 431 nsew signal input
rlabel metal2 s 171938 703520 172050 704960 6 la_oenb[112]
port 432 nsew signal input
rlabel metal2 s 510038 703520 510150 704960 6 la_oenb[113]
port 433 nsew signal input
rlabel metal2 s 137806 703520 137918 704960 6 la_oenb[114]
port 434 nsew signal input
rlabel metal2 s 31546 703520 31658 704960 6 la_oenb[115]
port 435 nsew signal input
rlabel metal2 s 380594 703520 380706 704960 6 la_oenb[116]
port 436 nsew signal input
rlabel metal3 s -960 324308 480 324548 4 la_oenb[117]
port 437 nsew signal input
rlabel metal3 s 583520 601748 584960 601988 6 la_oenb[118]
port 438 nsew signal input
rlabel metal2 s 481702 -960 481814 480 8 la_oenb[119]
port 439 nsew signal input
rlabel metal3 s 583520 437188 584960 437428 6 la_oenb[11]
port 440 nsew signal input
rlabel metal2 s 124926 -960 125038 480 8 la_oenb[120]
port 441 nsew signal input
rlabel metal3 s -960 79508 480 79748 4 la_oenb[121]
port 442 nsew signal input
rlabel metal3 s -960 432428 480 432668 4 la_oenb[122]
port 443 nsew signal input
rlabel metal2 s 341310 -960 341422 480 8 la_oenb[123]
port 444 nsew signal input
rlabel metal2 s 558982 703520 559094 704960 6 la_oenb[124]
port 445 nsew signal input
rlabel metal3 s -960 376668 480 376908 4 la_oenb[125]
port 446 nsew signal input
rlabel metal3 s -960 336548 480 336788 4 la_oenb[126]
port 447 nsew signal input
rlabel metal2 s 8362 703520 8474 704960 6 la_oenb[127]
port 448 nsew signal input
rlabel metal2 s 46358 703520 46470 704960 6 la_oenb[12]
port 449 nsew signal input
rlabel metal2 s 235050 -960 235162 480 8 la_oenb[13]
port 450 nsew signal input
rlabel metal2 s 282062 703520 282174 704960 6 la_oenb[14]
port 451 nsew signal input
rlabel metal3 s 583520 641868 584960 642108 6 la_oenb[15]
port 452 nsew signal input
rlabel metal3 s 583520 305268 584960 305508 6 la_oenb[16]
port 453 nsew signal input
rlabel metal3 s -960 316148 480 316388 4 la_oenb[17]
port 454 nsew signal input
rlabel metal2 s 542882 -960 542994 480 8 la_oenb[18]
port 455 nsew signal input
rlabel metal3 s 583520 248828 584960 249068 6 la_oenb[19]
port 456 nsew signal input
rlabel metal3 s 583520 545988 584960 546228 6 la_oenb[1]
port 457 nsew signal input
rlabel metal2 s 278198 703520 278310 704960 6 la_oenb[20]
port 458 nsew signal input
rlabel metal3 s -960 152268 480 152508 4 la_oenb[21]
port 459 nsew signal input
rlabel metal2 s 349038 -960 349150 480 8 la_oenb[22]
port 460 nsew signal input
rlabel metal2 s 185462 -960 185574 480 8 la_oenb[23]
port 461 nsew signal input
rlabel metal3 s 583520 193068 584960 193308 6 la_oenb[24]
port 462 nsew signal input
rlabel metal2 s 41206 -960 41318 480 8 la_oenb[25]
port 463 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_oenb[26]
port 464 nsew signal input
rlabel metal3 s 583520 176748 584960 176988 6 la_oenb[27]
port 465 nsew signal input
rlabel metal2 s 578302 703520 578414 704960 6 la_oenb[28]
port 466 nsew signal input
rlabel metal3 s 583520 361028 584960 361268 6 la_oenb[29]
port 467 nsew signal input
rlabel metal2 s 68254 -960 68366 480 8 la_oenb[2]
port 468 nsew signal input
rlabel metal3 s -960 216188 480 216428 4 la_oenb[30]
port 469 nsew signal input
rlabel metal3 s -960 15588 480 15828 4 la_oenb[31]
port 470 nsew signal input
rlabel metal3 s -960 244068 480 244308 4 la_oenb[32]
port 471 nsew signal input
rlabel metal2 s 421166 -960 421278 480 8 la_oenb[33]
port 472 nsew signal input
rlabel metal3 s 583520 445348 584960 445588 6 la_oenb[34]
port 473 nsew signal input
rlabel metal2 s 536442 703520 536554 704960 6 la_oenb[35]
port 474 nsew signal input
rlabel metal3 s -960 596988 480 597228 4 la_oenb[36]
port 475 nsew signal input
rlabel metal2 s 300738 703520 300850 704960 6 la_oenb[37]
port 476 nsew signal input
rlabel metal2 s 544170 703520 544282 704960 6 la_oenb[38]
port 477 nsew signal input
rlabel metal2 s 72762 703520 72874 704960 6 la_oenb[39]
port 478 nsew signal input
rlabel metal3 s -960 300508 480 300748 4 la_oenb[3]
port 479 nsew signal input
rlabel metal3 s 583520 116908 584960 117148 6 la_oenb[40]
port 480 nsew signal input
rlabel metal3 s 583520 293028 584960 293268 6 la_oenb[41]
port 481 nsew signal input
rlabel metal3 s 583520 465748 584960 465988 6 la_oenb[42]
port 482 nsew signal input
rlabel metal2 s 209934 703520 210046 704960 6 la_oenb[43]
port 483 nsew signal input
rlabel metal2 s 501022 -960 501134 480 8 la_oenb[44]
port 484 nsew signal input
rlabel metal3 s -960 653428 480 653668 4 la_oenb[45]
port 485 nsew signal input
rlabel metal3 s -960 99908 480 100148 4 la_oenb[46]
port 486 nsew signal input
rlabel metal2 s 486854 703520 486966 704960 6 la_oenb[47]
port 487 nsew signal input
rlabel metal3 s 583520 681988 584960 682228 6 la_oenb[48]
port 488 nsew signal input
rlabel metal3 s 583520 20348 584960 20588 6 la_oenb[49]
port 489 nsew signal input
rlabel metal3 s -960 11508 480 11748 4 la_oenb[4]
port 490 nsew signal input
rlabel metal2 s 577014 -960 577126 480 8 la_oenb[50]
port 491 nsew signal input
rlabel metal3 s 583520 112828 584960 113068 6 la_oenb[51]
port 492 nsew signal input
rlabel metal2 s 117198 -960 117310 480 8 la_oenb[52]
port 493 nsew signal input
rlabel metal2 s 178378 -960 178490 480 8 la_oenb[53]
port 494 nsew signal input
rlabel metal3 s 583520 36668 584960 36908 6 la_oenb[54]
port 495 nsew signal input
rlabel metal3 s 583520 273308 584960 273548 6 la_oenb[55]
port 496 nsew signal input
rlabel metal3 s 583520 622148 584960 622388 6 la_oenb[56]
port 497 nsew signal input
rlabel metal2 s 228610 703520 228722 704960 6 la_oenb[57]
port 498 nsew signal input
rlabel metal2 s 202206 703520 202318 704960 6 la_oenb[58]
port 499 nsew signal input
rlabel metal2 s 99810 703520 99922 704960 6 la_oenb[59]
port 500 nsew signal input
rlabel metal2 s 220238 -960 220350 480 8 la_oenb[5]
port 501 nsew signal input
rlabel metal3 s 583520 690148 584960 690388 6 la_oenb[60]
port 502 nsew signal input
rlabel metal3 s -960 155668 480 155908 4 la_oenb[61]
port 503 nsew signal input
rlabel metal2 s 65678 703520 65790 704960 6 la_oenb[62]
port 504 nsew signal input
rlabel metal3 s -960 51628 480 51868 4 la_oenb[63]
port 505 nsew signal input
rlabel metal3 s 583520 609908 584960 610148 6 la_oenb[64]
port 506 nsew signal input
rlabel metal2 s 350326 703520 350438 704960 6 la_oenb[65]
port 507 nsew signal input
rlabel metal2 s 312330 703520 312442 704960 6 la_oenb[66]
port 508 nsew signal input
rlabel metal2 s 426318 703520 426430 704960 6 la_oenb[67]
port 509 nsew signal input
rlabel metal2 s 460450 703520 460562 704960 6 la_oenb[68]
port 510 nsew signal input
rlabel metal2 s 464314 703520 464426 704960 6 la_oenb[69]
port 511 nsew signal input
rlabel metal3 s -960 252228 480 252468 4 la_oenb[6]
port 512 nsew signal input
rlabel metal2 s 247930 703520 248042 704960 6 la_oenb[70]
port 513 nsew signal input
rlabel metal3 s -960 224348 480 224588 4 la_oenb[71]
port 514 nsew signal input
rlabel metal2 s 7074 -960 7186 480 8 la_oenb[72]
port 515 nsew signal input
rlabel metal2 s 573150 -960 573262 480 8 la_oenb[73]
port 516 nsew signal input
rlabel metal2 s 387034 -960 387146 480 8 la_oenb[74]
port 517 nsew signal input
rlabel metal3 s 583520 200548 584960 200788 6 la_oenb[75]
port 518 nsew signal input
rlabel metal2 s 316194 703520 316306 704960 6 la_oenb[76]
port 519 nsew signal input
rlabel metal3 s 583520 265148 584960 265388 6 la_oenb[77]
port 520 nsew signal input
rlabel metal3 s -960 581348 480 581588 4 la_oenb[78]
port 521 nsew signal input
rlabel metal2 s 30258 -960 30370 480 8 la_oenb[79]
port 522 nsew signal input
rlabel metal3 s -960 260388 480 260628 4 la_oenb[7]
port 523 nsew signal input
rlabel metal3 s -960 171988 480 172228 4 la_oenb[80]
port 524 nsew signal input
rlabel metal2 s 236338 703520 236450 704960 6 la_oenb[81]
port 525 nsew signal input
rlabel metal3 s 583520 4708 584960 4948 6 la_oenb[82]
port 526 nsew signal input
rlabel metal2 s 280774 -960 280886 480 8 la_oenb[83]
port 527 nsew signal input
rlabel metal3 s -960 492948 480 493188 4 la_oenb[84]
port 528 nsew signal input
rlabel metal3 s 583520 533748 584960 533988 6 la_oenb[85]
port 529 nsew signal input
rlabel metal3 s 583520 669748 584960 669988 6 la_oenb[86]
port 530 nsew signal input
rlabel metal2 s 565422 -960 565534 480 8 la_oenb[87]
port 531 nsew signal input
rlabel metal3 s -960 584748 480 584988 4 la_oenb[88]
port 532 nsew signal input
rlabel metal3 s -960 131868 480 132108 4 la_oenb[89]
port 533 nsew signal input
rlabel metal3 s 583520 637788 584960 638028 6 la_oenb[8]
port 534 nsew signal input
rlabel metal2 s 152618 703520 152730 704960 6 la_oenb[90]
port 535 nsew signal input
rlabel metal3 s -960 39388 480 39628 4 la_oenb[91]
port 536 nsew signal input
rlabel metal2 s 550610 -960 550722 480 8 la_oenb[92]
port 537 nsew signal input
rlabel metal2 s 308466 703520 308578 704960 6 la_oenb[93]
port 538 nsew signal input
rlabel metal3 s 583520 220948 584960 221188 6 la_oenb[94]
port 539 nsew signal input
rlabel metal2 s 103674 703520 103786 704960 6 la_oenb[95]
port 540 nsew signal input
rlabel metal3 s -960 372588 480 372828 4 la_oenb[96]
port 541 nsew signal input
rlabel metal3 s -960 556868 480 557108 4 la_oenb[97]
port 542 nsew signal input
rlabel metal2 s 90794 -960 90906 480 8 la_oenb[98]
port 543 nsew signal input
rlabel metal3 s 583520 517428 584960 517668 6 la_oenb[99]
port 544 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_oenb[9]
port 545 nsew signal input
rlabel metal3 s -960 220268 480 220508 4 pxl_done
port 546 nsew signal output
rlabel metal2 s 182242 -960 182354 480 8 pxl_start_in_path
port 547 nsew signal input
rlabel metal3 s -960 292348 480 292588 4 pxl_start_out_path
port 548 nsew signal input
rlabel metal3 s -960 613308 480 613548 4 serial_data_rlbp_out
port 549 nsew signal output
rlabel metal2 s 320058 703520 320170 704960 6 user_clock2
port 550 nsew signal input
rlabel metal3 s 583520 702388 584960 702628 6 user_irq[0]
port 551 nsew signal output
rlabel metal3 s -960 592908 480 593148 4 user_irq[1]
port 552 nsew signal output
rlabel metal3 s -960 660908 480 661148 4 user_irq[2]
port 553 nsew signal output
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 554 nsew power bidirectional
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 554 nsew power bidirectional
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 554 nsew power bidirectional
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 554 nsew power bidirectional
rlabel metal4 s 1794 -7654 2414 711590 6 vccd1
port 554 nsew power bidirectional
rlabel metal4 s 37794 -7654 38414 711590 6 vccd1
port 554 nsew power bidirectional
rlabel metal4 s 73794 -7654 74414 711590 6 vccd1
port 554 nsew power bidirectional
rlabel metal4 s 109794 -7654 110414 711590 6 vccd1
port 554 nsew power bidirectional
rlabel metal4 s 145794 -7654 146414 78000 6 vccd1
port 554 nsew power bidirectional
rlabel metal4 s 145794 142000 146414 198000 6 vccd1
port 554 nsew power bidirectional
rlabel metal4 s 145794 262000 146414 711590 6 vccd1
port 554 nsew power bidirectional
rlabel metal4 s 181794 -7654 182414 78000 6 vccd1
port 554 nsew power bidirectional
rlabel metal4 s 181794 142000 182414 198000 6 vccd1
port 554 nsew power bidirectional
rlabel metal4 s 181794 262000 182414 711590 6 vccd1
port 554 nsew power bidirectional
rlabel metal4 s 217794 -7654 218414 711590 6 vccd1
port 554 nsew power bidirectional
rlabel metal4 s 253794 -7654 254414 711590 6 vccd1
port 554 nsew power bidirectional
rlabel metal4 s 289794 -7654 290414 711590 6 vccd1
port 554 nsew power bidirectional
rlabel metal4 s 325794 -7654 326414 711590 6 vccd1
port 554 nsew power bidirectional
rlabel metal4 s 361794 -7654 362414 711590 6 vccd1
port 554 nsew power bidirectional
rlabel metal4 s 397794 -7654 398414 711590 6 vccd1
port 554 nsew power bidirectional
rlabel metal4 s 433794 -7654 434414 711590 6 vccd1
port 554 nsew power bidirectional
rlabel metal4 s 469794 -7654 470414 711590 6 vccd1
port 554 nsew power bidirectional
rlabel metal4 s 505794 -7654 506414 711590 6 vccd1
port 554 nsew power bidirectional
rlabel metal4 s 541794 -7654 542414 711590 6 vccd1
port 554 nsew power bidirectional
rlabel metal4 s 577794 -7654 578414 711590 6 vccd1
port 554 nsew power bidirectional
rlabel metal5 s -8726 2866 592650 3486 6 vccd1
port 554 nsew power bidirectional
rlabel metal5 s -8726 38866 592650 39486 6 vccd1
port 554 nsew power bidirectional
rlabel metal5 s -8726 74866 592650 75486 6 vccd1
port 554 nsew power bidirectional
rlabel metal5 s -8726 110866 592650 111486 6 vccd1
port 554 nsew power bidirectional
rlabel metal5 s -8726 146866 592650 147486 6 vccd1
port 554 nsew power bidirectional
rlabel metal5 s -8726 182866 592650 183486 6 vccd1
port 554 nsew power bidirectional
rlabel metal5 s -8726 218866 592650 219486 6 vccd1
port 554 nsew power bidirectional
rlabel metal5 s -8726 254866 592650 255486 6 vccd1
port 554 nsew power bidirectional
rlabel metal5 s -8726 290866 592650 291486 6 vccd1
port 554 nsew power bidirectional
rlabel metal5 s -8726 326866 592650 327486 6 vccd1
port 554 nsew power bidirectional
rlabel metal5 s -8726 362866 592650 363486 6 vccd1
port 554 nsew power bidirectional
rlabel metal5 s -8726 398866 592650 399486 6 vccd1
port 554 nsew power bidirectional
rlabel metal5 s -8726 434866 592650 435486 6 vccd1
port 554 nsew power bidirectional
rlabel metal5 s -8726 470866 592650 471486 6 vccd1
port 554 nsew power bidirectional
rlabel metal5 s -8726 506866 592650 507486 6 vccd1
port 554 nsew power bidirectional
rlabel metal5 s -8726 542866 592650 543486 6 vccd1
port 554 nsew power bidirectional
rlabel metal5 s -8726 578866 592650 579486 6 vccd1
port 554 nsew power bidirectional
rlabel metal5 s -8726 614866 592650 615486 6 vccd1
port 554 nsew power bidirectional
rlabel metal5 s -8726 650866 592650 651486 6 vccd1
port 554 nsew power bidirectional
rlabel metal5 s -8726 686866 592650 687486 6 vccd1
port 554 nsew power bidirectional
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 555 nsew power bidirectional
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 555 nsew power bidirectional
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 555 nsew power bidirectional
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 555 nsew power bidirectional
rlabel metal4 s 10794 -7654 11414 711590 6 vccd2
port 555 nsew power bidirectional
rlabel metal4 s 46794 -7654 47414 711590 6 vccd2
port 555 nsew power bidirectional
rlabel metal4 s 82794 -7654 83414 711590 6 vccd2
port 555 nsew power bidirectional
rlabel metal4 s 118794 -7654 119414 78000 6 vccd2
port 555 nsew power bidirectional
rlabel metal4 s 118794 142000 119414 198000 6 vccd2
port 555 nsew power bidirectional
rlabel metal4 s 118794 262000 119414 711590 6 vccd2
port 555 nsew power bidirectional
rlabel metal4 s 154794 -7654 155414 78000 6 vccd2
port 555 nsew power bidirectional
rlabel metal4 s 154794 142000 155414 198000 6 vccd2
port 555 nsew power bidirectional
rlabel metal4 s 154794 262000 155414 711590 6 vccd2
port 555 nsew power bidirectional
rlabel metal4 s 190794 -7654 191414 78000 6 vccd2
port 555 nsew power bidirectional
rlabel metal4 s 190794 142000 191414 198000 6 vccd2
port 555 nsew power bidirectional
rlabel metal4 s 190794 262000 191414 711590 6 vccd2
port 555 nsew power bidirectional
rlabel metal4 s 226794 -7654 227414 711590 6 vccd2
port 555 nsew power bidirectional
rlabel metal4 s 262794 -7654 263414 711590 6 vccd2
port 555 nsew power bidirectional
rlabel metal4 s 298794 -7654 299414 711590 6 vccd2
port 555 nsew power bidirectional
rlabel metal4 s 334794 -7654 335414 711590 6 vccd2
port 555 nsew power bidirectional
rlabel metal4 s 370794 -7654 371414 711590 6 vccd2
port 555 nsew power bidirectional
rlabel metal4 s 406794 -7654 407414 711590 6 vccd2
port 555 nsew power bidirectional
rlabel metal4 s 442794 -7654 443414 711590 6 vccd2
port 555 nsew power bidirectional
rlabel metal4 s 478794 -7654 479414 711590 6 vccd2
port 555 nsew power bidirectional
rlabel metal4 s 514794 -7654 515414 711590 6 vccd2
port 555 nsew power bidirectional
rlabel metal4 s 550794 -7654 551414 711590 6 vccd2
port 555 nsew power bidirectional
rlabel metal5 s -8726 11866 592650 12486 6 vccd2
port 555 nsew power bidirectional
rlabel metal5 s -8726 47866 592650 48486 6 vccd2
port 555 nsew power bidirectional
rlabel metal5 s -8726 83866 592650 84486 6 vccd2
port 555 nsew power bidirectional
rlabel metal5 s -8726 119866 592650 120486 6 vccd2
port 555 nsew power bidirectional
rlabel metal5 s -8726 155866 592650 156486 6 vccd2
port 555 nsew power bidirectional
rlabel metal5 s -8726 191866 592650 192486 6 vccd2
port 555 nsew power bidirectional
rlabel metal5 s -8726 227866 592650 228486 6 vccd2
port 555 nsew power bidirectional
rlabel metal5 s -8726 263866 592650 264486 6 vccd2
port 555 nsew power bidirectional
rlabel metal5 s -8726 299866 592650 300486 6 vccd2
port 555 nsew power bidirectional
rlabel metal5 s -8726 335866 592650 336486 6 vccd2
port 555 nsew power bidirectional
rlabel metal5 s -8726 371866 592650 372486 6 vccd2
port 555 nsew power bidirectional
rlabel metal5 s -8726 407866 592650 408486 6 vccd2
port 555 nsew power bidirectional
rlabel metal5 s -8726 443866 592650 444486 6 vccd2
port 555 nsew power bidirectional
rlabel metal5 s -8726 479866 592650 480486 6 vccd2
port 555 nsew power bidirectional
rlabel metal5 s -8726 515866 592650 516486 6 vccd2
port 555 nsew power bidirectional
rlabel metal5 s -8726 551866 592650 552486 6 vccd2
port 555 nsew power bidirectional
rlabel metal5 s -8726 587866 592650 588486 6 vccd2
port 555 nsew power bidirectional
rlabel metal5 s -8726 623866 592650 624486 6 vccd2
port 555 nsew power bidirectional
rlabel metal5 s -8726 659866 592650 660486 6 vccd2
port 555 nsew power bidirectional
rlabel metal5 s -8726 695866 592650 696486 6 vccd2
port 555 nsew power bidirectional
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 556 nsew power bidirectional
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 556 nsew power bidirectional
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 556 nsew power bidirectional
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 556 nsew power bidirectional
rlabel metal4 s 19794 -7654 20414 711590 6 vdda1
port 556 nsew power bidirectional
rlabel metal4 s 55794 -7654 56414 711590 6 vdda1
port 556 nsew power bidirectional
rlabel metal4 s 91794 -7654 92414 711590 6 vdda1
port 556 nsew power bidirectional
rlabel metal4 s 127794 -7654 128414 78000 6 vdda1
port 556 nsew power bidirectional
rlabel metal4 s 127794 262000 128414 711590 6 vdda1
port 556 nsew power bidirectional
rlabel metal4 s 163794 -7654 164414 78000 6 vdda1
port 556 nsew power bidirectional
rlabel metal4 s 163794 262000 164414 711590 6 vdda1
port 556 nsew power bidirectional
rlabel metal4 s 199794 -7654 200414 711590 6 vdda1
port 556 nsew power bidirectional
rlabel metal4 s 235794 -7654 236414 711590 6 vdda1
port 556 nsew power bidirectional
rlabel metal4 s 271794 -7654 272414 711590 6 vdda1
port 556 nsew power bidirectional
rlabel metal4 s 307794 -7654 308414 711590 6 vdda1
port 556 nsew power bidirectional
rlabel metal4 s 343794 -7654 344414 711590 6 vdda1
port 556 nsew power bidirectional
rlabel metal4 s 379794 -7654 380414 711590 6 vdda1
port 556 nsew power bidirectional
rlabel metal4 s 415794 -7654 416414 711590 6 vdda1
port 556 nsew power bidirectional
rlabel metal4 s 451794 -7654 452414 711590 6 vdda1
port 556 nsew power bidirectional
rlabel metal4 s 487794 -7654 488414 711590 6 vdda1
port 556 nsew power bidirectional
rlabel metal4 s 523794 -7654 524414 711590 6 vdda1
port 556 nsew power bidirectional
rlabel metal4 s 559794 -7654 560414 711590 6 vdda1
port 556 nsew power bidirectional
rlabel metal5 s -8726 20866 592650 21486 6 vdda1
port 556 nsew power bidirectional
rlabel metal5 s -8726 56866 592650 57486 6 vdda1
port 556 nsew power bidirectional
rlabel metal5 s -8726 92866 592650 93486 6 vdda1
port 556 nsew power bidirectional
rlabel metal5 s -8726 128866 592650 129486 6 vdda1
port 556 nsew power bidirectional
rlabel metal5 s -8726 164866 592650 165486 6 vdda1
port 556 nsew power bidirectional
rlabel metal5 s -8726 200866 592650 201486 6 vdda1
port 556 nsew power bidirectional
rlabel metal5 s -8726 236866 592650 237486 6 vdda1
port 556 nsew power bidirectional
rlabel metal5 s -8726 272866 592650 273486 6 vdda1
port 556 nsew power bidirectional
rlabel metal5 s -8726 308866 592650 309486 6 vdda1
port 556 nsew power bidirectional
rlabel metal5 s -8726 344866 592650 345486 6 vdda1
port 556 nsew power bidirectional
rlabel metal5 s -8726 380866 592650 381486 6 vdda1
port 556 nsew power bidirectional
rlabel metal5 s -8726 416866 592650 417486 6 vdda1
port 556 nsew power bidirectional
rlabel metal5 s -8726 452866 592650 453486 6 vdda1
port 556 nsew power bidirectional
rlabel metal5 s -8726 488866 592650 489486 6 vdda1
port 556 nsew power bidirectional
rlabel metal5 s -8726 524866 592650 525486 6 vdda1
port 556 nsew power bidirectional
rlabel metal5 s -8726 560866 592650 561486 6 vdda1
port 556 nsew power bidirectional
rlabel metal5 s -8726 596866 592650 597486 6 vdda1
port 556 nsew power bidirectional
rlabel metal5 s -8726 632866 592650 633486 6 vdda1
port 556 nsew power bidirectional
rlabel metal5 s -8726 668866 592650 669486 6 vdda1
port 556 nsew power bidirectional
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 557 nsew power bidirectional
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 557 nsew power bidirectional
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 557 nsew power bidirectional
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 557 nsew power bidirectional
rlabel metal4 s 28794 -7654 29414 711590 6 vdda2
port 557 nsew power bidirectional
rlabel metal4 s 64794 -7654 65414 711590 6 vdda2
port 557 nsew power bidirectional
rlabel metal4 s 100794 -7654 101414 711590 6 vdda2
port 557 nsew power bidirectional
rlabel metal4 s 136794 -7654 137414 78000 6 vdda2
port 557 nsew power bidirectional
rlabel metal4 s 136794 262000 137414 711590 6 vdda2
port 557 nsew power bidirectional
rlabel metal4 s 172794 -7654 173414 78000 6 vdda2
port 557 nsew power bidirectional
rlabel metal4 s 172794 262000 173414 711590 6 vdda2
port 557 nsew power bidirectional
rlabel metal4 s 208794 -7654 209414 711590 6 vdda2
port 557 nsew power bidirectional
rlabel metal4 s 244794 -7654 245414 711590 6 vdda2
port 557 nsew power bidirectional
rlabel metal4 s 280794 -7654 281414 711590 6 vdda2
port 557 nsew power bidirectional
rlabel metal4 s 316794 -7654 317414 711590 6 vdda2
port 557 nsew power bidirectional
rlabel metal4 s 352794 -7654 353414 711590 6 vdda2
port 557 nsew power bidirectional
rlabel metal4 s 388794 -7654 389414 711590 6 vdda2
port 557 nsew power bidirectional
rlabel metal4 s 424794 -7654 425414 711590 6 vdda2
port 557 nsew power bidirectional
rlabel metal4 s 460794 -7654 461414 711590 6 vdda2
port 557 nsew power bidirectional
rlabel metal4 s 496794 -7654 497414 711590 6 vdda2
port 557 nsew power bidirectional
rlabel metal4 s 532794 -7654 533414 711590 6 vdda2
port 557 nsew power bidirectional
rlabel metal4 s 568794 -7654 569414 711590 6 vdda2
port 557 nsew power bidirectional
rlabel metal5 s -8726 29866 592650 30486 6 vdda2
port 557 nsew power bidirectional
rlabel metal5 s -8726 65866 592650 66486 6 vdda2
port 557 nsew power bidirectional
rlabel metal5 s -8726 101866 592650 102486 6 vdda2
port 557 nsew power bidirectional
rlabel metal5 s -8726 137866 592650 138486 6 vdda2
port 557 nsew power bidirectional
rlabel metal5 s -8726 173866 592650 174486 6 vdda2
port 557 nsew power bidirectional
rlabel metal5 s -8726 209866 592650 210486 6 vdda2
port 557 nsew power bidirectional
rlabel metal5 s -8726 245866 592650 246486 6 vdda2
port 557 nsew power bidirectional
rlabel metal5 s -8726 281866 592650 282486 6 vdda2
port 557 nsew power bidirectional
rlabel metal5 s -8726 317866 592650 318486 6 vdda2
port 557 nsew power bidirectional
rlabel metal5 s -8726 353866 592650 354486 6 vdda2
port 557 nsew power bidirectional
rlabel metal5 s -8726 389866 592650 390486 6 vdda2
port 557 nsew power bidirectional
rlabel metal5 s -8726 425866 592650 426486 6 vdda2
port 557 nsew power bidirectional
rlabel metal5 s -8726 461866 592650 462486 6 vdda2
port 557 nsew power bidirectional
rlabel metal5 s -8726 497866 592650 498486 6 vdda2
port 557 nsew power bidirectional
rlabel metal5 s -8726 533866 592650 534486 6 vdda2
port 557 nsew power bidirectional
rlabel metal5 s -8726 569866 592650 570486 6 vdda2
port 557 nsew power bidirectional
rlabel metal5 s -8726 605866 592650 606486 6 vdda2
port 557 nsew power bidirectional
rlabel metal5 s -8726 641866 592650 642486 6 vdda2
port 557 nsew power bidirectional
rlabel metal5 s -8726 677866 592650 678486 6 vdda2
port 557 nsew power bidirectional
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 558 nsew ground bidirectional
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 558 nsew ground bidirectional
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 558 nsew ground bidirectional
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 558 nsew ground bidirectional
rlabel metal4 s 24294 -7654 24914 711590 6 vssa1
port 558 nsew ground bidirectional
rlabel metal4 s 60294 -7654 60914 711590 6 vssa1
port 558 nsew ground bidirectional
rlabel metal4 s 96294 -7654 96914 711590 6 vssa1
port 558 nsew ground bidirectional
rlabel metal4 s 132294 -7654 132914 78000 6 vssa1
port 558 nsew ground bidirectional
rlabel metal4 s 132294 262000 132914 711590 6 vssa1
port 558 nsew ground bidirectional
rlabel metal4 s 168294 -7654 168914 78000 6 vssa1
port 558 nsew ground bidirectional
rlabel metal4 s 168294 262000 168914 711590 6 vssa1
port 558 nsew ground bidirectional
rlabel metal4 s 204294 -7654 204914 711590 6 vssa1
port 558 nsew ground bidirectional
rlabel metal4 s 240294 -7654 240914 711590 6 vssa1
port 558 nsew ground bidirectional
rlabel metal4 s 276294 -7654 276914 711590 6 vssa1
port 558 nsew ground bidirectional
rlabel metal4 s 312294 -7654 312914 711590 6 vssa1
port 558 nsew ground bidirectional
rlabel metal4 s 348294 -7654 348914 711590 6 vssa1
port 558 nsew ground bidirectional
rlabel metal4 s 384294 -7654 384914 711590 6 vssa1
port 558 nsew ground bidirectional
rlabel metal4 s 420294 -7654 420914 711590 6 vssa1
port 558 nsew ground bidirectional
rlabel metal4 s 456294 -7654 456914 711590 6 vssa1
port 558 nsew ground bidirectional
rlabel metal4 s 492294 -7654 492914 711590 6 vssa1
port 558 nsew ground bidirectional
rlabel metal4 s 528294 -7654 528914 711590 6 vssa1
port 558 nsew ground bidirectional
rlabel metal4 s 564294 -7654 564914 711590 6 vssa1
port 558 nsew ground bidirectional
rlabel metal5 s -8726 25366 592650 25986 6 vssa1
port 558 nsew ground bidirectional
rlabel metal5 s -8726 61366 592650 61986 6 vssa1
port 558 nsew ground bidirectional
rlabel metal5 s -8726 97366 592650 97986 6 vssa1
port 558 nsew ground bidirectional
rlabel metal5 s -8726 133366 592650 133986 6 vssa1
port 558 nsew ground bidirectional
rlabel metal5 s -8726 169366 592650 169986 6 vssa1
port 558 nsew ground bidirectional
rlabel metal5 s -8726 205366 592650 205986 6 vssa1
port 558 nsew ground bidirectional
rlabel metal5 s -8726 241366 592650 241986 6 vssa1
port 558 nsew ground bidirectional
rlabel metal5 s -8726 277366 592650 277986 6 vssa1
port 558 nsew ground bidirectional
rlabel metal5 s -8726 313366 592650 313986 6 vssa1
port 558 nsew ground bidirectional
rlabel metal5 s -8726 349366 592650 349986 6 vssa1
port 558 nsew ground bidirectional
rlabel metal5 s -8726 385366 592650 385986 6 vssa1
port 558 nsew ground bidirectional
rlabel metal5 s -8726 421366 592650 421986 6 vssa1
port 558 nsew ground bidirectional
rlabel metal5 s -8726 457366 592650 457986 6 vssa1
port 558 nsew ground bidirectional
rlabel metal5 s -8726 493366 592650 493986 6 vssa1
port 558 nsew ground bidirectional
rlabel metal5 s -8726 529366 592650 529986 6 vssa1
port 558 nsew ground bidirectional
rlabel metal5 s -8726 565366 592650 565986 6 vssa1
port 558 nsew ground bidirectional
rlabel metal5 s -8726 601366 592650 601986 6 vssa1
port 558 nsew ground bidirectional
rlabel metal5 s -8726 637366 592650 637986 6 vssa1
port 558 nsew ground bidirectional
rlabel metal5 s -8726 673366 592650 673986 6 vssa1
port 558 nsew ground bidirectional
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 559 nsew ground bidirectional
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 559 nsew ground bidirectional
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 559 nsew ground bidirectional
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 559 nsew ground bidirectional
rlabel metal4 s 33294 -7654 33914 711590 6 vssa2
port 559 nsew ground bidirectional
rlabel metal4 s 69294 -7654 69914 711590 6 vssa2
port 559 nsew ground bidirectional
rlabel metal4 s 105294 -7654 105914 711590 6 vssa2
port 559 nsew ground bidirectional
rlabel metal4 s 141294 -7654 141914 78000 6 vssa2
port 559 nsew ground bidirectional
rlabel metal4 s 141294 142000 141914 198000 6 vssa2
port 559 nsew ground bidirectional
rlabel metal4 s 141294 262000 141914 711590 6 vssa2
port 559 nsew ground bidirectional
rlabel metal4 s 177294 -7654 177914 78000 6 vssa2
port 559 nsew ground bidirectional
rlabel metal4 s 177294 142000 177914 198000 6 vssa2
port 559 nsew ground bidirectional
rlabel metal4 s 177294 262000 177914 711590 6 vssa2
port 559 nsew ground bidirectional
rlabel metal4 s 213294 -7654 213914 711590 6 vssa2
port 559 nsew ground bidirectional
rlabel metal4 s 249294 -7654 249914 711590 6 vssa2
port 559 nsew ground bidirectional
rlabel metal4 s 285294 -7654 285914 711590 6 vssa2
port 559 nsew ground bidirectional
rlabel metal4 s 321294 -7654 321914 711590 6 vssa2
port 559 nsew ground bidirectional
rlabel metal4 s 357294 -7654 357914 711590 6 vssa2
port 559 nsew ground bidirectional
rlabel metal4 s 393294 -7654 393914 711590 6 vssa2
port 559 nsew ground bidirectional
rlabel metal4 s 429294 -7654 429914 711590 6 vssa2
port 559 nsew ground bidirectional
rlabel metal4 s 465294 -7654 465914 711590 6 vssa2
port 559 nsew ground bidirectional
rlabel metal4 s 501294 -7654 501914 711590 6 vssa2
port 559 nsew ground bidirectional
rlabel metal4 s 537294 -7654 537914 711590 6 vssa2
port 559 nsew ground bidirectional
rlabel metal4 s 573294 -7654 573914 711590 6 vssa2
port 559 nsew ground bidirectional
rlabel metal5 s -8726 34366 592650 34986 6 vssa2
port 559 nsew ground bidirectional
rlabel metal5 s -8726 70366 592650 70986 6 vssa2
port 559 nsew ground bidirectional
rlabel metal5 s -8726 106366 592650 106986 6 vssa2
port 559 nsew ground bidirectional
rlabel metal5 s -8726 142366 592650 142986 6 vssa2
port 559 nsew ground bidirectional
rlabel metal5 s -8726 178366 592650 178986 6 vssa2
port 559 nsew ground bidirectional
rlabel metal5 s -8726 214366 592650 214986 6 vssa2
port 559 nsew ground bidirectional
rlabel metal5 s -8726 250366 592650 250986 6 vssa2
port 559 nsew ground bidirectional
rlabel metal5 s -8726 286366 592650 286986 6 vssa2
port 559 nsew ground bidirectional
rlabel metal5 s -8726 322366 592650 322986 6 vssa2
port 559 nsew ground bidirectional
rlabel metal5 s -8726 358366 592650 358986 6 vssa2
port 559 nsew ground bidirectional
rlabel metal5 s -8726 394366 592650 394986 6 vssa2
port 559 nsew ground bidirectional
rlabel metal5 s -8726 430366 592650 430986 6 vssa2
port 559 nsew ground bidirectional
rlabel metal5 s -8726 466366 592650 466986 6 vssa2
port 559 nsew ground bidirectional
rlabel metal5 s -8726 502366 592650 502986 6 vssa2
port 559 nsew ground bidirectional
rlabel metal5 s -8726 538366 592650 538986 6 vssa2
port 559 nsew ground bidirectional
rlabel metal5 s -8726 574366 592650 574986 6 vssa2
port 559 nsew ground bidirectional
rlabel metal5 s -8726 610366 592650 610986 6 vssa2
port 559 nsew ground bidirectional
rlabel metal5 s -8726 646366 592650 646986 6 vssa2
port 559 nsew ground bidirectional
rlabel metal5 s -8726 682366 592650 682986 6 vssa2
port 559 nsew ground bidirectional
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 560 nsew ground bidirectional
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 560 nsew ground bidirectional
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 560 nsew ground bidirectional
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 560 nsew ground bidirectional
rlabel metal4 s 6294 -7654 6914 711590 6 vssd1
port 560 nsew ground bidirectional
rlabel metal4 s 42294 -7654 42914 711590 6 vssd1
port 560 nsew ground bidirectional
rlabel metal4 s 78294 -7654 78914 711590 6 vssd1
port 560 nsew ground bidirectional
rlabel metal4 s 114294 -7654 114914 711590 6 vssd1
port 560 nsew ground bidirectional
rlabel metal4 s 150294 -7654 150914 78000 6 vssd1
port 560 nsew ground bidirectional
rlabel metal4 s 150294 142000 150914 198000 6 vssd1
port 560 nsew ground bidirectional
rlabel metal4 s 150294 262000 150914 711590 6 vssd1
port 560 nsew ground bidirectional
rlabel metal4 s 186294 -7654 186914 78000 6 vssd1
port 560 nsew ground bidirectional
rlabel metal4 s 186294 142000 186914 198000 6 vssd1
port 560 nsew ground bidirectional
rlabel metal4 s 186294 262000 186914 711590 6 vssd1
port 560 nsew ground bidirectional
rlabel metal4 s 222294 -7654 222914 711590 6 vssd1
port 560 nsew ground bidirectional
rlabel metal4 s 258294 -7654 258914 711590 6 vssd1
port 560 nsew ground bidirectional
rlabel metal4 s 294294 -7654 294914 711590 6 vssd1
port 560 nsew ground bidirectional
rlabel metal4 s 330294 -7654 330914 711590 6 vssd1
port 560 nsew ground bidirectional
rlabel metal4 s 366294 -7654 366914 711590 6 vssd1
port 560 nsew ground bidirectional
rlabel metal4 s 402294 -7654 402914 711590 6 vssd1
port 560 nsew ground bidirectional
rlabel metal4 s 438294 -7654 438914 711590 6 vssd1
port 560 nsew ground bidirectional
rlabel metal4 s 474294 -7654 474914 711590 6 vssd1
port 560 nsew ground bidirectional
rlabel metal4 s 510294 -7654 510914 711590 6 vssd1
port 560 nsew ground bidirectional
rlabel metal4 s 546294 -7654 546914 711590 6 vssd1
port 560 nsew ground bidirectional
rlabel metal4 s 582294 -7654 582914 711590 6 vssd1
port 560 nsew ground bidirectional
rlabel metal5 s -8726 7366 592650 7986 6 vssd1
port 560 nsew ground bidirectional
rlabel metal5 s -8726 43366 592650 43986 6 vssd1
port 560 nsew ground bidirectional
rlabel metal5 s -8726 79366 592650 79986 6 vssd1
port 560 nsew ground bidirectional
rlabel metal5 s -8726 115366 592650 115986 6 vssd1
port 560 nsew ground bidirectional
rlabel metal5 s -8726 151366 592650 151986 6 vssd1
port 560 nsew ground bidirectional
rlabel metal5 s -8726 187366 592650 187986 6 vssd1
port 560 nsew ground bidirectional
rlabel metal5 s -8726 223366 592650 223986 6 vssd1
port 560 nsew ground bidirectional
rlabel metal5 s -8726 259366 592650 259986 6 vssd1
port 560 nsew ground bidirectional
rlabel metal5 s -8726 295366 592650 295986 6 vssd1
port 560 nsew ground bidirectional
rlabel metal5 s -8726 331366 592650 331986 6 vssd1
port 560 nsew ground bidirectional
rlabel metal5 s -8726 367366 592650 367986 6 vssd1
port 560 nsew ground bidirectional
rlabel metal5 s -8726 403366 592650 403986 6 vssd1
port 560 nsew ground bidirectional
rlabel metal5 s -8726 439366 592650 439986 6 vssd1
port 560 nsew ground bidirectional
rlabel metal5 s -8726 475366 592650 475986 6 vssd1
port 560 nsew ground bidirectional
rlabel metal5 s -8726 511366 592650 511986 6 vssd1
port 560 nsew ground bidirectional
rlabel metal5 s -8726 547366 592650 547986 6 vssd1
port 560 nsew ground bidirectional
rlabel metal5 s -8726 583366 592650 583986 6 vssd1
port 560 nsew ground bidirectional
rlabel metal5 s -8726 619366 592650 619986 6 vssd1
port 560 nsew ground bidirectional
rlabel metal5 s -8726 655366 592650 655986 6 vssd1
port 560 nsew ground bidirectional
rlabel metal5 s -8726 691366 592650 691986 6 vssd1
port 560 nsew ground bidirectional
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 561 nsew ground bidirectional
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 561 nsew ground bidirectional
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 561 nsew ground bidirectional
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 561 nsew ground bidirectional
rlabel metal4 s 15294 -7654 15914 711590 6 vssd2
port 561 nsew ground bidirectional
rlabel metal4 s 51294 -7654 51914 711590 6 vssd2
port 561 nsew ground bidirectional
rlabel metal4 s 87294 -7654 87914 711590 6 vssd2
port 561 nsew ground bidirectional
rlabel metal4 s 123294 -7654 123914 78000 6 vssd2
port 561 nsew ground bidirectional
rlabel metal4 s 123294 142000 123914 198000 6 vssd2
port 561 nsew ground bidirectional
rlabel metal4 s 123294 262000 123914 711590 6 vssd2
port 561 nsew ground bidirectional
rlabel metal4 s 159294 -7654 159914 78000 6 vssd2
port 561 nsew ground bidirectional
rlabel metal4 s 159294 142000 159914 198000 6 vssd2
port 561 nsew ground bidirectional
rlabel metal4 s 159294 262000 159914 711590 6 vssd2
port 561 nsew ground bidirectional
rlabel metal4 s 195294 -7654 195914 711590 6 vssd2
port 561 nsew ground bidirectional
rlabel metal4 s 231294 -7654 231914 711590 6 vssd2
port 561 nsew ground bidirectional
rlabel metal4 s 267294 -7654 267914 711590 6 vssd2
port 561 nsew ground bidirectional
rlabel metal4 s 303294 -7654 303914 711590 6 vssd2
port 561 nsew ground bidirectional
rlabel metal4 s 339294 -7654 339914 711590 6 vssd2
port 561 nsew ground bidirectional
rlabel metal4 s 375294 -7654 375914 711590 6 vssd2
port 561 nsew ground bidirectional
rlabel metal4 s 411294 -7654 411914 711590 6 vssd2
port 561 nsew ground bidirectional
rlabel metal4 s 447294 -7654 447914 711590 6 vssd2
port 561 nsew ground bidirectional
rlabel metal4 s 483294 -7654 483914 711590 6 vssd2
port 561 nsew ground bidirectional
rlabel metal4 s 519294 -7654 519914 711590 6 vssd2
port 561 nsew ground bidirectional
rlabel metal4 s 555294 -7654 555914 711590 6 vssd2
port 561 nsew ground bidirectional
rlabel metal5 s -8726 16366 592650 16986 6 vssd2
port 561 nsew ground bidirectional
rlabel metal5 s -8726 52366 592650 52986 6 vssd2
port 561 nsew ground bidirectional
rlabel metal5 s -8726 88366 592650 88986 6 vssd2
port 561 nsew ground bidirectional
rlabel metal5 s -8726 124366 592650 124986 6 vssd2
port 561 nsew ground bidirectional
rlabel metal5 s -8726 160366 592650 160986 6 vssd2
port 561 nsew ground bidirectional
rlabel metal5 s -8726 196366 592650 196986 6 vssd2
port 561 nsew ground bidirectional
rlabel metal5 s -8726 232366 592650 232986 6 vssd2
port 561 nsew ground bidirectional
rlabel metal5 s -8726 268366 592650 268986 6 vssd2
port 561 nsew ground bidirectional
rlabel metal5 s -8726 304366 592650 304986 6 vssd2
port 561 nsew ground bidirectional
rlabel metal5 s -8726 340366 592650 340986 6 vssd2
port 561 nsew ground bidirectional
rlabel metal5 s -8726 376366 592650 376986 6 vssd2
port 561 nsew ground bidirectional
rlabel metal5 s -8726 412366 592650 412986 6 vssd2
port 561 nsew ground bidirectional
rlabel metal5 s -8726 448366 592650 448986 6 vssd2
port 561 nsew ground bidirectional
rlabel metal5 s -8726 484366 592650 484986 6 vssd2
port 561 nsew ground bidirectional
rlabel metal5 s -8726 520366 592650 520986 6 vssd2
port 561 nsew ground bidirectional
rlabel metal5 s -8726 556366 592650 556986 6 vssd2
port 561 nsew ground bidirectional
rlabel metal5 s -8726 592366 592650 592986 6 vssd2
port 561 nsew ground bidirectional
rlabel metal5 s -8726 628366 592650 628986 6 vssd2
port 561 nsew ground bidirectional
rlabel metal5 s -8726 664366 592650 664986 6 vssd2
port 561 nsew ground bidirectional
rlabel metal5 s -8726 700366 592650 700986 6 vssd2
port 561 nsew ground bidirectional
rlabel metal3 s 583520 256988 584960 257228 6 wb_clk_i
port 562 nsew signal input
rlabel metal3 s -960 348788 480 349028 4 wb_rst_i
port 563 nsew signal input
rlabel metal3 s 583520 385508 584960 385748 6 wbs_ack_o
port 564 nsew signal output
rlabel metal2 s 198342 703520 198454 704960 6 wbs_adr_i[0]
port 565 nsew signal input
rlabel metal2 s 54086 703520 54198 704960 6 wbs_adr_i[10]
port 566 nsew signal input
rlabel metal3 s -960 472548 480 472788 4 wbs_adr_i[11]
port 567 nsew signal input
rlabel metal2 s 64390 -960 64502 480 8 wbs_adr_i[12]
port 568 nsew signal input
rlabel metal3 s -960 360348 480 360588 4 wbs_adr_i[13]
port 569 nsew signal input
rlabel metal3 s 583520 662268 584960 662508 6 wbs_adr_i[14]
port 570 nsew signal input
rlabel metal3 s 583520 613988 584960 614228 6 wbs_adr_i[15]
port 571 nsew signal input
rlabel metal2 s 443706 -960 443818 480 8 wbs_adr_i[16]
port 572 nsew signal input
rlabel metal3 s 583520 557548 584960 557788 6 wbs_adr_i[17]
port 573 nsew signal input
rlabel metal3 s 583520 345388 584960 345628 6 wbs_adr_i[18]
port 574 nsew signal input
rlabel metal3 s 583520 88348 584960 88588 6 wbs_adr_i[19]
port 575 nsew signal input
rlabel metal2 s 206070 703520 206182 704960 6 wbs_adr_i[1]
port 576 nsew signal input
rlabel metal2 s 406998 703520 407110 704960 6 wbs_adr_i[20]
port 577 nsew signal input
rlabel metal2 s 390898 -960 391010 480 8 wbs_adr_i[21]
port 578 nsew signal input
rlabel metal2 s 557694 -960 557806 480 8 wbs_adr_i[22]
port 579 nsew signal input
rlabel metal3 s 583520 276708 584960 276948 6 wbs_adr_i[23]
port 580 nsew signal input
rlabel metal3 s -960 552788 480 553028 4 wbs_adr_i[24]
port 581 nsew signal input
rlabel metal2 s 375442 -960 375554 480 8 wbs_adr_i[25]
port 582 nsew signal input
rlabel metal2 s 72118 -960 72230 480 8 wbs_adr_i[26]
port 583 nsew signal input
rlabel metal3 s -960 19668 480 19908 4 wbs_adr_i[27]
port 584 nsew signal input
rlabel metal3 s 583520 525588 584960 525828 6 wbs_adr_i[28]
port 585 nsew signal input
rlabel metal2 s 498446 703520 498558 704960 6 wbs_adr_i[29]
port 586 nsew signal input
rlabel metal2 s 265318 -960 265430 480 8 wbs_adr_i[2]
port 587 nsew signal input
rlabel metal2 s 331006 703520 331118 704960 6 wbs_adr_i[30]
port 588 nsew signal input
rlabel metal3 s 583520 405228 584960 405468 6 wbs_adr_i[31]
port 589 nsew signal input
rlabel metal2 s 531290 -960 531402 480 8 wbs_adr_i[3]
port 590 nsew signal input
rlabel metal2 s 323922 703520 324034 704960 6 wbs_adr_i[4]
port 591 nsew signal input
rlabel metal3 s -960 108068 480 108308 4 wbs_adr_i[5]
port 592 nsew signal input
rlabel metal2 s 216374 -960 216486 480 8 wbs_adr_i[6]
port 593 nsew signal input
rlabel metal2 s 34122 -960 34234 480 8 wbs_adr_i[7]
port 594 nsew signal input
rlabel metal3 s 583520 96508 584960 96748 6 wbs_adr_i[8]
port 595 nsew signal input
rlabel metal3 s 583520 288948 584960 289188 6 wbs_adr_i[9]
port 596 nsew signal input
rlabel metal2 s 27682 703520 27794 704960 6 wbs_cyc_i
port 597 nsew signal input
rlabel metal2 s 574438 703520 574550 704960 6 wbs_dat_i[0]
port 598 nsew signal input
rlabel metal3 s -960 356268 480 356508 4 wbs_dat_i[10]
port 599 nsew signal input
rlabel metal3 s -960 408628 480 408868 4 wbs_dat_i[11]
port 600 nsew signal input
rlabel metal3 s -960 388228 480 388468 4 wbs_dat_i[12]
port 601 nsew signal input
rlabel metal2 s 26394 -960 26506 480 8 wbs_dat_i[13]
port 602 nsew signal input
rlabel metal2 s 144246 -960 144358 480 8 wbs_dat_i[14]
port 603 nsew signal input
rlabel metal3 s 583520 457588 584960 457828 6 wbs_dat_i[15]
port 604 nsew signal input
rlabel metal3 s -960 43468 480 43708 4 wbs_dat_i[16]
port 605 nsew signal input
rlabel metal2 s 293010 703520 293122 704960 6 wbs_dat_i[17]
port 606 nsew signal input
rlabel metal2 s 456586 703520 456698 704960 6 wbs_dat_i[18]
port 607 nsew signal input
rlabel metal3 s -960 577268 480 577508 4 wbs_dat_i[19]
port 608 nsew signal input
rlabel metal2 s 102386 -960 102498 480 8 wbs_dat_i[1]
port 609 nsew signal input
rlabel metal3 s 583520 505868 584960 506108 6 wbs_dat_i[20]
port 610 nsew signal input
rlabel metal2 s 479126 703520 479238 704960 6 wbs_dat_i[21]
port 611 nsew signal input
rlabel metal3 s -960 264468 480 264708 4 wbs_dat_i[22]
port 612 nsew signal input
rlabel metal3 s 583520 629628 584960 629868 6 wbs_dat_i[23]
port 613 nsew signal input
rlabel metal3 s 583520 309348 584960 309588 6 wbs_dat_i[24]
port 614 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 wbs_dat_i[25]
port 615 nsew signal input
rlabel metal2 s 410862 703520 410974 704960 6 wbs_dat_i[26]
port 616 nsew signal input
rlabel metal2 s 19954 703520 20066 704960 6 wbs_dat_i[27]
port 617 nsew signal input
rlabel metal2 s 208646 -960 208758 480 8 wbs_dat_i[28]
port 618 nsew signal input
rlabel metal3 s 583520 497708 584960 497948 6 wbs_dat_i[29]
port 619 nsew signal input
rlabel metal2 s 539018 -960 539130 480 8 wbs_dat_i[2]
port 620 nsew signal input
rlabel metal3 s 583520 280788 584960 281028 6 wbs_dat_i[30]
port 621 nsew signal input
rlabel metal3 s -960 248148 480 248388 4 wbs_dat_i[31]
port 622 nsew signal input
rlabel metal3 s 583520 100588 584960 100828 6 wbs_dat_i[3]
port 623 nsew signal input
rlabel metal2 s 106250 -960 106362 480 8 wbs_dat_i[4]
port 624 nsew signal input
rlabel metal2 s 326498 -960 326610 480 8 wbs_dat_i[5]
port 625 nsew signal input
rlabel metal3 s 583520 373268 584960 373508 6 wbs_dat_i[6]
port 626 nsew signal input
rlabel metal2 s 399914 703520 400026 704960 6 wbs_dat_i[7]
port 627 nsew signal input
rlabel metal3 s 583520 686068 584960 686308 6 wbs_dat_i[8]
port 628 nsew signal input
rlabel metal3 s 583520 104668 584960 104908 6 wbs_dat_i[9]
port 629 nsew signal input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_o[0]
port 630 nsew signal output
rlabel metal3 s 583520 461668 584960 461908 6 wbs_dat_o[10]
port 631 nsew signal output
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[11]
port 632 nsew signal output
rlabel metal3 s 583520 694228 584960 694468 6 wbs_dat_o[12]
port 633 nsew signal output
rlabel metal2 s 384458 703520 384570 704960 6 wbs_dat_o[13]
port 634 nsew signal output
rlabel metal3 s 583520 144788 584960 145028 6 wbs_dat_o[14]
port 635 nsew signal output
rlabel metal2 s 365138 703520 365250 704960 6 wbs_dat_o[15]
port 636 nsew signal output
rlabel metal2 s 436622 -960 436734 480 8 wbs_dat_o[16]
port 637 nsew signal output
rlabel metal3 s -960 135948 480 136188 4 wbs_dat_o[17]
port 638 nsew signal output
rlabel metal2 s 432758 -960 432870 480 8 wbs_dat_o[18]
port 639 nsew signal output
rlabel metal2 s -10 -960 102 480 8 wbs_dat_o[19]
port 640 nsew signal output
rlabel metal2 s 508750 -960 508862 480 8 wbs_dat_o[1]
port 641 nsew signal output
rlabel metal3 s -960 256308 480 256548 4 wbs_dat_o[20]
port 642 nsew signal output
rlabel metal3 s -960 524908 480 525148 4 wbs_dat_o[21]
port 643 nsew signal output
rlabel metal2 s 92082 703520 92194 704960 6 wbs_dat_o[22]
port 644 nsew signal output
rlabel metal3 s -960 167908 480 168148 4 wbs_dat_o[23]
port 645 nsew signal output
rlabel metal2 s 132654 -960 132766 480 8 wbs_dat_o[24]
port 646 nsew signal output
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_o[25]
port 647 nsew signal output
rlabel metal2 s 255014 703520 255126 704960 6 wbs_dat_o[26]
port 648 nsew signal output
rlabel metal2 s 114622 703520 114734 704960 6 wbs_dat_o[27]
port 649 nsew signal output
rlabel metal2 s 345174 -960 345286 480 8 wbs_dat_o[28]
port 650 nsew signal output
rlabel metal2 s 369002 703520 369114 704960 6 wbs_dat_o[29]
port 651 nsew signal output
rlabel metal3 s 583520 240668 584960 240908 6 wbs_dat_o[2]
port 652 nsew signal output
rlabel metal3 s -960 404548 480 404788 4 wbs_dat_o[30]
port 653 nsew signal output
rlabel metal3 s 583520 569788 584960 570028 6 wbs_dat_o[31]
port 654 nsew signal output
rlabel metal2 s 140382 -960 140494 480 8 wbs_dat_o[3]
port 655 nsew signal output
rlabel metal2 s 242778 -960 242890 480 8 wbs_dat_o[4]
port 656 nsew signal output
rlabel metal3 s -960 35988 480 36228 4 wbs_dat_o[5]
port 657 nsew signal output
rlabel metal3 s 583520 541908 584960 542148 6 wbs_dat_o[6]
port 658 nsew signal output
rlabel metal2 s 383170 -960 383282 480 8 wbs_dat_o[7]
port 659 nsew signal output
rlabel metal2 s 358054 703520 358166 704960 6 wbs_dat_o[8]
port 660 nsew signal output
rlabel metal2 s 354190 703520 354302 704960 6 wbs_dat_o[9]
port 661 nsew signal output
rlabel metal3 s -960 601068 480 601308 4 wbs_sel_i[0]
port 662 nsew signal input
rlabel metal2 s 16090 703520 16202 704960 6 wbs_sel_i[1]
port 663 nsew signal input
rlabel metal2 s 455298 -960 455410 480 8 wbs_sel_i[2]
port 664 nsew signal input
rlabel metal3 s -960 140028 480 140268 4 wbs_sel_i[3]
port 665 nsew signal input
rlabel metal3 s -960 541228 480 541468 4 wbs_stb_i
port 666 nsew signal input
rlabel metal3 s 583520 369188 584960 369428 6 wbs_we_i
port 667 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 7913910
string GDS_FILE /home/mxmont/Documents/Universidad/IC-UBB/MixPix/CARAVEL_WRAPPER/MixPix/openlane/user_project_wrapper/runs/22_10_28_22_25/results/signoff/user_project_wrapper.magic.gds
string GDS_START 4284704
<< end >>

